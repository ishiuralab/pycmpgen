module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [14:0] src16;
    reg [13:0] src17;
    reg [12:0] src18;
    reg [11:0] src19;
    reg [10:0] src20;
    reg [9:0] src21;
    reg [8:0] src22;
    reg [7:0] src23;
    reg [6:0] src24;
    reg [5:0] src25;
    reg [4:0] src26;
    reg [3:0] src27;
    reg [2:0] src28;
    reg [1:0] src29;
    reg [0:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3])<<27) + ((src28[0] + src28[1] + src28[2])<<28) + ((src29[0] + src29[1])<<29) + ((src30[0])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe76232cd64a7bf3b37de3c88c980134bb83797d1a16c4821861c9fb2d4e27f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11a6a56639c187d042023b8730ed175ef3be986c7c228c7d71d3b4544cd74dbb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b8fde9cdb65626fc4f11e48c0f9a89d6873c90a9b6e0bb49ec07ab3034d1588;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dd16593e1431da7276023bee461ca01d3573266ddf67fd78808ebd1792603e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hacacf73d915d79ec8fbc6121acf7ea8482dafa7aae4d48ec59457bd53e4d89b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfffe1125d485b0d6938fe668141d4b4e177db969e4e92cc14172fc80a3102161;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70c59588211536b09c581e756ffcae86f5217d31c7d89b44d681d790724a4fc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h300a6b2895858bccc7156dca81b56528134d74d1d19d42fe501b08b76a27b7b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78d7740df76ff433a9224e64488e14fd66c0dffe8ba9e9c2cd6bab9996de2691;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha963a6f84dab604397131ee62a8e1700caf1665741f764b9c35a1a52070e2a9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9eb6156ef3f327b9fca9528a2a1e3e3c4331bce15ae6f0b55771ae5a0134aed6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1dd724fa518177d4000d047996709f90f71544267843ff0f4278736596e0e985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39bf342da518e087148ab934f9498510a91afeaeece7f5cb2387466961c01972;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd65d8d2a74081c0f089cc45128535d34ab4679f59aa7718f969259b500f2051c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hadd7204e39c20135d906c4bcd280ea2345f50d7a9ed7d38a55a3804ab738f1c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdf7552554d2eef869656340729d94b1e4238dd80e4adf675aadc142c88a4cb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7010c2431a67e2302025bc82224ea4bd0bda9f140bd351da81b592a4a96fc086;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f84ba4014c6d7e0cebd80a3be6d3e0b390f773b2907edd0305bf3e40358e0c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he888991b007ec6b1ab4fb79b597a33cfcc900041a3c4b17b862e791c15c14b63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc7fac3afce4af4afcdb6973b11e40477413fd0fe0174eff254eea0646ae2d7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd710482bde6c13655bc05f39897fb50e2e0c35a9d766e9c1389dd88f99f8c24c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c8829050dd9b8f3a44570ba3df7975a898f23301ce59444a8ce7293bca2690f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5084845a8cb25c136a7c365b4bdd2a39147b7a1f4913f39ad5634ee000c093de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56f4099e14b9f5d4a4ced0a8fe680f04f0be3eceef7fa740822e26987efed883;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63ef3941c3755ef86ff6d92f9495140d6d7d8f7a846f80f0da548ad8714dcd43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9be7acba31b32196c56fabcf379b4d1eb89827df07e6bebb54468a6439db7760;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd9ed15dc666955d060428246be7d3f0a0f6f0ada5ef284157abdddcc54aa727;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h438bce784bcad15b26064f92e01a3f3183b7b646b7908c97179ce25bf1e1114c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb10430aecf31bf3e1d2a8238152ca5807c4016e4e2ee6a8fb60cd4224fde5206;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf41248c410d5b9a4edabdc1b8fbe94130f06be9df86bf0c0cf38b22ce1525207;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b28294a2bcfe022cfa80584cfe2f3665a3c94e39a08beb6993dc8244e48cc0f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78bfbd7a9cfabe5b61fb2d7493589f5a267a239c80431f79f6039ad4ab9d4122;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb88b94d88aca1d1078cb23aaa397aa3bc46c7f2947d0daaae4542438eb9ba01d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha703276933f78153b1f3c3a17a9018531fa4e078dc619ba508627205d8f0ac7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2a6702e132f1dbef66c101be72039a53628aa224fd7db9513843238431d14f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75c7315b2afb69b775a1a189888fa0bb1b6df2f92ad1def3a8a8b8bbe14126c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1642e3332bab8ef3f78f458078b9ee542274f4d4b7b80c14081df7dd42e0d926;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1560838d3131dee930aac84bfac02b108f9150588cbf02009bb5074bbff1513;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haffdd879f30feda8ae7534955011e4ce8f5ce962f623b27781c2e1f1efaf1748;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67193da2369b14694f04f94c7a77ec795f8d1e0f0b5ad253ce7d1d98f3e4783b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd22a8aee530157ad38c6a02bed9f118e597b335e4befce50e328c80a66f9ae54;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h269a7d8e60d1e3ddf571ecfb988826f7ad54ef21f68e8ff3eea900e144f9b4cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h177c33e996d87670dca3d2b82d521802c9b43d0da8589565b3a0e0393f903f0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4615cab00ee30b16f2dfac026f690477eaf6feae719559a0f332d766e69c393e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ea215e362bf586441e1a3bb228d9ea5233b5a3059cf2dd537d745fec0f349ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd108f35f39075e07b8e5bb4a536d95d383f4f6f26bc5c4679ba8bdaadcff5ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97107db243ada118e9c70f3799082f91598183e7042cadf07140424e1a2517b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha95f796c290e3cf7388d1c50335d26a4c54b1dc3cb73a93a64a0550181c3f145;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63383065164dd6c15697c272538d2bf1e2256db16fc862532a11c844634dcb14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h509cadd08a57f0c6653ec8ba221f38149013f3cb6e1da2c7ec6660aed23d5e01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd15e762ae14f4a6b18c71dd81b6e34512e2f2bf05410c228470b8848f9ec0b88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62cd6482a146f7f1e1038684dc294f06589fbefedcd5d485d71a7aea87707724;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a731c81b13ccd97f646d91c8e171888747370e1a4102a0e86040fa54179a949;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42709130ee9f48acf79242eafe0c4970beb512eedc964d064f1d47f7344a840e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9e84e9582fd311242fb1cde832aa2fbb97f04b2fc8aa48184b80524230e2242;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2b1140a750240fb796ada55bf4ab47f2cb3fafd3090ddb5fcd1787d791d2332;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1f050d3bb42f797780e68d6184cf79431c6e840fb285633e858e00dd43fc3d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50914779a6377965f0a64d4f122836d6f6f0c1be52f203838937313bde843914;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbb56af4891181c439d1374608c35b2265b96b4fa1900de2af420106882f532a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c28c9deb973587b7ed8c77b9ed15134441a347550773ed128cb8c3cd69de75f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3629b66e4d166d6fbc5185a7e5bba2eb5ad53c331d4b66a7e4b70499aca7ef43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6697d0cc37298452ff3cdc21513b3a5218575408f81bd06fb2b2f05710f95215;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a8bc1603c2c84aa8c0992a3e740a33e35ffbcb0c896e95d27ed769d9bb88a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3b3a97c84636eceafddeac93f21507e93723efae1d922a5addf0712dedecbdb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1513f785c0a7cbcb188130e32aea5b59d1485e5ea6c21f15476490935cf991d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e7bfd02fb5ff3dcf784dae6bc708d838c1bcb30b7f9a6c04ae4f04061872322;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h571c525a24f7e6bdefa636d2b2a428b4367ba1532ef84a7f765f5030317ac7c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5161c5ce62d5ce604abdc5335fb060a5b4e7aee010468b6156dd5445aa330471;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3831c1eeebb3b004157bf5bc2a6bbe3e0803a04bfa92417d4b87104ec10b9f15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h506f54e5d2624b88c0345af126af610ea404356c90b5cd5eeb1ac1335b8d13ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fff700d84350f3c0ee3357c32e60f23f517842d0ecf35844d9ad56edd7b10b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44040cc710e87b19fe1edfa8fd5b4d98d42f94386cce72a0f7541101ee9afd7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e985fbdf68b45da7f6eade5a944aeccf36dea0df8f3357c0acb790683890a62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28d97291c3e4ddbbf99e765a628878f9b720e9a1439ad10707416758bc25a9b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h685711e9490149b74820c57872e8c104e74567ef8c35f5869081fbcbadac5d0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a1700a9d683a746cc15f1f22a75d08b59e4bca146da96abb90e914781ac10bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72924b438f5a6948703bb53297913c7830bd65402271225988a4603180cf1aff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98bee16fee1d2b03465778fa74623d8745701fcfe714dc7a633f7bb8555326d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21c82e86bed148a6e6ae2897febc6a0d1fbfc9e68863731292bbde8f8075ac35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3a3acc60dcf6eee23287bb154bde7cd8e9ab82edce779b3a8882eed19abbf19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac9e0ac13d39fbd88c48f6c4f3e8ac54f0498fc2ddc9a220091429093d96b1cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1309f606adf114edfec262a26bbe7e4b6876207c87f993882af1ba5b95c8d38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h646e6671b3a4f7a6036942265acb75c5f6f93807833341adc06800efa5023d8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5b2374dc1c4c4404009bdd84604fbaee2601c68316ac580f40dd33497854c7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a15cc05eb38dcd44c3fa63fdece0b589f7acafa1bd801efb3dd694a33700357;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44aac88792be83796682ee292fda84bd747194a0f62084b8736fe477a5cbffb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30b3b5ed0949a9bf58bbffd6aa1cea4b9027c7a34bbfc5f1a8cf919accb429fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc653c64f4af6b3c5e56b8261b675130e136966d99c88e85ff4f85f1fe795ba24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5fdf226cfc1c740c7b73c65b37ff46faa00ba893cd9f66cd1dff0492a3d07d23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd87c6a43a5d4c5a7b433eebfeb95ac7dab42eabb9b1d1b3b52040e38222e0933;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h213e3f758f251de8e280982f513e97475dbdde6d2afb39825504350396cece8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe571763158073f0748d755c2439af821b87db79d35713e0eb998fa22af85bcf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33304acd83c1048eab01c8cfeea3d5f7a09f2edb5da51d2d7b2946dc7d4de051;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56796f05973ebb897ecf45bbbec807ea6325b3b73ffbbdd58a037a2c706001a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11b446db5b2bebe672523c3d20177f24aaf0c6b8cbf70062fbbc32be4a95c5a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4049dbf6ad73157515202d621f60aebff2c5be68db835d5fc21f929f963e9e7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0c831c431cd3aa7e9f786e8f90ae3e2d0d862d11d7d10052a6907a5d9b7670b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55ecf8fc70d0b4a695168c7729fbde768971f281d5ebad7825b3c4bf69399cda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93482d364edf21c81be73f899b59d4a64c40ed78828dcc37f58a14b58a0e5f43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h193ecd78631ee7f4101bccabb7018d4c142c99874e3e9f7cbbaa8027970dda4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeb217514da6a6f86fb5a869997215bef3edf01a0f0e3a496758be82b66928d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23af7528e7bb3bc830236ce1a74c4603dec42c24d28d58a19cd3593f0bb47420;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b40c2c6cb8e954861344e598ccf5505cec661c22ea504171da86fa542f34998;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb739a8a1c6512dfe5cb102a65927d00e584bf7096d6c20f7fd9ab6d6341d2eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda3b33372d72071eeca537f6a538b39074e7b9206ceccd39de10803fea5c69be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he670609a5ca190010e96dcbd56e137803e267e93078d7dca770209cd1336ada2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49f7a2c68b2b488b17ac59d9ee4709eb3d3529fd4a574ffcd3f0acee41e856dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb812ec998c642e683f5f9f6ecd585a9977aeaa1062437ce72f79c223eb5cb0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h668385bfe99069c23117874e46fbca24e27800bd1a0628252f6679fac5e165e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bbfb57c7e3f312de24f69dfce214fa8c3703272d7ef11e8c408ea9d58bae202;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8df3aaebdd25505a36f67d6aac8f27a1bdfaed0e979f35d4fa9e70cda0f12bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75826104e2a6165babb648a63e1da638dd43b2f85cc5e43c138dd32388e0a373;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6af2e0caf85ca0d355fc81526a989556c7d96434ca79c440db8f711179a8361;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3059dc7199e636ad46ef7474f12794a410fa33f5d817980c9b1ea376d6cd025;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78f1c9fe24ffed4e283d8697eb5ee0c91bf56ba1dc05db65b341f1257bde1c57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe68c3e2e7d77afe5817114423b48fc58fc7eb9a4644b0a1a05ca5528430cc64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56c3218129a32bf0c8e1015c2f74992c08fd60947277c2399324a8d1a6fef8c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43f2e098f47d4f4ae19428593e34ff41d4ab495a83688b5116beec29150e4a56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2bbbb612d1ec0b1973b99a35396ecee254c3852a875fa5d51be5558902c70ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h464a2b668ea27d5c1174684b44392af5a6b329da238b348afea74d2db3c807c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc07e29b30ce6a65ba540c8a4572975ef85076c0396f0ad0fdce92e5f2f18defb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea7c54230566b73d47348a2ab253abaa8b6776a9296dfc41fb3eeddc1f2e990a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96972e0ab58c00fc6ede51c3f46bbb1cde42ad38560a0cd00361ef87aaeffe2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94f5ab9e7d2edb0ca9876a105aafd2fa985129606f2dd2d50593f408301b8d74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he42aaf0736e9d4173a3ef2c9f8592a23c46d9d2a176fc578972ce2776bb43dcf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fe4dfdf467ce4f7ec4790c1022136a133ec01e092c380bfc2c8b6bde6b19a19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d78f542e55cad159eb1e1060349f1381851249fb8c88712bda02bca5fafc90c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha024151f4ccebe3db1849661f7edcc9e65d15c335d700585e7370cc547df55a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14fa2a69f09df18a7e14ab0900e47ddd93887280b38d916d1aef4f3c5cf17c85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6f0143d341fed1c05bc34c660bc17b5b3f2255ca6e2928d2d7fd95a56c6f282;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5bb9495172fb664b81904ee2939d1d8a42dbfa8eee59e0abd8966d83112b80c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c1b5434a73bbdeff57758016c836a833a419b29a77d7e3a9e6e050c9d5c9079;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d0d16060976db351d140812d6ff5a4cd4858fd489d0119869af556b083ca996;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15f39e0701a8c2eb10dbecb86148db285c6fdc61211178052d9f331345bd9373;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f822dbb908baa56d45a930cb67069f7d3405d050e89c9d54f0312f2d7711f4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h907e7a34f72cb9dd06af9345319e8fd85d80c236071f08dc46db7805fec6de4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc11a637c99b7fd69993c645674402c9635701ddf5c725c39aa4f6e42e352f663;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ff4973905728a2f7453c645c86d19c67c37cf5fa3b64d022f1597337456e65b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37e7775513bddeb86ab0edeaeedf36332908348e48864ae57ed049c3ae26f30b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8f238fa79d185eec1aa148807883d42a744571d594d4722a444553f380f6dcc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4dd6d8192c5f4cd8903551a0be2602e8abf806f4fcaef56f92c777a9d16b65c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c0620d1b2685368abdc51a5cf71077037f19af9afd90dcf0da5fd5bc69b7d24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84b9dadde908b1960ed6c0e34f7355d9d547ed7988b84e334b9590ded43a2dad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha01e5be3ecd3cfa57be8476fd4316f15bca87656179eaf3518251f847f3ed917;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h704d8cf4d048ad6c97a729bd9c5c9ddd39548be280b267bc8d55094bf3fcf019;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5dbfa56d300abae6d61b415ad06afa5cacdd97582f24b19e998acb5cfb1fccd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h450ba2f733f6d8d76403a6fb462c2c579a16f416253d6251376cb1e56454e768;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6492eee3804d70c2c67f9ea7330be2ec2b207876f38be15501c9e349fd1e7054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54416b733f93a6032a291f998e1199ca21f88d128f5d0be02291ded193157726;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f0608ab6b16fa0d34609794213d9772812bdc28d9005ec39535b0ea824f06e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f9ad694fa61a74c9c59dd6dc769455ba225bb0dce7d5b8d0d3464b0043e680f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21ee6fc4538d99fbc8cd91e36f694db2a1742c31d184b153ff143bac7f7caf6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2445502d618dc84e336385a4db80dc0a580490648be538928ea4f4fe9bb193d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf15b054b3e354cdfd2d20748211057d08daa0c260c09d11c4b8c22877a3383da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c64f55db30e165e6494abb2d080af420db9ee90ab13af6a6658e246099fc038;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd91ba49dc80f43a7844e75d9193be1637742d6da6c838c00d91b10d2972d9b76;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he87bf4b2c2713a821589fe2246863525606dba9bcc0cf9378104c5bad003c2e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e5f2ff9ca1f9f87ac701eb67aeed44b901d593fb54e2e7e41974a2ff09080d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7434da94f33fb6a014e5724ff6a17aa47c344cc64ea1b8f9b19c84a732728525;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53d3e23e4c482defaf3123e599433908c01c2f8f92bd46eb6d9556d7d075ff45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c2f42f9497603446a8b33384cdf029638056a0d358739039a19c6e6c9334e68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37686122064a2cd0a1d5aa19a49d476047170b3046d64bc0960abe9029a142a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b7c0bd053cd9a6921f1c9a568255bb7195fcc9a08f6d1a2d57d5bc402ac090a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71b963772b3aedcbc1a0916bd5d426c714914769a33230374351316fde80abbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79447d707dca058492e6a17eb343ad47cb27e14aa0a96f149b6006489f233dcc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e246ae1e03804d7497e848a1a58311b189afe00b8b4ac22b299dfccd0424780;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28aa15c963530bfdcce71d564bb2dc121af2353156b69dd61e9b232e97398541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefae48359baa2feee49b9ea0f5ccb435a67a441cc52a435b0832f249d614d8bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c90060c489a239952948ed6996676f13477f3533bf0d81624e726ca7764fff6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h343008112b20a6fd7eee5903ef70f07b4d468958f5fd70039bc7bc87148ec654;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70809653c0cf82f05d5a7c02eaa34c7c1422991768612f72eca7c512ca93b51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7dd92a918a70d7d629a1d002da4e7f0dd541b2c6dadf647eaf52122594b84ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he84afb4bf350dbfeb3bcdf577d37aa060a7e1d827675444371e2a65611307053;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e68f06c78125a5fd327300d09e9cee920d619c73859b54d4a055d5e15b21dee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6222ecf2d71ccdfe2efcae571c763dfb7f022741f94f4523383eab8859ff828;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8d27f0ce80c92fee9fac93d3e8770e8cb95e9fa3093a0fbaac1305cab364730;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b15f29f7c12d2007cae68d00d5b7ebc9b50f4446bf67590394e283b137c8b0f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca553a03b83db9967a037981f609a06b3984006b606cd5dc4aec68a5487aa559;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfc56cf8ba60805a10dd2f8cf3169f35ee79e6b768265a74cd602f53c0098d08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he309b5066b8cb226e359c6ce44c1bd5525fcfad283b301b3c71f640277c5401;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeaa2f2b2d7e039dad99900736b6cfece3afd3551568b6cb2eccb0e3bf8f93af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h105c0c9bec0c200a8c295fff26c077448958788767ca28785b5538f0a593a33c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6a33bef939c55506ed138348814138807f6d90315fed5ed35ffa3fd4c91b97b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4685e751da3fc83365fa74650e9da3f10a6125e922b12469d781b4566ee5ba07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7101b5878f3ed68e70aed20d23eb50bd404a387b908a13400d8eb3ae8ef33ffc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23269f744f282649d15c7ca7e1ea782acc0628df055722cad44a9a81f6c960ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7a91e9ab2e6912bbbc3771fb7393cbd07fbfb37b5c9a304346153459744bb02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef698cb696de397db40d68955c2b73fcaa3fdde31150c35b68e0b0600c779c10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49e3e63e2d6467a27eaaf10019f23a31c331ec947693d5de51e7d898b4429fe7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7effb8c315dc533ec83d5c66ce8b5e7f82073b19c1d23bc3ed9d6dbda148e6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2cf8c8b6f2db18fcdc892ddc5fc619338a12b7e9d3566b28fa1b7ed5ec0dc6ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35aef5edd26fa2cda39dc5683071f1661009ddd2f2103106ef7973dc7dedfdea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51ae740f0a90241149da707431cae58405fd5c893217395ff2b8d6a50d078b4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h964c007112c8f281b752ba0d6cf58bf3b6dd28dd5dac7d836d4465e2f58814a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61f37ad5ce389d760b6bcba49850e0c0896704dad0f1992e7b6a9eb2f7fad26a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc78f209d8201fdccb422a75c31c2a8f809a3d85b755c7f1da6d97824de78a33b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b3896b5deff9160c373113e919e684c89f819ac59d3eadc5538abc147b379f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ad70b52f00cd903834b2931c419b3c3030c6a316cde63e9ab7da748ff406626;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80f1e3afbb78e141652fa24f27eb9feb7a7e1039624c18034c95393c90394e03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd967d7616bc3be399898a5b1779710c47060bc89002202dd730bd5fdc624ce80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h278fbaab8d7f1cf39ec136ddc5fda7941227e047782e8514a83d716eb8a98a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbf9df0f0f392b521e0ab66d8ad616508441045afcfcbca64d9f1cff5ec8ae5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h539ca2bf998c10aeae47bf3f07afe93264605ad691d446eeecca75e2ea7b94a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83b4869619ae78dc5c33a948b75d44e974839ceb79d815d9fd02c25f08580af9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8d8072cd285b6f7dc3e51584eda1212cb632e4dd6a71dbe69f8b20d130d40f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa4f90ac176a960a3380bb07793340bfe331a153cea4870bd7f5151fc94a8704;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0a5551e78c6e7ce09cabefe2e6188af5dc081b92499b0a86365e11128e5a092;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf44a9326176f5407dc0cb061b445f605649419cf01f3f0959ffefcc76f36ee60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h662654ae603d9b8ca3508f9bc923d4c811795a2a5ec009ede41ea31819cbe59e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c7436c11f968c0fd8d99487cdd16c032dac0a1f2a54ee4ed9a6a963dd75eaa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf09c2add8bd0494ec452acaec5d010fdb600a5cbde4950f26fcaec36cebaa839;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha079920bd10bcc533effab210696146af1812c40aeede06b3096ce6ecf277b41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdedd1a74e8ac1e962fa11d0c0e07da87e7687ca0117691c894997728cabf09b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h427fbeb1772b9c2d1a04b932cd5f0a6f164bc06bf50a4b0bf298ad039ad12f90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1df944527dc3b962110c03f2f0f0db8e4847c34327183cc0b081257e2af7424b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb82af4976ff5cbc8c94d8331517e7f175d16db3fc2fd1b65acef97546c784134;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24252e8c474f6ad0616b2d55b43d23608bed7171e27bfcc4df0e9a70a8f91b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd33c9d420e061ca0933b039351afcd592faf49ef50f0ed7e66fd9d0c99200b25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd33fc332dd3f3c5efb5e4a94800edb2e60653c3094a665774885430c0e31f0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29014cacf423e2d039e424d85d6dddc0e7259a87a3e7d77a685e2f0ced0536d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e9ac818a3553920926d384e5029d77bee793cab6b3709b6d932fd782d66b27b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac26fa88b9b6b4661220a9312ecec00aceea634fb1b9268952121e7b70e531d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fe2b11098f48b188e59c92025b71a7e974152760fe5fe9e106ebe4f22a50dcb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62a492fed6ca1893cee67611bafdc9853ad07335fe8f362b03f20942524559ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27e6100abe6fa1fbb322962fe5903aa7d66775d1da96316b394f27bcec0b8433;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88ce9d28a3a35e7b2cf806489d1304509c6b8827cfc63612fa3f1a44f3be7a5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58d7a214cb79bae2df94ea37c7b45fb3c23fbf9c04c9919b125b041cfeef6006;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb551b843e28f7d29eba7c1523449eea0949b72f717dbf83e4578c8a83fd64d24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf091f577b23246a6dcaefff2786f81bdc6ddb8369747572c2d4949f185ef8e08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h940a742449838d555814f3f80dc6b9d2f2c8e3266ef2dabf48781f75ddd08de2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0e1ffeef2a313cc7da2229ac1e433e7799e80c921887406bcfb9685d0197c8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbeb731af1c07029485b6824c1409bd5b14f2a412d048256bc15d2cebea109e50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e59985b88565dc1a5898132446369cf94334721ef9ef7c365ceaeb7af134ef4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c74f210f6651fefa410ba5de5cddfb45e98943429c3b5f83664e594531f7ff2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cc9fb238d5e41d701bd0cd118018516300f78b5a49fed99e2ca933b548185ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9180607385442ebb0736d0ea647302bd07de6e91d2ef11c7e1a814c9db99e76a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4718637916a8b0b357fe4edfecfc88d9808d0883d26c6e57d92f34f5c7d0c70a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h130d2d6c037ad96b06d77a6cd4f6c8555cb25d29b1718d8201054ff6f94f3275;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69e73a8dfc9add274c49e6f2391ba0ca6cc924476479e003359bc7b3dde4aca0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dfd43dc01e5684d26c3b7de30076baf7b597a6426b25f37949b04478ee29b14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h824e9c03a891e07c1a5e74583cedc403f836cbad6140de6dbff560e218457af6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha27c3a76bc99104821baa31fdf51c82e4f14144cf3d55b212f5d956c4b96b7ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36d4561dc3be1f8a5d49ff9ba26ebaedc34e838788defb5fe75483c98aaf9139;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3175d740ec4226fb2077d1cd8b67035b5622f4af7271ef87822b054333d2a3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf48f31c4060cba1abedad588383be85579240045b9c7499d727236534c0c92b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7ba5978986f9bfb62581b143c2cf42248587eb77126f3387164c647846fbf71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc603eb6a5c648c937ab1aa9e1f955aa10597ebb670de330351f8555d8eb3947e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc755e4456de6330a88e6b1868b26ca05b915acce77997b8370430ad69003169a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3957b1ade86d13cdbeef1e1ee669fcca99b404ba6916f7aa6e67537be397bfb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ed6e1f25badcd37ac87b4562b73dfe0ff36eec8f367c8f63d2440f360ca10b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6920036cf7a3e58965781c16eb64efa60e78f9c185fb87824d9ecf2508e9692b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5599c188a271ed73d739e7aaca88f51c58835a0fec0deac07182e771c3821e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c5014dbcbfbbfc044c7ee39cfcc092e1e95d28f68d6fec0bfacedde617f265b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcda0808dfff74c7ca42bed7649b937d102c120c66a0769940e709eafe0bbe9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h874e873096c1e24af8ddebedaedb1e5875c5cbe07584620f7c65a3a58977abe3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb350f2881c93e578dc9468acd1ac9e03c96bcdb8d1c36a0cdfcf4f3d2c1d7a9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67dc02be512b3806d738495cfbd2f90127b31ba64dc73bb620554890001c49df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6295fbe07973c6a6141e55fb9f84cb94a31db55ce5ba1dcb5e954049925dac60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf664bd16eb6c9f9a80e0b79e823ce8a95fc76fce6d8f384924ec96baf1dd4b38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha931537acb1fe89b85dc97f423f87e4cd99bd9ba2e055466ad2f8e09482a72db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f6aaa0cc5342e673cf42effc86241207e96a9a69ac3f6b411bfd0fe27d4bca5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha93081153fbfcb5b6aedf5287875e194d0612fb620528cff2832bc9317821553;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf8e210c4efcce7d4d6d2f1bf219144ff20388bd2ab0e7ee66242a3a727fda7e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7da126992bfe536e6a5c97d1251f6aaef5f16eeeb835e1e7d1c765ae2029fd4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7284f570a75614c68177165c94c3f730d6909ff11563dc6a85b2a79d9daeb626;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h797e232071f31e7810422281b16039bbd0eb08891e7756f984060e62979b3878;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h342ab6f257607f92af2d74aaeb0f7fc3e04d1eb2338bcabc323fda3ea75594f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f7d1789ad870f8a4a7d9038bcef8840413f7aca526734421d7d2206cd364c5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hadb5e5389b99ce7f1f9ce9c8d4cd9b93a820bd10544b10d3f1ab0546fa073873;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h423f68a3accfb245f4227ed9a026587ca8647297257ba9f393e84b0dcf080e2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8b1e13fb6d77b74c1ef63f7e48fafeb29dad6a2b887080fc82ebef6b3032c63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a29dae483ab75664544a31061266d22cfd5d8368fb0192fdd70aabe83c86d5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8074c46cd2a694a9b0a786fa15337dce90bff49b57a133294346993451090cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h978ffaa75b513cce4ae79af89e22e50f0e027cf08d2375fc8648b0a2bb74418c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fdffa1f411519823962699f52e1502efd1954ac4bd3167cb2681f3d151d84eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h601ec8f265392dd5f701e7ae07f1452eb194ae6e252984ece1e69c95e63c9f92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78a939544787b3bb087fa51db32d4f210ae8e7c334f81d679796c637e706ff78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31e0610f019f578900d63b2e92606ef45aea3841bc19adec1b505e7b617e14b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd43eb86e177ce176a86ec1a86c54eb01cc6dc7b2020041c762c09badecd1f4a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1504a3c93151550c6b00dcfbe5a69cceb67bcd428e98f6a72d9faf5814b039d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ca8339cdb8bb2a9d2aa975292ab7bf1f91f4f3ab71d5115c66c0bcf5a6c0477;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b219587da4f1ed6535e3159986ba59d77ec17bb74e4f13366b5c6f2867e3a3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59a7acc040b2ce8f840947771dfa8fdeb17ae3610421781f5fde82e3754c6138;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3acb0dd60cb65030b06d45e787c3cb3826da7ac098a4aec234c921ca02a6f28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae44958a6e907825970c9f3b3941783c893629707f12fec17936b7fd633d4098;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74d9e00f5ad657293d5ac71e74337afced12da7f3db0fe45972aa949d61af098;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74b3c56f32204030822be97514b2bbd70004aab5bd2930e456d9f949a72bbe3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce550afa87b1a1715f89c8dac1fe93585c24d2cc7cf5a59218cce91a7b21456b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb02d621cd335fcfafe795cb5c0604d72010295713d2286721ceff61b4459a890;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12669f756ed259d40c9468a4cafc09f6fe07d9cdef6672bdbf64034648a2610a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbce3d414498d1375c2bd411056658c6166ac46bb6617ccd752016f819bbddb4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58e920de10b1323ea2e4a3664fa37bc99e63c392f90775bbc51444b7cf140b19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hace21ca27f8836806db0ace1543aa7dd7471181114d4fe51c83c38a8db75855f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cd46f79fa3839918678dc6fafd12243db01d7d7e8760f87b15cabd3a1621a73;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7f6d01f5cbe4f78d11ba9eb8cddc7b2f62c4108a72f895c0031ce374e603f9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fa4de83451b4e052b1c715b952d4c68f57a5c9eb8bfdf2d7af739e34e71b481;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43bc13fdd9c6b76f7abe90bf673f556f29ef28333da31de770936ea7ee502084;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdef96e6590e737708037893a3f5de6ed2480c3f7dd211d46ce4d0c7e42feb44d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62716b94067d5a268565a008d4ff640f8977f1e60eeb2a0b221df3a0666bc9ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc5fe32669c73e39748d71f3afe1a066d353f12d762d4e61835acbb0551a1d9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha393359dcfb117b379bf493320c896667c159f5d0613b168bc61cdcef0231452;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97ed9120427f8f75429bcbce3d1270d1c46c2723555fce4acc02146af9a2b131;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47628431d99702cea77783a05b65a8d34d5a39b351d921e161aea6261ea66842;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ae6b6029d09a708ff5a27692abc16b22ecef9d9019b52225987b63b84e40387;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10182b6e4a86a140d398647a9c0df5b8fec0446ec1d5a765d5bb8f52ea038aba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd15ed60a93b48ae0db7deeeb577da6632bf6c334ec2c7c4a9cb0aeb4b130924;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd31f9679ad076b58a8e75542dd03e73a0c9c7c380b99ea5b5153ccc3a8f97dfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd2a163d3804966267146a5779285fe45d1e817ccaac9db8b608dfabda32627e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9e89143e8ff161c67e78d404708505e7904bd132b7b876fe7c8eb8ed5926342;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80e0c88bdf2b293b7a06c1960db335577e395302ff23d31e935906e78a574a6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ae976080b5863efe4fec36ddb1c97a28be7a5efcb31dd949d7da8f33096a1e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h858ae10e13a91059f769386565bbf51d4ea678aa37482aa742034f22884efd1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e547e4c25f61b84aaa1a23089f22b8a5d586cf2f27be1036acc62c119a598da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96b22e2825dd4a24dd516dfa98410e601f834e5683672d9f1b875e13de81587e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he33da421967854a9436176dad874add182e7f558b7d500120418f407d52faa93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37cea5da2b9603330855697cd8352bf4e08a8a348d0ca30f6c21c3ee2fc95134;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda1ac740c0245d7930164313e9fc49f6eac9adcfdd8e2132ab23f39210f56f50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h569cb4879729244d4c58c9663034e2f3a62d423395779e6fcb03b09abb0e7bf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2bea07cc71d34141c787cb2af401c1a5320e5fbc41190b96b6d63cf5358fe8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e073ed8ba1687aa37046556cbed89d3567b75d533511d68beaad638ae4597e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa1181b7ed9117ee4bcb976a624431dab5999c9f94a76adfecae0d3dfc286dce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5e668973473ef91c786bd27c187a97ad249ca5fb4d64314f1ef3518ac3d8429;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5abab4e391c39d653f2ebb0a7de20f8604e7c001bce3d091b2df935e25a262d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e712d39bf17d54e92812212ff802b5405556cc3a79415a2eae72ceaab529287;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdfb09fcea6c91438cef9901f220073d3a91521d2fda47c95a1c7f3cb4c18f46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1d5e401af870dcb3d9fa563a68bbfc7aa4aae5d6932f1607dec5633ac9ec668;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd488750a20906dfd54aabf5a693e33bb516595715c6bc185cda631c57436ceb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc57af05738a87b3951a9d0c0c4577ec912a997f7bb46e1ed8a134157a84c81db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f5d5924f4b40ac3af78a3ad9365c682e29b577f279f7bf792431d715d7c68f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha60dfb34090f116492c5192e0e0f114c483caddb64dec2a91c57cf4e01633467;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41d581b3c12debf80429b98f0b4ab1802497b6e0f6e1dc887d07a1d2bf2cd0b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5716e6d455e1a82647dd3fd7f65cec0fdc543637c484dcdc35a266ef9e252733;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b3e5efec301506edacd0966984715a43dba34b5792802f32f11a51ea631f11e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h278b397002af8397ce649104ca35b45607af12c2a8d78d88d73ebb9603a72c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc66b150bedcd361971fec22d36a3a512d21bb5e841157730d7a5c28458ff1faa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h724d2de313381c54bd69eef7b874b973c3cb92b7bd3f5df8738bc387e8465f30;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h554f10f873d3935cdef9ae36a29ed1786aa2668f2deae91c3b4ac2f6fe6da42d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58a4f47d06d3719da31b221a728cfe851fd1d1ed06a1653df53635cb39fdff2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab9733593591c6aab6e45c93cf64019ebb97fd144e71ccf1aaf6a0b03ad62fd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda56be2f78216f8179d6e6a44c93051887c8fb58b5bd8dc5434c39e8dc49738f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e34f2b55d69a9f37a08dfad8b285626ee78787768053c4517f79183494e75c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a0a1c8d86168db4595b11f23ccb400a98a4f8c6a79f294b4f0e6399788e730f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc951a386f88e9f1230383c8f0de63b7fb66a8e731faea848cacb5f835417368d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a4fbf76d9f17819481f2cd345cba0524d7f1713430e1db389bac19927deff18;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd52519c96471ba2e665c27658f1bb5e7ab5f257a1c21fd096a8e9d7b8788ce00;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37f7828161e60ef305da98f430c6978ef80a1555df43e45067430943ca45f356;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbec548294a8676f89474f2ab2faf5b2b24b1f4fa5e8cafc0a1c003e00278ef3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9eada8c5ba048e650a207299b7b7dc5d2893c404d5f5698d82f7f0746f5f5783;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19bf7fab310f59ae01bafdd266405078ce7adf03de66baffbb982aab629a6f3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6c553264f7ede62737a3f45f35f6eef493cd7285d158298cdb86b0be77412ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf728816568523a8d394c53f17f40c9fcf5b777bf15aff20dd9bc61cac7421ce0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1272f5fd88be70c7389a15dda9b87e5ea9931b595f794d7de3af4528e3b97f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e436dfd7d71c77d2629fc9db3c1e095c00fc9195ca06902aa414926fbf5dc9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83f1125b98492c6912b30ac8638a0b76253e9f1c02b62404bf1c5f9ebd67224b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha486ecf3e949016e1b7fc29f8d48d821d6fd6f1d95137cc8b2d7b429bc6c2584;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f3598b92f51be0a84a51e34d20d891e9b42c5be87ac1d51c30ab1240995097d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha775f3cb9f17037161829cc9399be6c8bd21d4f667d22d274ab0e5b45e81ad83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcac9b2251e77e38e06558aa9e9e569c217b2009125e0835c5292eb6982da5dbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3b9ac38dd1783d521a2addb60e2152cb24853999f8d9fb0e39a5d6fced1ad04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb18fa7fab6fe67cece41d6c317e9db54dede407183a0b098bfa912be7013e196;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa916367d9f4fb6efce42b06627596e2fa4095d31d313862505cd2fd15dfb1bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h854f95ac7baf3ec9e431615bff77d6f643e59dd346f76bddfe65e73d9b1af548;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e4759af185bd79d2941292529b3d794be499d1e4ae1cf25e998635ace025579;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8920a84fdfd3681250e40dacd94fac87d44246621884dfeb096bc0ba723da0e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1209b176174d6cf0f4ce6dcbbc2cf77002e8cda6a1cb9f74b211defa86b2e51e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bc51021d460ef1cc72a7587af8a73d949ce9c1589e22b05c2c18b9c3e94a5d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6e08a6756506f6d269e783e791ae401501e4526b358a9542c2f5e99c5504d90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h686625d81e435c1f6c894b439afbc71ad4d64a667223daeb6c1bd19c87319f7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a07e44497aaa5d8220f74b6cf0997d942f3c10c6d3f2230848eaae6b2104ca5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30a44468ff068ed707b63e82f24caea62dc017244dda4c2d5148e36f0ee0ec0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9a7e496c796e4905b16373b64107ac6f03e3047be49a1191d9fac75b05db91b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5fcb5356624860b673de1570357e75d9e0c190220342dd51c9466ade9e5fcbbe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdae76583480789703ab68b68f53c9fcb90062a1bc0b141f206c21f6e080cbdb3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5270dfd16b29f46523334edf33805e6e254c9a16934eab2a769814ff34d7fef2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb74639750e3d6fd0d74dd1e1bd217efd637f0295f285a6b46e36ea8d6f7b058;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7473bc7dddaea8ec70088b7ee900c13766f7c996f49ad6102e82b5c240bf1b8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa08f1a1439d0f16062c5e8416ddf87896ec79d049cfe7243216c5de02fb0678;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9c3a1fc503514a36835d0760a8087b8dea2f9bbbb30065ba880db2dbe440b7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha552331bb709b34a7dff33dfe4b5d6c82169e5c0f67f7f0e24db6c82e2e6f26b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3209d2436c07decd8ec19c95032db89abdff8f38628289b92268a3968400cd0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he04e620af6bf7d1981725bd7629855a4f8ec53a39394a565e65ad07c38271fd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5289c7c8faa71480dd7132db4ede13bba48d3a03201dfd0950fc187823b6b5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5749c8bafd0e19e3922064fcfd000f9636ee8c55e68dc7d01d280766d757d9b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2eb0ec51f60d3a7b89ba17897e7576856253f2a0c6428c3d6a9ca4c65b6c68c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h939b965debf5b9cc61dae362cb309e65d11fd14585f263065380243b01b39393;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51e226c16743b5bfaa984d307bc7b489feae289b7807e2c2c0fee94225bdaa4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23076e593b9f78af70e9070432782dd732e013307a1445e3999c69385665d46a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea62082b30096a7301cab949f9387df4003abb33398f77a7b243d76e98b36ec3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf117139fbc3a01029ffe9d380880116766341fa03505540a3c9da467e8ada275;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4b648763938b00a044530d7bb154adf2aee3cde4800fad0fc222ab59900897b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1837ba88eed663be15e51829ce118b50a4915145b88398f4b7e4a8454224dbb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd272854031389055669642b95b150e0f7c80aed805281c497dcb247029d27515;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he725ce23b9e1a9fd9ac4bfd2a90c1d0ae2c862a239a99dddd0581059e818a736;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11548b457d9e75374e1f1d894e03db910b57e96fdc4991bd40f397f61a5c4167;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba7286e575b27c6bcc4a491f37d70b7652195cb6b050542f9992a0b2d3db19bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h278eed41a4616e457be9272223e4750577a69f69c53971af7cc0b9b6fd3cee69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3360ebc09ccc8eb3d70b68eb7c4a2cd35185a91f2ed8f986b70255fffb9850a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64527fee96f67c6eaa7f6e1a29dc29238c1a3f326b1b75cd7cb004201a27c0ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff0901aff494a04d287787e3b8caaf928bed07ced62c674abb138dd3f5ee207a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25c069d0db9467a10e194043793f6004c136e4786aa0f3bf82fd4c01a08b8776;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdac6ca8901f38b4c6b3471798bbc75abc11be63fa0a96bd8b3fd347a519fe564;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h313f02bdd509289d11c3aad5c7219f3a02e56aa3fe34c7656841b2e84443cd58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f540e49ff23fa8cd31fbddda3092e7dee91704abef72db6850a4368d15cfd46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf3e76b527939e6af2716b721d71b2b8ca9965c57dd6d780dd323af511cc792f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2891dd0017319da21c639eb4baab3276f6bd098de79c1634cbc35ab63d368443;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b720d62c0e66ac421f0c37ec7ddeaed39617c7c100a87f75b3f153645b80229;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55b2907cd7af29e83956f2e4d50767bba22892ca068c9942b49e1989602e157a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9dcfae68d5077fd23ef486383ae61d262c6c0a40b36e281ec8da338ae8df82d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d2a0ed4b262372acfbc9b3f37a5d6c938ca768eac31c27200acb7f66eb0230b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h456306043f4a4393acbbe693b53e95c71ca2a4b43deb86a2892ff2c2dcbdf0c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd016e89a255761b69310d09e52b771b2b639002fbdfb5e925062f0040eafd68d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h924ba34eb76cb629eb34ab0900735a9b0cd72673dce79bc748f472225209a271;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7143f025d59067be0d0f9ab73492dd8f96a3e590d33b5a23a69b0bf846e1e60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha562abd31c9e36195fa59791c7afa85df5a95911230bdfb92e25f421faa8d164;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64fdec881af184f44227e73fa8f17e5a1b1b41cc0b9518a71f89ae0ab499558a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3aa2fd2002d850f16a16daa025b8626fa39327b07aa499d194f05d3afa4674d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ee86009f942a5963cf3f2e4c2ca93bb43d9e0efdbd1a3175a345f5d4b7bccfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87a2d64a506b9daac3dfe6aa4069d99edebe528b72acdc62dde033c5763e400a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68ff36e1a84ce50b9b584ee85c7661fe329b2f1ba6a2a14510be313f609468ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce3607018d09be1d24adc94790c3719d975073de03c206d5bb082c1537baf3d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1f018d54a968acc5f8de0adfd7766e37e53b08769fb4f4723a799219c6e26a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a90ead41f1b9d2f4d5422bb4281aa3afb06c738b4e74a51f633d574c50f4569;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4b349d04e72f7b6bea523e7347625f837894e1a7db47e4fc87e0dc291fab37c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89ed089b7b232bb4791bb6598d6f4da2c6cb73e3d1739679c70f71822902eeea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9738b533513c8ce1f5867131ea5f839cecb2d5140268f1637916b4ef453730c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2bab261ace202462838b6b5633f47c8c1cfff8e923797484e1b7478167a3a20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd7fd05d3a472ccf71571ae0e6d7c9d8282c4aaf6e22c8c4d85801e5193d7c56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b2bbaa19f87d0a158098efa675f5915d4effa0b00155ea38d8337da5633d567;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ae2b7664fd0ea9e1c2a44cc747966bf48ddcadec19f54316579e1e529d7f516;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a51cadad48caabd4ffc79e5fe56febfb15ac8c81a467589af603aad7a4e6740;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd667a3477db82f4282248d8e32ab494bb842b3905ff246b70598cefc77a98f10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h165aff9fdffcebb67ad5756d90ef95a986e21bb816c40fdd6bd2989cb8d18c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddd13cf6c92451ad663d54656224de18daaf4744e30f3692a0c8bc1b315d45f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf21cdf42dd631a483a925e948779eecb2d51dad1ae23e296c4e6894bbb639da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31f31f50e979325dbab4913427aa5d161724239f2a36ec185ebb4d351a2f9f7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72da4fd32d722655b604811068e374a35a2e02660f5d069cfe8b7e756a608a6d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48919f3a4df7d489acfd0c35e3fb8661d03ca9f21d184ec684cfbab15877b131;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafda1c3eccae58ec2ed07bb506fc81ddfc8b177dabeb456b871290a3de34a07b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d40dcdec0c1b71ca4e5f2f99879f4552eb0f8930bb25835d2b2d66af2a479b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60217d4f59ac70bde0a952a4e8af635f30410764787060be61af28eda5a96b29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40349fc304a808b2737bf40c35f0913d2a29453be3ba99b281814263f470b7c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h680bba06fb749281c067bbad809c2db8867592d86d55b58a5daa374d7ab7f09d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc34257feb298b390b0f224a02be0fc1d9332997eeea82b3a040f523878abb12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b533c36a74c92b7b07a5b8ebf26214ef1694f530bd9d9a0fdc6079c033870d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1db8b4faae00954f929731284053bd568e96a036f6a2593a655b0585cbe968e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a1121221c2dbf6bbf7548c381f2df278e5d34e2f1c9295cb147400746e2042a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde16b7398f87888f8204a93c117739133e2d50be04956de3d68b5aad978f4ca5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77bdf4475fb5379fbfe808884bd114d3c67157d4c6fee131213b0e736c5de51f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h546d8da2797dc7c5ce3a5089ae6c6bdd72d892ed1b881dadef0c3efb8f917336;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he320d620d036f484a1c391df3fd1eee4b9e68dfeb1142b4e37d1b7ea21e70c76;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc71e7e185dd94ec6f94138c747e1c0d32223710893510b10cb3cd2ca9ee28ac7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h660e8101286350cc2b21f67211cdc4cc2334cd9259bbc7d867be8b663f884b06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha069254f578343f93f4bce1806eb05c2a14f06aa4d594835ade9e2df32033a3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd26c465ab24f6a38f3dafce00362694d2c3a767950ad53137eea1e9f437ef8c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0c08721ca2dd9d410ed9e250866542541e4b67897094246d05ecee927ba16a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfab8110a1829b7ac5243e08310dc2cde002ee184c2fcb5d1844de3cac4d770a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3751f7a06d987eca648115714f5739cd12aebbf89e9d315f24d39254edd07fa5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1f67b3e45aae12c7aa912e87a6f790d361ae2a90cbda7518794be13d6cba5d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb43badcd21bc41962b4bdd8aabb88d53f87e4b84dce7db3e76a47f4797e4aa8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd1c3ea372bfb631d84e876ef4cab63cc06846b2cdc41f7ca72969d0766ed793;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h171de172d7432f1f3038f89cc12cb074c689789e253dd8d4386617bd621a6b38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd37ddc7b7b207b63dda74fe661e2043a3eb2458062f9d610deece5ce405abcc0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h897689eb758cd128eb06be69577649d022d8a78aba0b353da8a25a931f503e19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h858d4610ee96892a61848a87b0ec964422f7fcdf08417362a3807df60cbbaa36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9366414513490fc78c064dfcc3749842a6ab6539aad70af5e39944fddc478ecb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f630b2afc23238973a1250834f3df42e692604f61018d2b0882969db8d697aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf21eecf8e483543b0625943ddf812920dd6c7537bfcbf07983fb8f2b5d7b818f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd40908cd9d23bd82b77a953e939d285cee31d1809912de060a8582339a602aca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42e3bb67c66f86e9beb12cc7792c4f3ae91a2c2e64b19c49f5da3e6dbf304661;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81c22087b7f47f111341cc6a2cf4bcf980af753fdf1e76b2d055547a3b155c8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1eed6b3d0a4d0711ac05d825adb3f8b28c13b985569ad765164b91d47229fe4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdec2e463658a1e9cb784fc559ce6a4844e49a34919d06541ee83ffd64eb7abc9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcddd0f4422241e61757454d0908b256a6ab15dbfd3e1a8f4ad0041ad8574f9a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h714d2a541115fe202e5b3777cbcbf50d94eb9b2c99238052b1588a851f320b5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff4f63f0100b7c4aea28c84356c712c934b424ff393217ac467c651cc9d70652;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6c4fff5f84d10cb3a02b87f6fb2295e958105a97de55e940894776b56626734;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88d93a6b2cbb737fdadda5efc99e9507bfed1543deae23665734a3e359503046;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3dbc13f689b6c30d51e4cac0e267b1c4eb37a596bd50694ad7636d07983849d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b45ab25bf08bcfae7feda7c578839e19e147c6a37ab78092f0e0b9c6d090564;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57709d596c634c7b55a7e4bf84782bbf1fbb86894285dfea8d56cd54c37e3fda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha85502f1019687a040d1f45c2c421adf475c465584335c26dbd3381184467968;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeeed6b455b0bde051ecece95df77d2377e9b958977af94bfc52cd66c0c388d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h430d611bb23171f864400d33cc9db3c6946bf56c253270a70f297cfd3980c45b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd699fc8fb0202517ed6111d6b597de98629a6cf92b0c1439cd5aa2459a4e2b70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb44774fb937b7aa69fe467c3ecfdb5912d05d52852084c78ff0feecd1f2af4ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he02f7f4c1c28f431f4ea209eb0f0d3ddeac1ef2368290416aac9d10c688186df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfffa1afeae344ccd770f9539378a3ccbe8dc5c146930e64552071655cf2277c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd39abdb64617aa570eb1739e5cda506f6f7d603c2770707785b7051d2079703;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12fd4c200ed76f65db1a7477f5f2a73841c75b3c11610a53011cdbf330c0d5b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he81a7374a360c8019fa127b47a1b626bc82cec6a83acd0a211261b0d5772dc32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8070df1d26c44eac1506ab3f04c292ce9bfb365386ad1a5c515606b61b61ac20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a32c13fa4814db26182c36fed844a06d26165999120b80677735e1b20bdfe6d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7232345f0b901e7d2a90a6122beb7d8fd47a94eb3f687cf3fdcfc4ba336960cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9895b144b9cd4f78f26cd49ac5828047d4d7de10d07194737e5689be9de8809b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1327ee9289df7af26bc63b1406a3a50587b60ae76eada243b407cc4e954da160;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89f402edcbb1f55366de45fa7d4a5c317ca59eb8d870ad92d6bafff6750f3cfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1c7e012054271e0248ed4b5f4dbe489dc1a4f122d7cf0623e6ce61ead777f96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf93c5467406ed36aed9367e67ed6a3d5b3f0a23f2d55e13afffa1ae041d8b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e51ce940655f61bd2b5d733359093e3073c24bf008dfb09b238d72fe84abcaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd37d72c6545c36bcd350be4b2b283d9a2999e50438b50cb803587b3c5e1e00ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3bcc86f093eea450c4a346ec114af7ca9da45f5de95b08987c85ccf4e01adab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2bb97200539ef2e7f6a2ca8b0bc325cfac6c06dde37e2d71b7707c633439813;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75977c20177e55a5f17412e8733b399109bf1a898cd7718417cbcbdfe559656b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd35e4a3a94ab6f03c104390822406fbd7eeaf2e2020eba003644d1769e6d2d8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae0395090a49a3516bea59fb6af349f4195fbcef879e5290b1a4be326d5a0c37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9f1c00266e9feaa71ebe16a718c95b63ebd6e33b21a662ade5011ef13cd96e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a759ef01c643e80830298eb293669c6c7daa8dc536be3b360206840451a1ff6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfb9970ac4e58baebc80a010a78792a8ddadf3d79193414542665d6b6ba26862;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c2c97923390440abfcf380af9c2e4a14517bf8c0d948221e560f7017a56953c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6918d34a605a61cf9c56b2a4ec3107468e6f986fb9ec96cbceaa34b25bbdffdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he13e07b889c00f158e30eb437c0d99b28ff24e24b9e10bd7c2851ef9abdbf00d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9107a1f5f3c5e85ec1a12446755c710f8af2493000cce7733813fbe6dbd72c31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dd31b296fa44de5dee5c743ffc457c7ffbab75bffd6c213b48116dadf74bebc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habd8747b4fdd64d5107d7cb71db46ab275b93462df2b64767932232e518600c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b0cca811e4d5dd7ad9e65196214bec9df06906f53575ca38bf0bf9b7ed4cb13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8d50ff4c6be2f5864f5d7380e9c9a05b84a6173876c9e44b0b513229ec4e600;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffd7e7a794d5a98e2c0062dee7897256a61c13472f9b2b4a408ab63960ddcd68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h570419a50875ff72b1e8146ec423d2c5ed102732edff2e9fa3d22ddc66b86c2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7658f22f3ba6e344d54ae95b3faf1768db15573ed74f0854a6914b8f0ca27bc8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4922682c66a6ab5425d4a9c8446abd8c4984df5867d878669ed7dc72fc28e074;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef72a140aa8656d7d4edfbd2fd33141d2076004333e50eab4578d577a730e3f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc48567debcee23ddc96641f011203d3d6ce8ac048634d6d1c54ef800c699899f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39344073118a07f88c9183ede59780a141ff53dc264125bfbec7a813c3422c9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he969400ed16f955a70590a8e356d77b355397e003f4bd3df5fc392c0304ec423;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6209961be5637ecdcf58e3b2032348fdd88ecbda5bc4ba409a45c5b9b96645b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c2cdc291b92b24f4332683b670c7473e8dbe96ed56c243b288716f86d307e81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96bd0b7418cc5f16a9fb0d52d00fe2fc7dca8ca6e947a98cf9b7ee17b6a9a436;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5536d01e5cd1558db1faa48d83760d354e08e74577b106002702896e7e891569;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefcf88b7231e621d673e01d138fceaa782a6521fd8aa8371d112b8af0da99ce3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4172b00d6f1b8f25033f63fdb2f47b3cff73842f0365ad9ccb8dd8619680922;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47635db1fe51fb3fb6fbfbe0f8df0c1ff94415450733434570d5c60d6bb7175f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cc97a328b08de5b214220302c06df71494213ae5cc1b12947b2d61363b8f273;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9093e041cba70aed90a7b37a39ced834ea2bc4125f238db7233e74e849ce05d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1d7e31c94e9f0874f7b54abbda05e5334146b21a4e801b5eb7111ff5757ae5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc66ad2ed3ec7212db144c25208bbe2617059bef32e0bf8ab32a544a347ca7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h549e11e12f5679f52d20879e0319fb9a8c0c434fa7123e61a094c21af8d7feac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c1c23316a950804e9a460884400755e7de1b66dbbb601b0809d9b043aaf9b8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h298075444bde0151fe3431dede9527aab0fe44f2f570c5f815620256cf80dc62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd1c589f5c100d563db44fdba260b791e526fd28d456d9556533922130d790c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe36ec9a58b6bae9f5f1607d2419bedd18b3aea1490939023272864b8ec30aea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc738ba78bd380c52d4ab73e6084313a128879a199db92ccc60badd7ff4a59f12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf71ac44f53a267c382a9810d6ecbfd7340f5de33a696c5b62fcc26f82b121cbe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e0df883e4b87742c7cc95aa580f8df57df385324242828812404fd4eb921541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h581da15b4407f407ebb9361d7ea8325ac6d80581db5fb0a32a6a3d4a1a6d40b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he68ff090270008c535a6ddbb7f24951789330a4636b4749655e2026ea271df22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd094b62966ab46c95e2140e30de50dc7d5306ecbd551d509c25d73acbbc34616;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1b854b88689d76970a037bb9a9d68780ea9f66f0fe2160b66f16bbe05efa7bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e5a93bb53b20ab36710c0bf57b17dc7ed9005ea8118d378f897c50fb1ec80ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20bbfe9f58776f89df062c28901f8d8764f051f3a71e0fd68ca4995db864eddb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0d67bb506ebbdf6c3348d49ce111381303a71e99e35eb63fd35c086259c01a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23357516a5e3b98e453dbc249771a36a71b0af676ae0066ad13f0c7e151b750c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a863e0a4642733f0324b16040549d1bf487fb66ad877408c100dec468beee26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfadba2f612d2a68b7b3c4aeacb12561933474fb9247a238df21e6b7b43d1fa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdeedaf4d8d933f0f489fe6323cfa93c03e65c2527c128b7202c4eb262e090e35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec47d0f677f75017bf08e96b83e5325ad66f57fa23747e4cfe24695cd39c242d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8676936ad132c1b1f3767b4ee87da8e4346e65f664e873b32f368b1d35b62c42;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33a3e9de08e45115fec7889f76a1e3afc56ed89bf5918dae5117dd4274cff153;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a952110c51302d5bc0a9b006703e480fa19f8496a6600c9781cfb1939101ded;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h173094b1d2bd431c81b64d9d0fac341bed4c363f1ed018a1f9ef5934d976b7b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he41d905a3cd89e256d118189c3cab6b7d3589b1af414a98f6efac489a3679450;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44245a5ddf9dbfd54a0fc76d77192a56f654f96ddade1edfa59dcdb54dd4d4d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb99a91523f90c79ed576bec454391db1fc7a404a131e37599308c61247e32cd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h206263225834b65d54969dcae8e7ad52e784cc042e6a18f010ec91dc80c9070c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17ed530d6495cef7c1473a64bf35d39dcd28da03166b3bcf9c52c41e2d2dd0f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc8e5e35cd966453006920b768bcaffc2adf17f019b0da4dfc6bb8deafa03dbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd44b0579706b7388e436ce3bf18daf4a0fdda663dc0c2d76c909af0c916825d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5f6bb1517bce42d70708ec27d97c9c7aad588376777affa03df2414ddd6ed77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47a15396ba2a7bca453059a675f83c04b19152b62b0ab6435abb66f9864fc6f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h161d9a637b73a7c17cb48968284fb147434814d0b83dd7ffe2b83d69fcaea716;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d05a955dfee3bd9dd1029415a59baa4bf4e466075e6e6e86b3daf9225fc966a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h703fe3f9e2ee844c8028359c4783be2f2e4328b35ecd45ea6d1f2b78fb742f63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd024812067198815f2c304cebde3adf44988c72ec16417eb00c60048eb322d59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafa37722701dd23ecf1ca39f5532b2d59de2dbe71bcdcbe5664e1e7b5246fa5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he62f963cada21123e92b7bf5384e79e2ad97dbe05a25e287e87f331db55f630;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1eef0261e82f28bdfadbe1e54a0166fda45027d9314c7bb3163d1e6fff9769fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dd578bddc1309f8fd67b4262157d26b0919147a891ada48900dad195bae6217;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bd18f80703b0510716ad7ed4d501cde3fc15269c52ea200f8724df2772ee13d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d74b6e333d68f4f4fdee837d41dbbef6e403f5831e50d9339b01809b1685a8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd98e65eee0fe02329bc70177cb6d81dcb84f8b721435a96184fe47680d0092e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8515334012e1d80aa40586a1efbf416fa107414e398874bc0d4618f018c6f989;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8cd495cb85c58b13bf3a1e8b9fabb7710ca2d768b07f0ebdedf704f67ae85e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefb77cfe01c186199b5080371eaf9bf5f7f4ac5b46455c449ffde488ba44ee03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c6c487cd89565e6e6825f26f53bf6fcc2af60911281efd947132075fbf8219e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he60b8542189d79df3f75618dc5cf4094f9d42c1e564f12693b445527b41f21e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbea4a34bf1ee4ddfdb1dbb27de9d63b3704f30cc313f069f888f9cc3f523394;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63da99e42308ad6d728c55849cce99ccf2ba2bde6bb450992a0c7fd6e2f19446;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab1ad7b699eadc80e3f071b859f99c23a38133c4f1537a830fa534180eb7f1ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae442e1c8ea4cf86beaa83d1d37d21f9598346f1761e4b6157a1c5f9cd97bd1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had326d7fb25c8da732ce603163a4860e94acdb6370d509cdf8b7a8919d239540;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8716dd83a4cbbeedf6f0ac6b02c5cdd8c8442bab1bb598e96c478988ba7e7645;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5931c4d7999b1647162ee6b507279b91162c4834e6ca19664e98f653732ab507;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb22fcffdb73dde48f1d0a94cd09491858ea469e31c32da1b8b13e0a5eaffeb23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h438a77440c42e5e40c4d93d10cc018d665d8298287ced2d44c523d993bae651f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcea9aaca99f44abdb52b2a8ad44f774144348c2e233c1e78375d80635ee94f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he04c1bec39d8e72ada98a6fd44bd4a2d2a77ff24596d737ad417326b4e040b03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66caa48fffca0f5a7ec2812442db8b1112ca1d3aad324ef996de2eb69d7e7b8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9539e7789f2fc34d26c8174aafceaba04a785ccfb6671524e589cd3cae1c3d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha793ec59685a59c2165977598c4c9a1db3cc439493544ea09bc8529b2a0750c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had12ba682acda653b4b39eddaa1c96c2fd6bee79a7907b56d9f95b38b6e1d069;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a63459e6bbb4a2ac2d8538b333e7390669154f2d4e138d816f2e2b87b0528c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5708e595c66033328ba509f79f87d20c8c3e88ea4be80f2efecd07fe21b37527;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h685e5b7c3c34147b7570653ed696f7e1f6d06f38572dbf3ac51a1ec5b50418cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e32a2924fb5db82082f599249447175ffbc2feadc7531dc314bc20fa48faaca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11f4a92e9aa006f98c4b37993d6eb2e7fe3c644d36c890b3e554d1b0faba1a58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80bfa0c83c065cfcf2dff9ffed34a6d58ec811e391a0ded294d555180bf710d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd430996bd5095b6b7b95b9bb96c330f7cead8b070ebed9d9459dde4c18c5dbce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h830dc02b7ca1a1f6ddf0fc0ca38f37d09bbbf98a1cd8d3392b37715423b0e589;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h746195a19301037d46582cc8fc1b1d690e5bb039d9eead2cf1b09044c654f640;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24e266ec68c8d66d235f2d130d7ec17ebfc400f83888a680c83f91b55e5e3202;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h124fabb8f383346adba4b96f9415e7aa4d33f820309637d242b2f9c97b01c760;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7985a13f4712313496b7e1974afcebbdcb357532700b162c355a14ad86ffe15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3964487a6564cc858ddbf8d7e9f6f34828c91ec59418f159158da5ee15b53caa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb74f9a73992d2ac56e0447305383531096bf34771aa14c0f51510a16ffe95ce8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57210ae48235bf076e0a896dba26da96d762b4c25ff382b56fd2b3f387217e4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h404bdee58279760bf794ab4f1e916ccacf840c12422a71b7b4f6f9d4f9429875;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf57ee997dfbb6092b6dd507be33296cb1ea338683c3648283ac1c8b32077a239;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dc21ccbd21c2cf0e751b969056c4f11b05ef09800e9f7ce6648e3114655334f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12c2ba1690fb59d247b5d2f94b1c7ff5686f5ca997b2690ad7625b887c1e2ffc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8978bdd798a4a8ce8a339eba8a61949ae072b9494e6f6e60d224eaab89a228d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1673214757772e945a68a8b8daa62d7c7b09da26d0264b9387b14c7ed34bb49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a0214b1ec28309fbc198941f592144b0839161d08b1b168bf6a8e0f373d642a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3aad0c0dad9f4958ba10de8d4e49c2c507af378c67497caa2dc65ad2001bcf4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha232a370003aef5aaa38c84a800d0cd1c018599f65aabeb725dde1595a6950da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h850bf882fb3cdaca1f78d9a1387f98d75f60a5b4b737e79de273cf2b5b946e16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb86ca827ad1e3885a4128425e3656abc718661985c6f9a17ef3313bc65e1dc01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52bd67cd8baa070bd2368f94f91b3979b51f4a055d5ea23ab9883044520870d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a97d3d2e19f966a95dbea588eb9281919a229c0c2bf16f88b4c0694a78771d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33bbef9f6d03b9986c45b7d616902d059b43dd58420c54574900c68a0c819aae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb5835c9fdea8e68a6e794d718d3d66ef3cac0f372bee075a6fc7b2a07efc531;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58863b5b5593844bc523410d0f9ef4e89b53b3cb40ceabadcd367cee36de1940;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h818869345e02d469e88e0f653c93f18c52f0b428deceee6e455e5919c2ff0e14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a1aefc9211b7aa7cbacdd775315df1efd2c16c7660018aed56c8ac8ef166a6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6bc3a93ff1fe7baa79bad8c22657de3e99f4c8492e710447f6e78c3fdd3a570;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcb88b265f70d49ee547d2e0b4a0ea2934c2c60bc89675337de238c39954b71a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3512dcaaab3e1e39e0594c89c672f1e259734c3b5a69b35716c68444268f2b77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b0af78df38a4b69c438d9e60ee06d478bddb705a0b1396a1b442298a55c9ba9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c244bb2d014ee140f272ed8c8a6a270a97713e1c9faa7a77f22727c60ed4c77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c4b8feeadc224d027934321e2dc9b5cccf13aa4a1267896a945df4a8eb4af7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d393f93aa81508cc8674e4d178f87ead9788e25c8ea6f97caa7a2094f148401;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99322f1bf85bca243dd5b60fe9faf40cd9cf33bf4aa7934d31ffec54abe518bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26cd5cdd308d5c6fe1c318cbf4f8e80914b406b57e49c36739b7d8a5a849c2b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32484627c4cb98a5e120aac62f44a9b08d0e072a8259f0eb2a2dbcbec81c475b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45f3af504e0e155bab0f8ffc71d67d2b3fda867270b5f5685c11a352ec92648a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79839dbafb17f913b9c31894bec17efaf92ad17920e74cc03996465189c0abab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6e7d8d0a8faa3f11dc74dd794c0ada3ad81e850c34e33e280f70b1257a3959a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64d5a27f2b0c48ab94bf2b588817073aa3392c51be022cd5613a03c2d08b697a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8577e5225ea1d7c89ef8f7a11ef069eb02ecbda4ad803f218f72c81800937097;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc3ea6195fd52bc34e6eb21bc52f7df9e77317cf84faf7d6c8997179d7f3a924;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b1370e626eec00547b94bba9245967ef50a7339d697690970eea4a49c74ea79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2bdea4a0cde3fba72782364835a95d6e9c7d79114c22a0f0a644f1d548d29f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8237d49f5f5dafcf750fa9a4e947c52454561da37723de331b9ef71255128240;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h420dc6138da7d7d5d39e75d58cb4dec3a1ff8e9a7ba14fe57b0f3a1e1506a843;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h432107d9a4e281586c6b63029c30735b3c10092f697bca053735cdb8688d7a5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78d2343160c26bb7c94c594fd281ca1066186a74220ff0f53ee016a55a526aa2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h468521b5e5a6fadecd771f1cb7e5c212878c68223129358dc5413467545bca7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5fd4d90314ff7e7620182dd446e3bf431b5d77694527e23f2d7c317ac75adcf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a2fe0dce13849bf8a5157b8f4ccd903e9ec7b27ced6c78ffc13532b42cc545b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he88d3f14c533bde6e7641396a7633f9b6e8b5e67e35c3f93f0bebee19214577f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9f3a3bd9cb8f9752737982d41b8375a90495ccc81a088c0261df8727b30f345;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37d592a5bd94f3a5429189425d66463744190f280827002d513c58f76df90834;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc17426485dd93c456ba8002fdb9996d15425a479fd042c7bb4079400c11db754;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd9f4c3b01eab15d7827306f62f8d7b6098433699731475c773bc0fa831acaa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h183245293b560beba1c8d1d451ef747212eefe2a65a156a94db7485980b82e61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4e6e5b6a045101faa86292c2ae1d688d153409da980b9bef474cfdd9c041f45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6294748a429d4f534a4f4b40c411aab4499b3922c1633f07728ff4f231aa7ba5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heacde76f287f941e883f4905aaf5502a3706484c1dfcbacb93a93de9476cb77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb39373acc1c9fe9c4ab53a6ca3ea0647f5bf457bb2077a7971ae2732569f1d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed81058f7047efed3d35368ba1ad45167e5793c0af15d5e4ad2a0ceae4d0115d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48dcfcdaba98b5ce720006bc249a0ee909a23edd3b5802cd6ea6092b82a1d483;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha83409c81089f84471a51b6647c42ccd5f5d62211ea6b81ceaa7f32ba4b6be40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefc6b92ac16ddfbac023a8075119d338a524cea94b73c4a0c6427f2702a6de99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32a24c21b738937bf56e3924d3f66556a8cf600eae7929475d748677e376b19e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h831b3bb82c249bd93a5f68527d73458d7660e4057a99f0cd771ecc11cca45492;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc728f6b7325c63e60c97da0ba9e33bdd4f141834722016e5879eb57e811279b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ce8055d5394e36722f49989f7ef8f13430c20c0e63816c8b1d623f6094dedd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b5b1f926acb4fd9aa77fd5e507c054f4e6ba3544a740ce1467ded8e028a97e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h985054b6eb81c2f4728181a2d8b33415be0ca9e6afab42f7638c510ad2c81bf8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67b06f7ad3ac33ed44b543a78c9c9d93e9e43cf5ecda1ecee23de3bd3078f562;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8077f419aaf34edd65133c7d0e1614d7761718485ad9f2f78fa75d91b9263bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1719e19b0083f2e0f513e93dcd6ae97b503bdf4c27b9118f4d0afcf531ee13bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72b5a5d14e852801d280c8db1e26a920d2963f68fcb3c2d827a54ce4f4f636f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c59a929820947045fbdbecec4b5246dbf4fa0936ed7bbc9bcb28bba7c0bbe0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b22f9ba40cc3eebfe8617c0917f9381155b778ca037cfb2e10ebde665e96dd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb89f6f42783902c24a6d2c19ac119f4aa571eb5d22add4fa162a7d521946b40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf6ff2f2a631f76ce2eaaffd793594db309f79a240e395603bd2e3c3e1179de5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb06497c3736d0afc2182a7d5fe3a3d7d2b5771ea9a7c72927141ffbd0fecc0d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeb73f7f6f988fd36e8a952419f39e6f2529c457f9d50e902782e2ad20e95103;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fe07125f6afbb865e96ebc9fec2b506ad02fc207d6c499bfcc0202f19498ca1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40924e06a8fd142ec467466e6e9d2a4c9193288c22aa8d6144c6fcbaa75ce3fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9097a91ef5507618c9b4a69705a111d2e1e022c5dc515cb134d6bf84ecae5e97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5877b11ad660b05f6e97abd04ca27626935ce61536ec7d9002b5d4c4e8e25b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b22a2078cc7786eeb4e18fce3767048148d34d7d741c58683bc5a3b2a2c923a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbac93cef327c7060cd629166643c2a30b46caf606eebbf5abc12934592ae9855;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3ead6e4bb36eea69a5f4a50311ee281bbd8c220fe9eb6bf2737eb69420bf91b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf113b964add1cc2179a8d0707035951691d07e39d4a7bed96bada5f11141e6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90f764d94300e690463d6fd8035ea3a1b6c1e936bd4ea0a64479aaefe853a7fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h821da935204da5f37c809608c393648979a2e303f2a2af9054d8c81ab28df80f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h300d7012f7b6350b51927ae13e1688612e0a0efd781482bceeb923233bf6892;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe7ccd11396a56478b9e85231a15c84a5c7a01d05101a0a44d468ef3c15a4fb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h144d61feb3d5c79274f1542f094dff731642dcb5422dbc13c6bdbd20ba3aee6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29c67f3ad1543f020f5d031237112a3eb68ebe959d20cc88d24b0749a2b27d91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h449928c6944ea0f5277954b6d633427a8097436830e9b96b498f55f8e2002357;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a5d4c71ab893aa7b9ed745189d99a599f3d84fe47562df20cdff5ebdab02977;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b248dd2d77349dbefa703ebc060d4696f647b8317c4b62a0ce6c4c60489e008;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4a0f0c4bccb8b87631a12507986933848892a461865decaec093fdf4a8c5614;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46e821d6a7cdb68b6e12f6267e4003676afe8fdb80a86924a391ffda93896541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7386ee1dde199e6702c4dccdbd894c5effbd023ad0981b171fdad44d308c2d3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94d13a39b5a06f8faee27956191f27c3c1fa2b92347443e0ee771354b3079efd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6e86a94a71ba38581b0191dc1a1361fcb84870a6573aabdca5c7d05ab8d7c67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98bbc09ae804c6cd5226efb0f275693d0b612cd542db2609999dc3df40995dcb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd60fa58f6b18c58be38d4e7a32ab639dd3965e245f5425e3db1d7ba53b8efee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce7eef10bc8d5eaa9b34400f3836bd2714637c7e6c41f7d05fb0ec0ce13ffbbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba8fd2c8ac0be89b289b3981036745ca0bf03c04e0e7a8bd33a9e262d1ddbf11;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1024a0f8019d5eb1750a6be48dcf23e73a8b7c5235462c95ec55f03f0e9326c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29e05c8b5014fa79312140b0e0eb38b57721785ee76ba32d65fb017b9a4ac63b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h347b4f26591fbbe0d8f124e500fe68058f0f069735230d5052458fad8b2b3df4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7a04d940baa1c06735d3537e1774a78db92e377acef16fbe53b9123ee552de3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49f12299f0d7a8194d0b081b935699734d021ed55a57b50516a697c26fb1ea0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha482da86f758574448c762b2b3486642700353fd87ca9c3601a18889ab2515c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b2832cb5c358d84d7fa692247d57dec68a1eb21d14f02794e70c19a69c2ba9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3459a275450e4f51635e7cad3fefdd375c5bff73ba438e86a7ee1ae7f04f6e9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e01b5f62195e5cdddc0c3b4947072c4f2b24ce3a70ef35ea8a38152e810f618;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfebf5df0014e1d5df97b1ce670e7ab5caeba3bbf32c6ed7af25de50e83a6f8a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f00fe65d90f47e6ec9bab9429a1a3cba97178dbc39ee14cab677795c70f5af6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c281c9a0286539941c6e5970b48fc150a4914da7cfaf7d5c2615a0ae29b7eff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he163d7b8069d277c616b4ade2606080e2becc6cd934d9dc125e4a3c7c01d2aaa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he694b9a68b0ffe4a593d5a20570cfdeedf51832c632f5fd87a0294f353801439;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4e8b5e2d3d78cd8703ec6a4bf374cbbc370cb696339a7bfdde632df3ff5a982;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91f296bc1b3e9e3e50a8b8c1311a4dca02f8a235f929ebc30e9372ce04b9270e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32caec59974d07655618dfd7704a0e7d4d031e88ae90a22e49f2ad71007d39b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e213d0c3599656ad14b07eed78b5cb5af295cee7efdcf53e69f7cdea158dd16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h711061f968d030adb407ba9c7954e757fcff62b41b4f1a134b8e90b92aa9194f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f232c9ac646fc7fb26bbfa9a82449f9b3bd896a45cbe63ad2537d2459cd2eac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc22ab5b7c3a7119259bdab486eedacaf16764782182b391f50939bc725cc95b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc2957f12e3ed56a88096e4342380996b45c683b19be0605b7807f089c507ae8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93733233b26d1720d146fc7cb8df92c5d5b287b658569e2f0bb6b80178a85bc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h609ba2fda46fd2041104a5168d6fcaa07a3973f0e570b4e7355496e7d7489057;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heaab7594b4566eeb45addaacc5c93f13ec2f5a85e26f45c64b1a7be90712695b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7b8be8d5b2b3bc48c01295172087b97d9d7d8a500c91e5846e36719b73c914b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25e91aed8906cdead022cc84e67125a380e414bf02f6d0fa9fe202cc73f7123e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h886b90a085557362f6b159dcf1b159aba82efd7ea90de47291072f838b4ff0f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5a6865ae8498cc85be3e5218d41e5426f36ed11ecbec2fbe0aaee685f10717b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf59b601a9a59789423f244465d7b6457cac648f0a1893390292026b21a3ec3c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a85435af49a83daf6a19f505ac1e6eae0fde14e165cd8987115880fbdc74fa4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbeeb61a7b140cbb1a698a759135b025c20322d979e07966ef5a72501302a93e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcae26e178df96d17a78953bc33e2162110bc182d6d434c79b42d6d478f3c3a27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h825ce2f62c4728b0c54c9fa8ac0f0299d10abc4b9578284c39292679b44543ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc442e311bbef89c5d1b71978b27a591c5952265a46d0b2596f3c28cef0e5277c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc90555d80015b311f3f6fddadc20d3c9e7a64631c9b4712dc92f0477dda2e90f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2cc5f6595baed76c7390633d6696ce67df6ffa4528a358b340d9ec09099d9a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c8a61d699052468d821a7cc57dabf44b11d4ee2e670271db4004c0bb5831015;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6302a07b7a55876b7b3134be8631651fee82b196c3b0e0147f7c557c9b4a0001;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h226831401475cf8ebc575088255c859b868825c8600f675cb221ef8532c37138;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd8d7efc2208a13fe472d7bcb77a750ae7a639a15fa24abbd29397a039922f17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75a9d8aa1c132375835fa91a691a852a0830e5a70ca54592073f702226f62c9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he08ef6e5ff6d01241ab379d11c108a79bf2d1eb2e9d22bf504f014325680fa00;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf84bf6e6fb9c9b81cb00151b8b89ca858c4f621e195e8cf8a6f013c5c0b11498;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2b98f1a6ca3136e50481236b4473604bd9d3a78ad2dcb0ae5d3c5cd02d2f93a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haef855a2b0ed8b0d8f8322e49299b997bf89804f2c218c14b361f694417ccc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1b79091d0e14caae10f5c70b83295dd125f1b99b03fda6e8d8986c29be176ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bb7945b911f8f8f9699819245cce99f4e294aebc482a476ff50fbe438622f6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e9fa86329a7d5be8dd5dadca49beb1472b842a191947be6b393c7b2542a9330;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30d9d33067f76cdb9d5134b9a9d4605cd088524f2f017968291d8ff5f60e77a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc41a68fd3c95c425bbb3ba329d860b609fdb014e710d5c4ed7a25bba9e004c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86e59df41e131684cde6ab888f7aac43d44625d2ee6892649931614da80e5114;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ca8fd108082990350511f4f01f4d921aa24789ce599090030649bd37896b123;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hecafcc43fb16834901ebfe935d15e185a367583b7f1a799b28c157f1d3e63f96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h245deebc9a0d392008198387ea980f6c0200c79e513a01ab758616dea5e108c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b9904d5f05a77d47ff0a209feacbf72d703ff8747c9cb2f009e2f85a97aa855;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23e24a547f91280485ba03d28548c2644a1a0a45a0d5a6b3efcfc6304d571e9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d1e16660e208f31aff8d873f285809d37624239c7c7d4fc199659bcd04d3f20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd60f8931da1a003aed72b7f7c21478ba2779989c07003153bee411baea06c2b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc41dae1655f55cd4613c12b0ec8d14f5095d5c50b6ca7a4acfaa0c3bb31e9d9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea557b1409924b208eaceddf34fd5a3dc5026272ecf0d6920887eee251cbc399;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e3e2c41ae1090b7311bfc25a3d702ce231919df600c6b436b1f24bb78ae027f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h933611a6b0bab94294e9ffd0a412552c49c376e97703e658fb901235bcf68e52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5218432d40986ff3e615f642b5d29c279ba89cb10b487f3424a90c268b6e5160;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h522ed363c932d8dbdf9761f8844ab1f6f6b740c2365ba20dd01d83e7a1726210;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he63d2da8ca29c4bfad48d759931c9ebf90a0ce2133cca312bbc23583d3d09965;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7aa2776bcadb7c12ca1d2ef3a23ac7b30eebb4a7579fb3547140308b0a1ea285;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d14e19dae0366aab3a527684ea585e33f67d44e6b88f2fa91a38b349bd9eaf5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6996bde9ca48d44e1cc35ef26744f03493a11c4132ed222ad4e12bd3a2a43ea9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17400cfef6feb5a7762099ba41954a3e3948d35c639f883f1eadcf9f5a5fe03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf956dd5887dd9e4bcfcb6c72d879dfb365fcb3de7d6638fcec9d180b733f74b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35d9e5a381210471c8553b60b9cacf62d4af84398ca2429bf706fbda0e3bafb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15691a430442419ddcd599be42aeb9ef4e6e70dc1e995d6ff66ee2cf378b25f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf457ad5c442d4e631963f610e868c330548aa18ef01812153d95927a6ffc655d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea9c5fafe1cb5e49773e2db0c164cc443efdc2c7a52f580b209b94c58482ace0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ed16313f9a889477bdf2ce89ff4af5bb86091c2e649bb6213417744874da3af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79be1e12695d47099a8e8a893c9846357b32bcb8eb0373623b4f688446be0c7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5d4f4d6974065bbd074f61d0afe518e30f1b3dc1ef9bb2ff3b7190154c178ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f88cc5e583e7ff378983e590eb9e176e5ec5aed655820470bd657e6803f780a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1800c2ed0bab17fa2d335d83b7709f498b4b7142f90a400425b73b980c4cb7bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca846a599f096674c51cf5a654e87a1a3b76c8a74d7bb74736d24a6eca3b16ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdae55e64b8e39355939b1fcb2e989a329aaf2b854d9fe27f34e76aaeee32e93d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73fd8eb582485e77d25cf76a50ea5237ee193249e3e36e9af09ee49c1ade8b24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e96703e9cbaddc03475acfecb956ba0f947eab483ea7eec35815a2535692481;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36f843b3babaf3f2d13447ace6eaf796d80d11b999a3c9f310ca0b8cf5b24272;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5332187d87e8e78c9119f0a053052a16f0bb333390a681db7b13035ecc2b8199;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he44dfa4fadaf69dfcbe9ca21b6c2817cf907a84fcf432905e89e27cadca95d54;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbd722ae2ca1ce9bc075246615a2f59bd2f99338eabd7425a43d286931f1aaea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9986fdb7229eefdf7070c5cb95c638fb32c7fbc65bd758754c545cf4dd851e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ef7650318c9c52e1af7d54f5ad6dc08ccdf63686e898d839ed3b5260d4e7b29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41ab8f076facb67678d7eb38d8866d23cfebe810fd1eaaf1c11d232614f23732;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22e3254e42ae96d9fd0630d3e3d5af66f1efd580417be33d45d607d12f01b22c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e1d71a66628e5b7eac6d3546d5736baf0de2b14addfc16fe27a78308dc5299;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he62fb4e364a756fbbf5a6b717c0755ea0b2130fbcff41b3f3421d02a096dcd1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd727ae422c9024f19b8670269575645ed0a4e88011814ae3095f2f46086d16c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2caf020e353c8b04c5851b56f073e44aac416e75c100e66cd04bba5cd921a24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2657a19a3fca1b68ba080ee3e6a20dc65131b26de524bda31d9b6f97487d69db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30979735d90949bd769340c076d8bdd69006b0cbc380c188d326a95252e605dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h602846bb811427bba2d73f92b7d6a30531f27eee3ce32b19a9fe3905b15168ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h499a71586ec5f08df090381eaa4edd02c144983393a4003a6bf2dc262ad4a14d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52c87a35bf8de7e3f0bfb5b4bfec0a9492f50a5542825436a31687b11b70be5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6540e13702ce4f227cc5ea7a9c4ca40a7ce7d5b5f0237f01274bd21159f3532b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a0cbc6b0e8edfa03e1fe7cdb03cd8a40d8f93e42227f22afe8ad9686f52bd72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1bd35d4a4f3db5b651cdd419eb86c8d7f558ff9f793c4b5593a5456466daa3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h167c6d8892fafbf691f9b01c2550682e606858866285c0f2c0e7c96f96a8c723;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ddaaa715a27232a6812e5613504a62b661c4e26f340539707414d206b261112;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a1d4ae2b856e81c7c92d2b21cc031f50d4a6388cb6b873fb32ff1816354e156;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fd3fd8419bcde69d4d313cdb8cc61e317ce0885dfae1583f1e9cc3ed3e7eaf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h215892a679eb08a47d729ba7dfc5c6dcd0620589cfaea796e0f1bfea246a9f90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e5aa9144e0275237038176c5dbe82f9c7be8ae5245591983398a8c7fc1f664;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eebb827d217700970caf870a7d748187d52824e86341e685cec27b9ac6ae819;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf880b81e01690500ab75b3049fbaa0a44ea6f2b38fc7e59a2be0821eb6f9e51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ff7e28b346ef81c5d3b7c2e648b6ca3b2153e0c4120ebb80092675ca22faea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56a437588436f8fa8ec2bc73c13172f8953a39e757cef6691724c030796e50c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e9d1570585f0c34a557c0444e3646b9eae1cbe4b205de5d8e87629c9ed4f175;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bf53faa86a2359cf221b6ec7c1d3884fd233e5ffa20fed04016b847d6a0df86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf24f41a0f7e0f06ac60aa150567ab42e1a0e5fdec2e051a49ec5b0ccf8c2d913;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cb6be9bed761e6813b8bed62f0b94d7493fef417afc0a5de8cba3df90099ee3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2b4664efdea5c72cdb24631303e2a2ae30f7a654c4e3083747370ca35c84140;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6573578a0f18a0184cafd1977e23ad51d58f14ba55602805fb9b740444720cbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c9ddf1c542e1252b57a3c5e61042b24b14800cbf03c180a6325bf732f128003;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bd72061b21d5d61dfd09d49d9b5ce9d9e1131359d080cbd2cf42fe0c733cd82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a289e01ac825651e51315645f09b7839a9701c5e2924468d9c4a19105dcfa60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdd94c7052eef917ddb6e2b5bced10949f3c1c750076946cb07d356d4b064af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h739280cb5663c11eecbbda38a8ed965917c4b2e46ffeb6e99a0bed0c6d828b5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f55b85bd5727a8e165e44333e6bd3230069f8978a3d281be6faffec2360c1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3a4bd62ae4b01e6ca7bba56a906bd22b7bc2a70466fb2d8c406af575b98baae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h149412ee01503d9cdbb2a720af1a28b29b7a14bbb4594d748919cfaa3702c75e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e6b5849f6547d8862b3758cc8853beb03061a25c7f66fd3e34021c90c8d3fa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf565913978c9b8ec71da5dff92a4ac820bc19c5855cfbffe9b9339851b622f3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc45f7940aaa8ae2906fafbda26f2e18db13411b80cd7fc2adfcad8695c8a2d14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1cb8ae8918083e056b52a306a17342e12d044c452a3eaa85a51a530ce34c133;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd31476d2dd62a160bfdc7d1e9c627e1ab70b2466d80d1315c3304d6f5f09bf0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h855497d947c26dfeceb59545f7bf306e4dbb7d5d8242e3cd1e40ebe063c8d168;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bcb386ea0e29f68ec234518586f0c7f306dab5e6c00422723687a5f8384dc0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1dd319d2f505c80f34efce6611520870a2d58611d79fe463b6a278c88e2b032;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb233a3bb52968788ce46ad5ccebcb8bda5a1b32175eaf066b47ede9519d5a80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb89d8644016517fc758eafe247abc3509b688bc518c03cd7c820775461b3994;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b79cab6c51fc615c0bd49ed11e7beb236a58b52f5c94351c8bbed7aab4366d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h665a0a4ca1f8fa55e2d11cbdd58d8914cdf674ae27078bda30e941e0e351168f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec85f26690d11b6312acc7c825c9026a73ca12f8133400e81496cea909c18826;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha270a7ac2065260e56ad177aab43517a848a165f9fdcfabb3a946a699698aa81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habdf719e165d2cc06c0cdcc9eedb34f2e84d20294b6b66d106a0c556e00d7db7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec5479d7607a4f5ed880ac65ec6cc76dc1694457949a30c5082c3f97dbec5c2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d40bb80ddf624462172b7f8c68a139e500cdbaf6753acf05c4a5b0525f5e126;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b5f92be29dcb50a6cdad28787567de2007c05d099d9bf0d914266033659927a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f27a3076c65fa1426bcebf89d2399992dc1bcf76fd9616e598af95456ee0710;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b03c44b8609f272f6ad44f472cfee0f6d4b9d82d97160c85014f83cd30823a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bd6ebf483af4516fd4c3cfa95a39385a0366d6fabdc837ff13e9be4bcc2190f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0c6ae1e86eded00dedf9785a7f21e5b6f791320d8af0d74e93ed3f494eef5a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h582dfca766a0249ee75eecf73ce414e9ff956d61f8465ed5c5ac3377ad82e098;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc0c7c6b69ccde4420469e50cdeff78e829df4881bb63d53a83d81bff1e454aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60474edc96c1841278f2e0c54475ae810cc1cab48613b966728d7ca2082bac44;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h295bd438269aef0077a75cad66e0d3a6e32ece3ec23e6cd74916ce4a39790b19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8803d09247b34fdafac8b78f0929ae273551a12aa9e89a48c23a51cba96815a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6165f1e4d44bc3b277053a2eb9fecb073220d936845c3c58ea903db9e0ad7572;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3b2e5fbd72bb56bc78ed7627a6569705d0255a1a4ec853d92099a45b066284a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7014a56495972565271f080e3743dfe16f5b48a55c5cdb5d694b63e18d9704a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcc34b858b82b401929d40660646a1a0610acf17b9f86c01f63eef8093be46f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha52880448e08a87a830a5cf51c3b72f09878fad804f0de95bcaf95ab7b64891b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9d810e641b4ab8acc29cbf8e1512f9362d90d2758ec4be66fccf8c0b893919e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89e4e0488698d8621cdb630d529f409892d8aa29f6278d3d4a8345d5adfcd687;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85f2ad442bc76d785b82b17a2c0db17597a5fd23890e553653b9592c44bd0a4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f0b0b0a668f35c47c05ae628d70c1358b64892062157b65708a02467466f70c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he853d5cecd3b26d3d114b090859727d57752121ca0568d3c5bae8cf57b3c9153;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28fe7e06ae8788405ed88741dd0ae7599b349e0551b49778d5accc3387980bbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4a03f9bab5911685ac6f1005bc27c6e701cfada3e49dcacbc17114be4c1e75b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98c66d70f00813011a676f6354d7f423ed58f8a8cd405ecf2ffeb81036056ae7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca9c904354194d0eec69a3168bc8b457bd1bf386f715bd7f462a23227b75d8b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe43f6223a18fa9235fbeccc609ef94500ad16f6f686c21f61b069cd9fa4f457;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedf62aaa7c39a22d62d38170b0dcb4315424d2ad67c7c882c09cf941cd26abbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h269844f9710e75ed0280fe6a69426fc5e64de46761ba59262c0a3a4e74264a63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c5ef2a3dea8899ac16d8efa1d1f1c069b3efc24ca86040dcaa224f6ba769504;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a1ee20f94f3b741a654085fd5b06cbc95816522759d4a6a18e6f16fb07822ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h121216f22a87eb6db37752f9c7b3ab160bb55526bfadff5f681874bf4f68a619;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7161f845ad4fbc36cb7efcfce3e7734df1b221ab91e8a5b4a2e7e8db91703b1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd94577fe3f5a69bcb212267a120f03297d55714a7da0a7507f96b137465bd052;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1bb66d16e7344e1ed0b3335bc63f046232c42e9014c7b9d36817ac34c0fef584;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1475063ae3c9396068fc13a689fd711b6a0703c1ad0fb7f2d5dccfebe7e198bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbb57e00a775eee1d87d3e5294427e22746e83c3a4bb76193803341573da6153;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40dfd0c77b4db7f461fc3ff7174be9d84f14de74c42848959c9dfe66227a7227;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h176e2fd818af9db4a9960534c80963c167d596bf593bb4a3e475c69d7512a198;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbae70b6b052dfc6e442af1504ed5ba39162f2b868cc7b210245b329f1f4befab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37b7515e172c561279bb65c6c919eafe11c1c95e67ee7b1f1bf7966f401efc21;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1221b2ecffcfb53b93b8bc90263848d6bb66d3ef26f63b94a09b2e24698d99a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ec25b1b553659156e1d2b4b1f5258ed75b88e54f06c03d590bb35d2539efbfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd60d70df92fbf5757f74cb5ce70b66b204ced3da9630f42ad0db6bb8ac15dc71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h467f090b5485a3ec0fa67739ff2a87f67cef5f92b1b18fa84088eef6da47ddf3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99ffaf824f602583c9c938b2962ff45dcacb5805b1278076de89304e5d6d1bed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40c8e584723c1fba3100b1d9b60a9a4e9e359646569695674fa9d29dbe229da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a5ae0a7891672b313212a5820e3c342ada815ce092f4de6f25a4753fc73fa06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69b1eeb694ed917f3ea15acf16bcdb481500abfe7dc7d4616cbaa50d5109dd5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he81fd7b8939f33180bde1d5045cac2c3f05f56d1af22839dbcc90cb7ade76b14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff9dc63e42b7dc3e296862cc8e2539a7ed094135fd17a60d14b5a7f08b6ae49f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1e43cd13a8ce0e6b5f8d9606ff32e9b3d2f843307f1db3323baa53f4be031da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe9f777d7b3d9acfe00f104cc7a2756429c0fc6b5eee57d81a795ce73d654175;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he539c495c822e06963b7c3a8e68fac4f99c93cc7f5dec9cd1d7e6af23d0bd084;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ed96dfaf0b49da0a3fd3ca6bace0e4503aeca369350913d282b4552e08d09e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42c85054c03693f65edadce7c3716fc77eebcc795f2fb6d6b053457ccf378393;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb72d91d1417f99175753146e164978061fd704020ec26300cbfb0e8cd634cdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe2aed1192cc2fa00f0e4f9d9597a505fcba592fec7bf9565ca684e60f0d775c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0fe88e3c37e5a7f1cc3e55aba8a93de5dbc41187201d1f34028bd9eaa69929;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he143d094fad1fa904a5ba4c4fab201209c37f6801121fd0e4685578a43a14524;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74379b4a91827ec011c8f3f5950564692ca31dc79c634b36d2dac82e7647cdff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3eaeac80dc9e21df336b03a214198489d78d481118303842b09a5ab74e4f9981;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe16111d88878976a483256a6e333ad9b5854553038eb5470376fb63a9048c20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd16307fc9bea8dc260493ac911f838dcf9f390c750283b238aae14a71d0bffa2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcbeaf4e6bce534f0607715f6886e8a5ae80719e191de022dacc2efb44247791;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2cb37ad32b78cd8b9c3079b531326669cf44d04a9978fe67152b1151e771703d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60fe618b8f0281ab5cc401374616badcc4a23014d95958a48873b262408e02fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76f8f7b729f5ece6aebd6f1fdf4d23ba25eb2a59c38514639f0ca51625945cdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81e65ef2d5c912aaf27aa6808a6183c8f8f50827404dae36ca2811616f3d4ccf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h110518df8b27ca4474e487abc8abf58504750813c8de0ddb5ada758591548b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d54f5127e2a1c0341ef8d9927cd6995ee38b91221ca85473af29a9c355d9aff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h677f02fdc95088b3b9ef356085cd4fc07a8096ffbb9e7e7dee351b63fff262bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ab1dca06bac7f5ae6a7c641e72e8a15488c7c6140ab6859212fb8b8d3f90e64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h303a36d7acc096fb2aa1b0490949bbd0d917d37537023fa290891e902ab4596d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heda547d59546525b2e8e89806ecc89bbc6f6dbcc43ccabfd5676e4b7ac41c528;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf636ca823172f0a293682576b27e0bc4c289ea675f6845e0dd040ee13da431dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58226871e7f22ece212cdeb3cb2227165b3e52182f5bdbbec4d4200ff6d179c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd27517313ee3f7fcc332df2e10dc0986daf9874ed2fa1833154576cd12676ea1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c1fda442069594f1c5dc4b730d143c15201d4916b8572a7ee93b626ddb98e78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h449be4af01006692e33c9defa5cf9329052c63449519285388b1fbcd9c594528;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1301659b35ed26da888c9f3d1e3f5dedb0e793ed9d178e3f51a5fa8ef63c68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9348047fdd91bda9652426e0fd243776ab06a89c2a3084f6511e091aea4309a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60473d46beeda81a9a95b4c2d58b5f5de83902eb0e0af238ecd87020709b3a0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f435967345a791b9f738e44baac127ec4bd740a23c912a449b817bdec2fef9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h457cd21e1214a5c8b6ebcccd6a82e9e13bacd8927f2f7a7dec259aaa8c0f0b4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cdabd8f7fa923758465bc587da73930c326acfda06261c77a64577eec25297e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26700d5d791dfb0869fe8a3cd3da6d2a2b6e3abfd0a313dcddf8c983697d05c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3153dc38b90a1d1b79ed4937f46a2c4449f7107e32322ac9dfc8c2fc8e220d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha81519a2b076579a6525eabfe175c6bd0af7b60fcd5120bb64f84c24b7f5d97e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9643bed5ba363b7eb4d4ecdacd51f3ce9b0651d04c438898ec0f1f20bb888b78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f817da7ec36a2f78b85bd3d4d3a63f9d13efdf8c01027048df3b0ced66395c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2b441c9b67d059b7c03f5708cd2a5e7a93e36dcf104a8d90150bc326ebe5601;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c4c32d15286c8448cefc12ef33a67067bb5b89a2b1ff69a1b219472b8c4b46e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8607c31edb36b765a949e458f2ceee4be97c5484c317fc6c80725cb45c0e8a31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78d78a29efb21a26b172a6ab5a33338fb2bc3c03d9ad0f290bc9556e0e1022e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd293334dc6e74342b963656b310f6af1287755737e6e8c977a6f1128be8b602;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b4a25a48f60486b38ee08eba0968542df6059f6ff94f669a03fce332d1dae34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6071c6b116b413573b2dff2f64a3b66c7e8f935285008d0e9bbe1f807d4d8521;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha229e82deacb80f61b59ed2f50a54c09942ec1f0a47af2f2ed704524f86fb7ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hace24d936d19903900ca965801d8fd39ca0dcf9fe82b97dd2a1e47cc6278ec8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h992bebede1cd9e93d843a2adcf97cbd8220d3352ab04bd58809ce12f782e3f04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6910598a5c8f67e092bfb66c8047f5ec1b36580f391204285d095cc28e321e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb57328701e8bbe68f54063d22591b287144bd49835a87e1afd86379119bca4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bf1a793a456d71c3329529650d840e685392f0ae6a61f3bc0854647759b597f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7d99709c151e766f39f6ab07586aae2d524c01a6830bc22d32392f51837ea25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4600f07cf5270c6acdc82aef75a1e7495c085d84e5e6275fdcf7640f9bd788e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e87f89200d5391f982bcba169b7a04a0d04a0adb4c86299f10ce8677c18b354;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e280f3d2b806b1265b01975965a1922ec5aab53254d17816cbf3f5ad31ce038;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4a2503076c53140f4c99ceb08fb1b605d7d42ee85970102be70b6ae8854e77a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h791003db5119e0e7fd715196bbe842e7eada9d5f3e6bc3e969360d49bda66aa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64d3feca9bda536ea6e2f90bb34416115102be91d4d04fae1646fdc4792bf467;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1419dc85e7f7f7f24443153e10199782c099fce80f24c46b153762081e4c1255;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae2c51e0aa3df9db820327b2ed5af54b6c2023ea2151560cf90dd72c8c872f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f614469a6bd5332c53bcac6e47ba9513c7bb5439176f89a2e155380ca93ac01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62cf0ceca7237ea1ae67e12e0ea18b0280a7fc366f9a8586c56783c0194409f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf99625b1ec7693de328f935ff82559b35c3a26171e5b740ae441fe5a967d4048;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he76524b4eac8383567be333f700afb71420f77ca430a7d8fcbb53725231fbd9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8797c6fdb3ac7f3dfc04e9aaff5846ae6539370b55a4fae33ce1e1b90ce0cee0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d3360a145843e3d88848709fc6e58210418c7302df27c404ad4f09f010bf4a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf010b106657429446563e9a1c81f2eee85c38523c6b31601b6c94205427509d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he75ebd3739fc16eb355dac9043905489b0064cfcdf0190c36f5c2ba1292e38c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5579762069460800ff9bbe437cf4432cb5a12eb3623a4e924c8656fe93452b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he94c469c39cc1150fc3027b92957f6442fd40e8eb75207956264b7a3a2389e6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba35ab88e7f73d4caff32c4de7939227fd48b5e7075771957ee56c82be6f9ade;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65d513fdfdebc64c419588e43dc981e2e4c7037545ed286496168dd651cba757;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2acdd0456bc55a8f97a7c3b0bf75c21da1a6bcc519b28a4c3ab6da11b805a11b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c2b788889c1810752aaaf32647f120e6501b1924c7295cfbd9ca795febc1389;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb6ba6e45e62c570b2d0b7af850a078f2f90ab75611cbd78479cad07f39b4e99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7dd6151ea4d038bd71ff5ec2ded2fa416b849512d78c898df5935ed1e559f2d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6eda2a989abb0aaac4f13cd44d2ac79d9aed0b27b89634ad433442129c0a44dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee3123fc7af7c1513fcdf402a37789efd5103698af0e395954b54f3565524a93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9b61bc2ef60ec179a3724ae8b1e8e64e542288c9e18817686971c0db0aeacec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a6d351562b651864e5aa10e337dd1779d41448827e563beafc8d4c64c9f2008;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97dcd05bb3d7724da5a9c0ee0f2e5602831302d3cac67292a672db14fc09aa5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34ace74e071eb6e0db468cb4c22d6dccfb5df4af137c724903e298710578468b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21935c93fc3fa7e27ffa0ff2e0ee6e514cfed51390bb739d34212259e4b0a90d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf446c65034c161edfb9bb3fa419af87537d9910d257a21587c8a2c86d1f91851;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb05ed176a7533ea18a3039e8543d97ae8e925fbfd8074e8a43f596aacc7baa2c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h601750c2d10cff0dab18cec39616227338834bccf968cc1096b63d3d43b48445;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72e7f70b704a34906b783bc596d47ab0e735fc8bb8110d6d1628b36ec3f9c633;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'headfd50da4c773dde4666310aed2ae8cebb25e77cd3c5cedbddd5a24c524aa3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1524ed483fb453cfff71b841d3d36043cafee29a48f664cc775ea3a9e73a211e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce69c0a4679d335aebcbb279111fb97e922c1e1c83b78b33b46bafe39af37054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93dbb7a2e70ab1b9541d8ff4fbcb1bce28b6608c82040c7b5fe1b3098f90d776;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h844e36c0ed43dbc6bb55053eebec01ca55647cc1245311f6e6374aae84be658a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38fedbea6bc733fff8e988f08df30bf98c1b24746f5bb7d80b42c731111a2abf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5a842f37b5c28013d796f101323443ef34be483a6517e10c40370e3951fc6a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc693d7f836fde9342efd44a7438ef33959d3a0e4b0f5df67e47d3356ff59fca8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hebb8068a2c7fe74d43e0929414bec7627ed2d1197fa5e25537e3573bfa2eaa27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e2f2108fc6da75c158a3f7dfb44de7fc9c4944ba9ed39e9c8f1c127159056f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h976a762e5f93379dcfaf5a83c56a87c070fd5e467df68ca964b57519e1fff094;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hecd168fa314157e6e548970af85ab8ce7f0abaa11ee9a9d236d9704b87835757;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc60ff857b98581a51ecf52cf524751ec8cf254a6bd178439c2a234d2a882b3aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7147e7ac591187b7cc077fd3a2656908c2a05b472de684e308fba598e136f407;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ee1e3d17f3fabdd9f426f3c86aaf8d957663091305cf1b287bd59db4dc23058;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4333abed9484bac939762b9e6762615e062c1593d3063c0de4e4762ce1012ce4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ad3847e73371c1faeb8580bb01d0ecf79e5e3834f51cf411c96f8533aa20cbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e7af0ccf96eb988e8b7fd1ecce1d0c46a8cf212dd6b40394669ed9d125e25cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hebfa5fbc6a1f7da37f9ff12b6df1ebc8acdff63126ebc6f357952194058a1684;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2532936061b9b76f80199abe379403441d18b187dc779587fb193844b74f6c1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85f900873f7bb7e4b5346a83667693d1bc8d5e7f51b2a5b42e88bf01807a44af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he71bf221b3ab7e3c3e70a67b63ac9e71b6977dc13746f54ed1445967940c6050;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d25d8b5dadbef8a5b31aa909cb610574a964e865bcb2e64dbd53cae91e332fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc61cfbad795f0102c301dfa19dc74dd73d082cb8f9a4762711c3c31378a0a8b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf78d96501bd2b67ac893bf0448a7f460d9fddf19f0658d49a580376bf8401dac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h848dfeaa8980aa1159e7311ae103ec5c298c9315c612de13f43ae13cccac063;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b77794019e082a9f843af52544aaadd65bb5be34e91d1c09d83e49778e26370;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcd9de1262dbe6722349383ad8f8ab37749e10c2edf03d291c0bbe0721256bc1;
        #1
        $finish();
    end
endmodule
