module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    compressor2_1_162_12 compressor2_1_162_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_162_12(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [0:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    rowadder2_1_19 rowadder2_1inst(
        .src0({comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], 1'h0, comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst0({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [0:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [30:0] stage1_0;
   wire [52:0] stage1_1;
   wire [65:0] stage1_2;
   wire [57:0] stage1_3;
   wire [138:0] stage1_4;
   wire [67:0] stage1_5;
   wire [111:0] stage1_6;
   wire [47:0] stage1_7;
   wire [72:0] stage1_8;
   wire [78:0] stage1_9;
   wire [58:0] stage1_10;
   wire [52:0] stage1_11;
   wire [52:0] stage1_12;
   wire [26:0] stage1_13;
   wire [18:0] stage2_0;
   wire [22:0] stage2_1;
   wire [26:0] stage2_2;
   wire [32:0] stage2_3;
   wire [44:0] stage2_4;
   wire [37:0] stage2_5;
   wire [49:0] stage2_6;
   wire [33:0] stage2_7;
   wire [41:0] stage2_8;
   wire [29:0] stage2_9;
   wire [29:0] stage2_10;
   wire [24:0] stage2_11;
   wire [27:0] stage2_12;
   wire [28:0] stage2_13;
   wire [8:0] stage2_14;
   wire [2:0] stage2_15;
   wire [11:0] stage3_0;
   wire [13:0] stage3_1;
   wire [18:0] stage3_2;
   wire [14:0] stage3_3;
   wire [18:0] stage3_4;
   wire [17:0] stage3_5;
   wire [17:0] stage3_6;
   wire [18:0] stage3_7;
   wire [16:0] stage3_8;
   wire [11:0] stage3_9;
   wire [13:0] stage3_10;
   wire [17:0] stage3_11;
   wire [9:0] stage3_12;
   wire [12:0] stage3_13;
   wire [10:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [15:0] stage4_2;
   wire [5:0] stage4_3;
   wire [6:0] stage4_4;
   wire [7:0] stage4_5;
   wire [5:0] stage4_6;
   wire [6:0] stage4_7;
   wire [9:0] stage4_8;
   wire [6:0] stage4_9;
   wire [5:0] stage4_10;
   wire [5:0] stage4_11;
   wire [8:0] stage4_12;
   wire [4:0] stage4_13;
   wire [8:0] stage4_14;
   wire [4:0] stage4_15;
   wire [2:0] stage4_16;
   wire [0:0] stage4_17;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [4:0] stage5_2;
   wire [5:0] stage5_3;
   wire [2:0] stage5_4;
   wire [5:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [5:0] stage5_8;
   wire [3:0] stage5_9;
   wire [2:0] stage5_10;
   wire [1:0] stage5_11;
   wire [2:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [4:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [0:0] stage5_18;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [0:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [0:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc615_5 gpc23 (
      {stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[12]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc615_5 gpc24 (
      {stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143]},
      {stage0_1[13]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc615_5 gpc25 (
      {stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148]},
      {stage0_1[14]},
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc615_5 gpc26 (
      {stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[15]},
      {stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc615_5 gpc27 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_1[16]},
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[0],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[1],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[2],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[3],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[4],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[5],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[6],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[7],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[8],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[9],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[10],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[11],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85]},
      {stage1_5[12],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100]},
      {stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage1_5[13],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106]},
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97]},
      {stage1_5[14],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112]},
      {stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage1_5[15],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118]},
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109]},
      {stage1_5[16],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124]},
      {stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115]},
      {stage1_5[17],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130]},
      {stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121]},
      {stage1_5[18],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136]},
      {stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127]},
      {stage1_5[19],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142]},
      {stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage1_5[20],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148]},
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage1_5[21],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154]},
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145]},
      {stage1_5[22],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160]},
      {stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151]},
      {stage1_5[23],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc615_5 gpc52 (
      {stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage0_4[0]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[24],stage1_4[52],stage1_3[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[25],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[26],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[27],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[28],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[29],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[30],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[31],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[32],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[33],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[34],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[35],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[36],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[37],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[38],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[39],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[15],stage1_7[16],stage1_6[16],stage1_5[40]}
   );
   gpc606_5 gpc69 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[16],stage1_7[17],stage1_6[17],stage1_5[41]}
   );
   gpc606_5 gpc70 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[17],stage1_7[18],stage1_6[18],stage1_5[42]}
   );
   gpc606_5 gpc71 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[18],stage1_7[19],stage1_6[19],stage1_5[43]}
   );
   gpc606_5 gpc72 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[19],stage1_7[20],stage1_6[20],stage1_5[44]}
   );
   gpc606_5 gpc73 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[20],stage1_7[21],stage1_6[21],stage1_5[45]}
   );
   gpc606_5 gpc74 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[21],stage1_7[22],stage1_6[22],stage1_5[46]}
   );
   gpc606_5 gpc75 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[22],stage1_7[23],stage1_6[23],stage1_5[47]}
   );
   gpc606_5 gpc76 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[23],stage1_7[24],stage1_6[24],stage1_5[48]}
   );
   gpc606_5 gpc77 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[24],stage1_7[25],stage1_6[25],stage1_5[49]}
   );
   gpc606_5 gpc78 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[25],stage1_7[26],stage1_6[26],stage1_5[50]}
   );
   gpc606_5 gpc79 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[26],stage1_7[27],stage1_6[27],stage1_5[51]}
   );
   gpc606_5 gpc80 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[27],stage1_7[28],stage1_6[28],stage1_5[52]}
   );
   gpc606_5 gpc81 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[28],stage1_7[29],stage1_6[29],stage1_5[53]}
   );
   gpc606_5 gpc82 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[29],stage1_7[30],stage1_6[30],stage1_5[54]}
   );
   gpc606_5 gpc83 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[30],stage1_7[31],stage1_6[31],stage1_5[55]}
   );
   gpc606_5 gpc84 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[31],stage1_7[32],stage1_6[32],stage1_5[56]}
   );
   gpc606_5 gpc85 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[32],stage1_7[33],stage1_6[33],stage1_5[57]}
   );
   gpc606_5 gpc86 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[33],stage1_7[34],stage1_6[34],stage1_5[58]}
   );
   gpc606_5 gpc87 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[34],stage1_7[35],stage1_6[35],stage1_5[59]}
   );
   gpc606_5 gpc88 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[35],stage1_7[36],stage1_6[36],stage1_5[60]}
   );
   gpc606_5 gpc89 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[36],stage1_7[37],stage1_6[37],stage1_5[61]}
   );
   gpc606_5 gpc90 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[37],stage1_7[38],stage1_6[38],stage1_5[62]}
   );
   gpc606_5 gpc91 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[38],stage1_7[39],stage1_6[39],stage1_5[63]}
   );
   gpc615_5 gpc92 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154]},
      {stage0_6[90]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[39],stage1_7[40],stage1_6[40],stage1_5[64]}
   );
   gpc615_5 gpc93 (
      {stage0_5[155], stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159]},
      {stage0_6[91]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[40],stage1_7[41],stage1_6[41],stage1_5[65]}
   );
   gpc606_5 gpc94 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[0],stage1_9[26],stage1_8[41]}
   );
   gpc606_5 gpc95 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[1],stage1_9[27],stage1_8[42]}
   );
   gpc606_5 gpc96 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[2],stage1_9[28],stage1_8[43]}
   );
   gpc606_5 gpc97 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[3],stage1_9[29],stage1_8[44]}
   );
   gpc606_5 gpc98 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[4],stage1_9[30],stage1_8[45]}
   );
   gpc606_5 gpc99 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[5],stage1_9[31],stage1_8[46]}
   );
   gpc606_5 gpc100 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[6],stage1_9[32],stage1_8[47]}
   );
   gpc606_5 gpc101 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[7],stage1_9[33],stage1_8[48]}
   );
   gpc606_5 gpc102 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[8],stage1_9[34],stage1_8[49]}
   );
   gpc606_5 gpc103 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[9],stage1_9[35],stage1_8[50]}
   );
   gpc606_5 gpc104 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[10],stage1_9[36],stage1_8[51]}
   );
   gpc606_5 gpc105 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[11],stage1_9[37],stage1_8[52]}
   );
   gpc606_5 gpc106 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[12],stage1_9[38],stage1_8[53]}
   );
   gpc606_5 gpc107 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[13],stage1_9[39],stage1_8[54]}
   );
   gpc606_5 gpc108 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[14],stage1_9[40],stage1_8[55]}
   );
   gpc606_5 gpc109 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[15],stage1_9[41],stage1_8[56]}
   );
   gpc606_5 gpc110 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[16],stage1_9[42],stage1_8[57]}
   );
   gpc606_5 gpc111 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[17],stage1_9[43],stage1_8[58]}
   );
   gpc606_5 gpc112 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[18],stage1_9[44],stage1_8[59]}
   );
   gpc606_5 gpc113 (
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[19],stage1_9[45],stage1_8[60]}
   );
   gpc606_5 gpc114 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[20],stage1_9[46],stage1_8[61]}
   );
   gpc606_5 gpc115 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[21],stage1_10[21],stage1_9[47],stage1_8[62]}
   );
   gpc606_5 gpc116 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[22],stage1_10[22],stage1_9[48],stage1_8[63]}
   );
   gpc606_5 gpc117 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[23],stage1_10[23],stage1_9[49],stage1_8[64]}
   );
   gpc606_5 gpc118 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[24],stage1_10[24],stage1_9[50],stage1_8[65]}
   );
   gpc606_5 gpc119 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[25],stage1_10[25],stage1_9[51],stage1_8[66]}
   );
   gpc606_5 gpc120 (
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[26],stage1_11[26],stage1_10[26],stage1_9[52]}
   );
   gpc606_5 gpc121 (
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[27],stage1_11[27],stage1_10[27],stage1_9[53]}
   );
   gpc606_5 gpc122 (
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[28],stage1_11[28],stage1_10[28],stage1_9[54]}
   );
   gpc606_5 gpc123 (
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[29],stage1_11[29],stage1_10[29],stage1_9[55]}
   );
   gpc606_5 gpc124 (
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[30],stage1_11[30],stage1_10[30],stage1_9[56]}
   );
   gpc606_5 gpc125 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[31],stage1_11[31],stage1_10[31],stage1_9[57]}
   );
   gpc606_5 gpc126 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[32],stage1_11[32],stage1_10[32],stage1_9[58]}
   );
   gpc606_5 gpc127 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[33],stage1_11[33],stage1_10[33],stage1_9[59]}
   );
   gpc606_5 gpc128 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[34],stage1_11[34],stage1_10[34],stage1_9[60]}
   );
   gpc606_5 gpc129 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[35],stage1_11[35],stage1_10[35],stage1_9[61]}
   );
   gpc606_5 gpc130 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[36],stage1_11[36],stage1_10[36],stage1_9[62]}
   );
   gpc606_5 gpc131 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[37],stage1_11[37],stage1_10[37],stage1_9[63]}
   );
   gpc606_5 gpc132 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[38],stage1_11[38],stage1_10[38],stage1_9[64]}
   );
   gpc606_5 gpc133 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[39],stage1_11[39],stage1_10[39],stage1_9[65]}
   );
   gpc606_5 gpc134 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[40],stage1_11[40],stage1_10[40],stage1_9[66]}
   );
   gpc606_5 gpc135 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[41],stage1_11[41],stage1_10[41],stage1_9[67]}
   );
   gpc606_5 gpc136 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[42],stage1_11[42],stage1_10[42],stage1_9[68]}
   );
   gpc606_5 gpc137 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[43],stage1_11[43],stage1_10[43],stage1_9[69]}
   );
   gpc606_5 gpc138 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[44],stage1_11[44],stage1_10[44],stage1_9[70]}
   );
   gpc606_5 gpc139 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[45],stage1_11[45],stage1_10[45],stage1_9[71]}
   );
   gpc606_5 gpc140 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[46],stage1_11[46],stage1_10[46],stage1_9[72]}
   );
   gpc606_5 gpc141 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[47],stage1_11[47],stage1_10[47],stage1_9[73]}
   );
   gpc606_5 gpc142 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[48],stage1_11[48],stage1_10[48],stage1_9[74]}
   );
   gpc606_5 gpc143 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[49],stage1_11[49],stage1_10[49],stage1_9[75]}
   );
   gpc606_5 gpc144 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[50],stage1_11[50],stage1_10[50],stage1_9[76]}
   );
   gpc606_5 gpc145 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[51],stage1_11[51],stage1_10[51],stage1_9[77]}
   );
   gpc606_5 gpc146 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[52],stage1_11[52],stage1_10[52],stage1_9[78]}
   );
   gpc1_1 gpc147 (
      {stage0_0[159]},
      {stage1_0[28]}
   );
   gpc1_1 gpc148 (
      {stage0_0[160]},
      {stage1_0[29]}
   );
   gpc1_1 gpc149 (
      {stage0_0[161]},
      {stage1_0[30]}
   );
   gpc1_1 gpc150 (
      {stage0_1[161]},
      {stage1_1[52]}
   );
   gpc1_1 gpc151 (
      {stage0_2[148]},
      {stage1_2[52]}
   );
   gpc1_1 gpc152 (
      {stage0_2[149]},
      {stage1_2[53]}
   );
   gpc1_1 gpc153 (
      {stage0_2[150]},
      {stage1_2[54]}
   );
   gpc1_1 gpc154 (
      {stage0_2[151]},
      {stage1_2[55]}
   );
   gpc1_1 gpc155 (
      {stage0_2[152]},
      {stage1_2[56]}
   );
   gpc1_1 gpc156 (
      {stage0_2[153]},
      {stage1_2[57]}
   );
   gpc1_1 gpc157 (
      {stage0_2[154]},
      {stage1_2[58]}
   );
   gpc1_1 gpc158 (
      {stage0_2[155]},
      {stage1_2[59]}
   );
   gpc1_1 gpc159 (
      {stage0_2[156]},
      {stage1_2[60]}
   );
   gpc1_1 gpc160 (
      {stage0_2[157]},
      {stage1_2[61]}
   );
   gpc1_1 gpc161 (
      {stage0_2[158]},
      {stage1_2[62]}
   );
   gpc1_1 gpc162 (
      {stage0_2[159]},
      {stage1_2[63]}
   );
   gpc1_1 gpc163 (
      {stage0_2[160]},
      {stage1_2[64]}
   );
   gpc1_1 gpc164 (
      {stage0_2[161]},
      {stage1_2[65]}
   );
   gpc1_1 gpc165 (
      {stage0_3[157]},
      {stage1_3[53]}
   );
   gpc1_1 gpc166 (
      {stage0_3[158]},
      {stage1_3[54]}
   );
   gpc1_1 gpc167 (
      {stage0_3[159]},
      {stage1_3[55]}
   );
   gpc1_1 gpc168 (
      {stage0_3[160]},
      {stage1_3[56]}
   );
   gpc1_1 gpc169 (
      {stage0_3[161]},
      {stage1_3[57]}
   );
   gpc1_1 gpc170 (
      {stage0_4[91]},
      {stage1_4[68]}
   );
   gpc1_1 gpc171 (
      {stage0_4[92]},
      {stage1_4[69]}
   );
   gpc1_1 gpc172 (
      {stage0_4[93]},
      {stage1_4[70]}
   );
   gpc1_1 gpc173 (
      {stage0_4[94]},
      {stage1_4[71]}
   );
   gpc1_1 gpc174 (
      {stage0_4[95]},
      {stage1_4[72]}
   );
   gpc1_1 gpc175 (
      {stage0_4[96]},
      {stage1_4[73]}
   );
   gpc1_1 gpc176 (
      {stage0_4[97]},
      {stage1_4[74]}
   );
   gpc1_1 gpc177 (
      {stage0_4[98]},
      {stage1_4[75]}
   );
   gpc1_1 gpc178 (
      {stage0_4[99]},
      {stage1_4[76]}
   );
   gpc1_1 gpc179 (
      {stage0_4[100]},
      {stage1_4[77]}
   );
   gpc1_1 gpc180 (
      {stage0_4[101]},
      {stage1_4[78]}
   );
   gpc1_1 gpc181 (
      {stage0_4[102]},
      {stage1_4[79]}
   );
   gpc1_1 gpc182 (
      {stage0_4[103]},
      {stage1_4[80]}
   );
   gpc1_1 gpc183 (
      {stage0_4[104]},
      {stage1_4[81]}
   );
   gpc1_1 gpc184 (
      {stage0_4[105]},
      {stage1_4[82]}
   );
   gpc1_1 gpc185 (
      {stage0_4[106]},
      {stage1_4[83]}
   );
   gpc1_1 gpc186 (
      {stage0_4[107]},
      {stage1_4[84]}
   );
   gpc1_1 gpc187 (
      {stage0_4[108]},
      {stage1_4[85]}
   );
   gpc1_1 gpc188 (
      {stage0_4[109]},
      {stage1_4[86]}
   );
   gpc1_1 gpc189 (
      {stage0_4[110]},
      {stage1_4[87]}
   );
   gpc1_1 gpc190 (
      {stage0_4[111]},
      {stage1_4[88]}
   );
   gpc1_1 gpc191 (
      {stage0_4[112]},
      {stage1_4[89]}
   );
   gpc1_1 gpc192 (
      {stage0_4[113]},
      {stage1_4[90]}
   );
   gpc1_1 gpc193 (
      {stage0_4[114]},
      {stage1_4[91]}
   );
   gpc1_1 gpc194 (
      {stage0_4[115]},
      {stage1_4[92]}
   );
   gpc1_1 gpc195 (
      {stage0_4[116]},
      {stage1_4[93]}
   );
   gpc1_1 gpc196 (
      {stage0_4[117]},
      {stage1_4[94]}
   );
   gpc1_1 gpc197 (
      {stage0_4[118]},
      {stage1_4[95]}
   );
   gpc1_1 gpc198 (
      {stage0_4[119]},
      {stage1_4[96]}
   );
   gpc1_1 gpc199 (
      {stage0_4[120]},
      {stage1_4[97]}
   );
   gpc1_1 gpc200 (
      {stage0_4[121]},
      {stage1_4[98]}
   );
   gpc1_1 gpc201 (
      {stage0_4[122]},
      {stage1_4[99]}
   );
   gpc1_1 gpc202 (
      {stage0_4[123]},
      {stage1_4[100]}
   );
   gpc1_1 gpc203 (
      {stage0_4[124]},
      {stage1_4[101]}
   );
   gpc1_1 gpc204 (
      {stage0_4[125]},
      {stage1_4[102]}
   );
   gpc1_1 gpc205 (
      {stage0_4[126]},
      {stage1_4[103]}
   );
   gpc1_1 gpc206 (
      {stage0_4[127]},
      {stage1_4[104]}
   );
   gpc1_1 gpc207 (
      {stage0_4[128]},
      {stage1_4[105]}
   );
   gpc1_1 gpc208 (
      {stage0_4[129]},
      {stage1_4[106]}
   );
   gpc1_1 gpc209 (
      {stage0_4[130]},
      {stage1_4[107]}
   );
   gpc1_1 gpc210 (
      {stage0_4[131]},
      {stage1_4[108]}
   );
   gpc1_1 gpc211 (
      {stage0_4[132]},
      {stage1_4[109]}
   );
   gpc1_1 gpc212 (
      {stage0_4[133]},
      {stage1_4[110]}
   );
   gpc1_1 gpc213 (
      {stage0_4[134]},
      {stage1_4[111]}
   );
   gpc1_1 gpc214 (
      {stage0_4[135]},
      {stage1_4[112]}
   );
   gpc1_1 gpc215 (
      {stage0_4[136]},
      {stage1_4[113]}
   );
   gpc1_1 gpc216 (
      {stage0_4[137]},
      {stage1_4[114]}
   );
   gpc1_1 gpc217 (
      {stage0_4[138]},
      {stage1_4[115]}
   );
   gpc1_1 gpc218 (
      {stage0_4[139]},
      {stage1_4[116]}
   );
   gpc1_1 gpc219 (
      {stage0_4[140]},
      {stage1_4[117]}
   );
   gpc1_1 gpc220 (
      {stage0_4[141]},
      {stage1_4[118]}
   );
   gpc1_1 gpc221 (
      {stage0_4[142]},
      {stage1_4[119]}
   );
   gpc1_1 gpc222 (
      {stage0_4[143]},
      {stage1_4[120]}
   );
   gpc1_1 gpc223 (
      {stage0_4[144]},
      {stage1_4[121]}
   );
   gpc1_1 gpc224 (
      {stage0_4[145]},
      {stage1_4[122]}
   );
   gpc1_1 gpc225 (
      {stage0_4[146]},
      {stage1_4[123]}
   );
   gpc1_1 gpc226 (
      {stage0_4[147]},
      {stage1_4[124]}
   );
   gpc1_1 gpc227 (
      {stage0_4[148]},
      {stage1_4[125]}
   );
   gpc1_1 gpc228 (
      {stage0_4[149]},
      {stage1_4[126]}
   );
   gpc1_1 gpc229 (
      {stage0_4[150]},
      {stage1_4[127]}
   );
   gpc1_1 gpc230 (
      {stage0_4[151]},
      {stage1_4[128]}
   );
   gpc1_1 gpc231 (
      {stage0_4[152]},
      {stage1_4[129]}
   );
   gpc1_1 gpc232 (
      {stage0_4[153]},
      {stage1_4[130]}
   );
   gpc1_1 gpc233 (
      {stage0_4[154]},
      {stage1_4[131]}
   );
   gpc1_1 gpc234 (
      {stage0_4[155]},
      {stage1_4[132]}
   );
   gpc1_1 gpc235 (
      {stage0_4[156]},
      {stage1_4[133]}
   );
   gpc1_1 gpc236 (
      {stage0_4[157]},
      {stage1_4[134]}
   );
   gpc1_1 gpc237 (
      {stage0_4[158]},
      {stage1_4[135]}
   );
   gpc1_1 gpc238 (
      {stage0_4[159]},
      {stage1_4[136]}
   );
   gpc1_1 gpc239 (
      {stage0_4[160]},
      {stage1_4[137]}
   );
   gpc1_1 gpc240 (
      {stage0_4[161]},
      {stage1_4[138]}
   );
   gpc1_1 gpc241 (
      {stage0_5[160]},
      {stage1_5[66]}
   );
   gpc1_1 gpc242 (
      {stage0_5[161]},
      {stage1_5[67]}
   );
   gpc1_1 gpc243 (
      {stage0_6[92]},
      {stage1_6[42]}
   );
   gpc1_1 gpc244 (
      {stage0_6[93]},
      {stage1_6[43]}
   );
   gpc1_1 gpc245 (
      {stage0_6[94]},
      {stage1_6[44]}
   );
   gpc1_1 gpc246 (
      {stage0_6[95]},
      {stage1_6[45]}
   );
   gpc1_1 gpc247 (
      {stage0_6[96]},
      {stage1_6[46]}
   );
   gpc1_1 gpc248 (
      {stage0_6[97]},
      {stage1_6[47]}
   );
   gpc1_1 gpc249 (
      {stage0_6[98]},
      {stage1_6[48]}
   );
   gpc1_1 gpc250 (
      {stage0_6[99]},
      {stage1_6[49]}
   );
   gpc1_1 gpc251 (
      {stage0_6[100]},
      {stage1_6[50]}
   );
   gpc1_1 gpc252 (
      {stage0_6[101]},
      {stage1_6[51]}
   );
   gpc1_1 gpc253 (
      {stage0_6[102]},
      {stage1_6[52]}
   );
   gpc1_1 gpc254 (
      {stage0_6[103]},
      {stage1_6[53]}
   );
   gpc1_1 gpc255 (
      {stage0_6[104]},
      {stage1_6[54]}
   );
   gpc1_1 gpc256 (
      {stage0_6[105]},
      {stage1_6[55]}
   );
   gpc1_1 gpc257 (
      {stage0_6[106]},
      {stage1_6[56]}
   );
   gpc1_1 gpc258 (
      {stage0_6[107]},
      {stage1_6[57]}
   );
   gpc1_1 gpc259 (
      {stage0_6[108]},
      {stage1_6[58]}
   );
   gpc1_1 gpc260 (
      {stage0_6[109]},
      {stage1_6[59]}
   );
   gpc1_1 gpc261 (
      {stage0_6[110]},
      {stage1_6[60]}
   );
   gpc1_1 gpc262 (
      {stage0_6[111]},
      {stage1_6[61]}
   );
   gpc1_1 gpc263 (
      {stage0_6[112]},
      {stage1_6[62]}
   );
   gpc1_1 gpc264 (
      {stage0_6[113]},
      {stage1_6[63]}
   );
   gpc1_1 gpc265 (
      {stage0_6[114]},
      {stage1_6[64]}
   );
   gpc1_1 gpc266 (
      {stage0_6[115]},
      {stage1_6[65]}
   );
   gpc1_1 gpc267 (
      {stage0_6[116]},
      {stage1_6[66]}
   );
   gpc1_1 gpc268 (
      {stage0_6[117]},
      {stage1_6[67]}
   );
   gpc1_1 gpc269 (
      {stage0_6[118]},
      {stage1_6[68]}
   );
   gpc1_1 gpc270 (
      {stage0_6[119]},
      {stage1_6[69]}
   );
   gpc1_1 gpc271 (
      {stage0_6[120]},
      {stage1_6[70]}
   );
   gpc1_1 gpc272 (
      {stage0_6[121]},
      {stage1_6[71]}
   );
   gpc1_1 gpc273 (
      {stage0_6[122]},
      {stage1_6[72]}
   );
   gpc1_1 gpc274 (
      {stage0_6[123]},
      {stage1_6[73]}
   );
   gpc1_1 gpc275 (
      {stage0_6[124]},
      {stage1_6[74]}
   );
   gpc1_1 gpc276 (
      {stage0_6[125]},
      {stage1_6[75]}
   );
   gpc1_1 gpc277 (
      {stage0_6[126]},
      {stage1_6[76]}
   );
   gpc1_1 gpc278 (
      {stage0_6[127]},
      {stage1_6[77]}
   );
   gpc1_1 gpc279 (
      {stage0_6[128]},
      {stage1_6[78]}
   );
   gpc1_1 gpc280 (
      {stage0_6[129]},
      {stage1_6[79]}
   );
   gpc1_1 gpc281 (
      {stage0_6[130]},
      {stage1_6[80]}
   );
   gpc1_1 gpc282 (
      {stage0_6[131]},
      {stage1_6[81]}
   );
   gpc1_1 gpc283 (
      {stage0_6[132]},
      {stage1_6[82]}
   );
   gpc1_1 gpc284 (
      {stage0_6[133]},
      {stage1_6[83]}
   );
   gpc1_1 gpc285 (
      {stage0_6[134]},
      {stage1_6[84]}
   );
   gpc1_1 gpc286 (
      {stage0_6[135]},
      {stage1_6[85]}
   );
   gpc1_1 gpc287 (
      {stage0_6[136]},
      {stage1_6[86]}
   );
   gpc1_1 gpc288 (
      {stage0_6[137]},
      {stage1_6[87]}
   );
   gpc1_1 gpc289 (
      {stage0_6[138]},
      {stage1_6[88]}
   );
   gpc1_1 gpc290 (
      {stage0_6[139]},
      {stage1_6[89]}
   );
   gpc1_1 gpc291 (
      {stage0_6[140]},
      {stage1_6[90]}
   );
   gpc1_1 gpc292 (
      {stage0_6[141]},
      {stage1_6[91]}
   );
   gpc1_1 gpc293 (
      {stage0_6[142]},
      {stage1_6[92]}
   );
   gpc1_1 gpc294 (
      {stage0_6[143]},
      {stage1_6[93]}
   );
   gpc1_1 gpc295 (
      {stage0_6[144]},
      {stage1_6[94]}
   );
   gpc1_1 gpc296 (
      {stage0_6[145]},
      {stage1_6[95]}
   );
   gpc1_1 gpc297 (
      {stage0_6[146]},
      {stage1_6[96]}
   );
   gpc1_1 gpc298 (
      {stage0_6[147]},
      {stage1_6[97]}
   );
   gpc1_1 gpc299 (
      {stage0_6[148]},
      {stage1_6[98]}
   );
   gpc1_1 gpc300 (
      {stage0_6[149]},
      {stage1_6[99]}
   );
   gpc1_1 gpc301 (
      {stage0_6[150]},
      {stage1_6[100]}
   );
   gpc1_1 gpc302 (
      {stage0_6[151]},
      {stage1_6[101]}
   );
   gpc1_1 gpc303 (
      {stage0_6[152]},
      {stage1_6[102]}
   );
   gpc1_1 gpc304 (
      {stage0_6[153]},
      {stage1_6[103]}
   );
   gpc1_1 gpc305 (
      {stage0_6[154]},
      {stage1_6[104]}
   );
   gpc1_1 gpc306 (
      {stage0_6[155]},
      {stage1_6[105]}
   );
   gpc1_1 gpc307 (
      {stage0_6[156]},
      {stage1_6[106]}
   );
   gpc1_1 gpc308 (
      {stage0_6[157]},
      {stage1_6[107]}
   );
   gpc1_1 gpc309 (
      {stage0_6[158]},
      {stage1_6[108]}
   );
   gpc1_1 gpc310 (
      {stage0_6[159]},
      {stage1_6[109]}
   );
   gpc1_1 gpc311 (
      {stage0_6[160]},
      {stage1_6[110]}
   );
   gpc1_1 gpc312 (
      {stage0_6[161]},
      {stage1_6[111]}
   );
   gpc1_1 gpc313 (
      {stage0_7[156]},
      {stage1_7[42]}
   );
   gpc1_1 gpc314 (
      {stage0_7[157]},
      {stage1_7[43]}
   );
   gpc1_1 gpc315 (
      {stage0_7[158]},
      {stage1_7[44]}
   );
   gpc1_1 gpc316 (
      {stage0_7[159]},
      {stage1_7[45]}
   );
   gpc1_1 gpc317 (
      {stage0_7[160]},
      {stage1_7[46]}
   );
   gpc1_1 gpc318 (
      {stage0_7[161]},
      {stage1_7[47]}
   );
   gpc1_1 gpc319 (
      {stage0_8[156]},
      {stage1_8[67]}
   );
   gpc1_1 gpc320 (
      {stage0_8[157]},
      {stage1_8[68]}
   );
   gpc1_1 gpc321 (
      {stage0_8[158]},
      {stage1_8[69]}
   );
   gpc1_1 gpc322 (
      {stage0_8[159]},
      {stage1_8[70]}
   );
   gpc1_1 gpc323 (
      {stage0_8[160]},
      {stage1_8[71]}
   );
   gpc1_1 gpc324 (
      {stage0_8[161]},
      {stage1_8[72]}
   );
   gpc1_1 gpc325 (
      {stage0_10[156]},
      {stage1_10[53]}
   );
   gpc1_1 gpc326 (
      {stage0_10[157]},
      {stage1_10[54]}
   );
   gpc1_1 gpc327 (
      {stage0_10[158]},
      {stage1_10[55]}
   );
   gpc1_1 gpc328 (
      {stage0_10[159]},
      {stage1_10[56]}
   );
   gpc1_1 gpc329 (
      {stage0_10[160]},
      {stage1_10[57]}
   );
   gpc1_1 gpc330 (
      {stage0_10[161]},
      {stage1_10[58]}
   );
   gpc1163_5 gpc331 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc332 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc333 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc334 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc335 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc336 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc337 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc606_5 gpc338 (
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc339 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc606_5 gpc340 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc606_5 gpc341 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc606_5 gpc342 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc606_5 gpc343 (
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc344 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52]},
      {stage1_3[6]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc345 (
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[8],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc346 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[9],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc347 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[50]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[10],stage2_5[10],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc348 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[51]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[11],stage2_5[11],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc349 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[52]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[12],stage2_5[12],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc350 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[53]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[13],stage2_5[13],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc351 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[54]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[14],stage2_5[14],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc352 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[55]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[15],stage2_5[15],stage2_4[21],stage2_3[21]}
   );
   gpc606_5 gpc353 (
      {stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[8],stage2_6[16],stage2_5[16],stage2_4[22]}
   );
   gpc606_5 gpc354 (
      {stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[9],stage2_6[17],stage2_5[17],stage2_4[23]}
   );
   gpc606_5 gpc355 (
      {stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[10],stage2_6[18],stage2_5[18],stage2_4[24]}
   );
   gpc606_5 gpc356 (
      {stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77], stage1_4[78], stage1_4[79]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[11],stage2_6[19],stage2_5[19],stage2_4[25]}
   );
   gpc606_5 gpc357 (
      {stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[12],stage2_6[20],stage2_5[20],stage2_4[26]}
   );
   gpc606_5 gpc358 (
      {stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[13],stage2_6[21],stage2_5[21],stage2_4[27]}
   );
   gpc606_5 gpc359 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[14],stage2_6[22],stage2_5[22],stage2_4[28]}
   );
   gpc606_5 gpc360 (
      {stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[15],stage2_6[23],stage2_5[23],stage2_4[29]}
   );
   gpc606_5 gpc361 (
      {stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[16],stage2_6[24],stage2_5[24],stage2_4[30]}
   );
   gpc606_5 gpc362 (
      {stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[17],stage2_6[25],stage2_5[25],stage2_4[31]}
   );
   gpc606_5 gpc363 (
      {stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[18],stage2_6[26],stage2_5[26],stage2_4[32]}
   );
   gpc606_5 gpc364 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126], stage1_4[127]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[19],stage2_6[27],stage2_5[27],stage2_4[33]}
   );
   gpc606_5 gpc365 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[12],stage2_7[20],stage2_6[28],stage2_5[28]}
   );
   gpc606_5 gpc366 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[13],stage2_7[21],stage2_6[29],stage2_5[29]}
   );
   gpc615_5 gpc367 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76]},
      {stage1_7[12]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[14],stage2_7[22],stage2_6[30]}
   );
   gpc615_5 gpc368 (
      {stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[15],stage2_7[23],stage2_6[31]}
   );
   gpc615_5 gpc369 (
      {stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85], stage1_6[86]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[16],stage2_7[24],stage2_6[32]}
   );
   gpc615_5 gpc370 (
      {stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90], stage1_6[91]},
      {stage1_7[15]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[5],stage2_8[17],stage2_7[25],stage2_6[33]}
   );
   gpc615_5 gpc371 (
      {stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage1_7[16]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[6],stage2_8[18],stage2_7[26],stage2_6[34]}
   );
   gpc615_5 gpc372 (
      {stage1_7[17], stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21]},
      {stage1_8[30]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[7],stage2_8[19],stage2_7[27]}
   );
   gpc615_5 gpc373 (
      {stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26]},
      {stage1_8[31]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[8],stage2_8[20],stage2_7[28]}
   );
   gpc615_5 gpc374 (
      {stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31]},
      {stage1_8[32]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[9],stage2_8[21],stage2_7[29]}
   );
   gpc615_5 gpc375 (
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage1_8[33]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[10],stage2_8[22],stage2_7[30]}
   );
   gpc615_5 gpc376 (
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_8[34]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[11],stage2_8[23],stage2_7[31]}
   );
   gpc615_5 gpc377 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_8[35]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[12],stage2_8[24],stage2_7[32]}
   );
   gpc606_5 gpc378 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[6],stage2_10[11],stage2_9[13],stage2_8[25]}
   );
   gpc606_5 gpc379 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[7],stage2_10[12],stage2_9[14],stage2_8[26]}
   );
   gpc606_5 gpc380 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[8],stage2_10[13],stage2_9[15],stage2_8[27]}
   );
   gpc606_5 gpc381 (
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[9],stage2_10[14],stage2_9[16],stage2_8[28]}
   );
   gpc606_5 gpc382 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[4],stage2_11[10],stage2_10[15],stage2_9[17]}
   );
   gpc606_5 gpc383 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[5],stage2_11[11],stage2_10[16],stage2_9[18]}
   );
   gpc606_5 gpc384 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[6],stage2_11[12],stage2_10[17],stage2_9[19]}
   );
   gpc606_5 gpc385 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[7],stage2_11[13],stage2_10[18],stage2_9[20]}
   );
   gpc606_5 gpc386 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[8],stage2_11[14],stage2_10[19],stage2_9[21]}
   );
   gpc606_5 gpc387 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[9],stage2_11[15],stage2_10[20],stage2_9[22]}
   );
   gpc606_5 gpc388 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[6],stage2_12[10],stage2_11[16],stage2_10[21]}
   );
   gpc606_5 gpc389 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[7],stage2_12[11],stage2_11[17],stage2_10[22]}
   );
   gpc615_5 gpc390 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40]},
      {stage1_11[36]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[8],stage2_12[12],stage2_11[18],stage2_10[23]}
   );
   gpc615_5 gpc391 (
      {stage1_10[41], stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45]},
      {stage1_11[37]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[9],stage2_12[13],stage2_11[19],stage2_10[24]}
   );
   gpc615_5 gpc392 (
      {stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_11[38]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[10],stage2_12[14],stage2_11[20],stage2_10[25]}
   );
   gpc615_5 gpc393 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55]},
      {stage1_11[39]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[11],stage2_12[15],stage2_11[21],stage2_10[26]}
   );
   gpc1163_5 gpc394 (
      {stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[0]},
      {1'b0},
      {stage2_15[0],stage2_14[6],stage2_13[12],stage2_12[16],stage2_11[22]}
   );
   gpc615_5 gpc395 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage1_12[42]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[1],stage2_14[7],stage2_13[13],stage2_12[17],stage2_11[23]}
   );
   gpc615_5 gpc396 (
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52]},
      {stage1_12[43]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12]},
      {stage2_15[2],stage2_14[8],stage2_13[14],stage2_12[18],stage2_11[24]}
   );
   gpc1_1 gpc397 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc398 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc399 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc400 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc401 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc402 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc403 (
      {stage1_0[24]},
      {stage2_0[12]}
   );
   gpc1_1 gpc404 (
      {stage1_0[25]},
      {stage2_0[13]}
   );
   gpc1_1 gpc405 (
      {stage1_0[26]},
      {stage2_0[14]}
   );
   gpc1_1 gpc406 (
      {stage1_0[27]},
      {stage2_0[15]}
   );
   gpc1_1 gpc407 (
      {stage1_0[28]},
      {stage2_0[16]}
   );
   gpc1_1 gpc408 (
      {stage1_0[29]},
      {stage2_0[17]}
   );
   gpc1_1 gpc409 (
      {stage1_0[30]},
      {stage2_0[18]}
   );
   gpc1_1 gpc410 (
      {stage1_1[36]},
      {stage2_1[6]}
   );
   gpc1_1 gpc411 (
      {stage1_1[37]},
      {stage2_1[7]}
   );
   gpc1_1 gpc412 (
      {stage1_1[38]},
      {stage2_1[8]}
   );
   gpc1_1 gpc413 (
      {stage1_1[39]},
      {stage2_1[9]}
   );
   gpc1_1 gpc414 (
      {stage1_1[40]},
      {stage2_1[10]}
   );
   gpc1_1 gpc415 (
      {stage1_1[41]},
      {stage2_1[11]}
   );
   gpc1_1 gpc416 (
      {stage1_1[42]},
      {stage2_1[12]}
   );
   gpc1_1 gpc417 (
      {stage1_1[43]},
      {stage2_1[13]}
   );
   gpc1_1 gpc418 (
      {stage1_1[44]},
      {stage2_1[14]}
   );
   gpc1_1 gpc419 (
      {stage1_1[45]},
      {stage2_1[15]}
   );
   gpc1_1 gpc420 (
      {stage1_1[46]},
      {stage2_1[16]}
   );
   gpc1_1 gpc421 (
      {stage1_1[47]},
      {stage2_1[17]}
   );
   gpc1_1 gpc422 (
      {stage1_1[48]},
      {stage2_1[18]}
   );
   gpc1_1 gpc423 (
      {stage1_1[49]},
      {stage2_1[19]}
   );
   gpc1_1 gpc424 (
      {stage1_1[50]},
      {stage2_1[20]}
   );
   gpc1_1 gpc425 (
      {stage1_1[51]},
      {stage2_1[21]}
   );
   gpc1_1 gpc426 (
      {stage1_1[52]},
      {stage2_1[22]}
   );
   gpc1_1 gpc427 (
      {stage1_2[53]},
      {stage2_2[14]}
   );
   gpc1_1 gpc428 (
      {stage1_2[54]},
      {stage2_2[15]}
   );
   gpc1_1 gpc429 (
      {stage1_2[55]},
      {stage2_2[16]}
   );
   gpc1_1 gpc430 (
      {stage1_2[56]},
      {stage2_2[17]}
   );
   gpc1_1 gpc431 (
      {stage1_2[57]},
      {stage2_2[18]}
   );
   gpc1_1 gpc432 (
      {stage1_2[58]},
      {stage2_2[19]}
   );
   gpc1_1 gpc433 (
      {stage1_2[59]},
      {stage2_2[20]}
   );
   gpc1_1 gpc434 (
      {stage1_2[60]},
      {stage2_2[21]}
   );
   gpc1_1 gpc435 (
      {stage1_2[61]},
      {stage2_2[22]}
   );
   gpc1_1 gpc436 (
      {stage1_2[62]},
      {stage2_2[23]}
   );
   gpc1_1 gpc437 (
      {stage1_2[63]},
      {stage2_2[24]}
   );
   gpc1_1 gpc438 (
      {stage1_2[64]},
      {stage2_2[25]}
   );
   gpc1_1 gpc439 (
      {stage1_2[65]},
      {stage2_2[26]}
   );
   gpc1_1 gpc440 (
      {stage1_3[47]},
      {stage2_3[22]}
   );
   gpc1_1 gpc441 (
      {stage1_3[48]},
      {stage2_3[23]}
   );
   gpc1_1 gpc442 (
      {stage1_3[49]},
      {stage2_3[24]}
   );
   gpc1_1 gpc443 (
      {stage1_3[50]},
      {stage2_3[25]}
   );
   gpc1_1 gpc444 (
      {stage1_3[51]},
      {stage2_3[26]}
   );
   gpc1_1 gpc445 (
      {stage1_3[52]},
      {stage2_3[27]}
   );
   gpc1_1 gpc446 (
      {stage1_3[53]},
      {stage2_3[28]}
   );
   gpc1_1 gpc447 (
      {stage1_3[54]},
      {stage2_3[29]}
   );
   gpc1_1 gpc448 (
      {stage1_3[55]},
      {stage2_3[30]}
   );
   gpc1_1 gpc449 (
      {stage1_3[56]},
      {stage2_3[31]}
   );
   gpc1_1 gpc450 (
      {stage1_3[57]},
      {stage2_3[32]}
   );
   gpc1_1 gpc451 (
      {stage1_4[128]},
      {stage2_4[34]}
   );
   gpc1_1 gpc452 (
      {stage1_4[129]},
      {stage2_4[35]}
   );
   gpc1_1 gpc453 (
      {stage1_4[130]},
      {stage2_4[36]}
   );
   gpc1_1 gpc454 (
      {stage1_4[131]},
      {stage2_4[37]}
   );
   gpc1_1 gpc455 (
      {stage1_4[132]},
      {stage2_4[38]}
   );
   gpc1_1 gpc456 (
      {stage1_4[133]},
      {stage2_4[39]}
   );
   gpc1_1 gpc457 (
      {stage1_4[134]},
      {stage2_4[40]}
   );
   gpc1_1 gpc458 (
      {stage1_4[135]},
      {stage2_4[41]}
   );
   gpc1_1 gpc459 (
      {stage1_4[136]},
      {stage2_4[42]}
   );
   gpc1_1 gpc460 (
      {stage1_4[137]},
      {stage2_4[43]}
   );
   gpc1_1 gpc461 (
      {stage1_4[138]},
      {stage2_4[44]}
   );
   gpc1_1 gpc462 (
      {stage1_5[60]},
      {stage2_5[30]}
   );
   gpc1_1 gpc463 (
      {stage1_5[61]},
      {stage2_5[31]}
   );
   gpc1_1 gpc464 (
      {stage1_5[62]},
      {stage2_5[32]}
   );
   gpc1_1 gpc465 (
      {stage1_5[63]},
      {stage2_5[33]}
   );
   gpc1_1 gpc466 (
      {stage1_5[64]},
      {stage2_5[34]}
   );
   gpc1_1 gpc467 (
      {stage1_5[65]},
      {stage2_5[35]}
   );
   gpc1_1 gpc468 (
      {stage1_5[66]},
      {stage2_5[36]}
   );
   gpc1_1 gpc469 (
      {stage1_5[67]},
      {stage2_5[37]}
   );
   gpc1_1 gpc470 (
      {stage1_6[97]},
      {stage2_6[35]}
   );
   gpc1_1 gpc471 (
      {stage1_6[98]},
      {stage2_6[36]}
   );
   gpc1_1 gpc472 (
      {stage1_6[99]},
      {stage2_6[37]}
   );
   gpc1_1 gpc473 (
      {stage1_6[100]},
      {stage2_6[38]}
   );
   gpc1_1 gpc474 (
      {stage1_6[101]},
      {stage2_6[39]}
   );
   gpc1_1 gpc475 (
      {stage1_6[102]},
      {stage2_6[40]}
   );
   gpc1_1 gpc476 (
      {stage1_6[103]},
      {stage2_6[41]}
   );
   gpc1_1 gpc477 (
      {stage1_6[104]},
      {stage2_6[42]}
   );
   gpc1_1 gpc478 (
      {stage1_6[105]},
      {stage2_6[43]}
   );
   gpc1_1 gpc479 (
      {stage1_6[106]},
      {stage2_6[44]}
   );
   gpc1_1 gpc480 (
      {stage1_6[107]},
      {stage2_6[45]}
   );
   gpc1_1 gpc481 (
      {stage1_6[108]},
      {stage2_6[46]}
   );
   gpc1_1 gpc482 (
      {stage1_6[109]},
      {stage2_6[47]}
   );
   gpc1_1 gpc483 (
      {stage1_6[110]},
      {stage2_6[48]}
   );
   gpc1_1 gpc484 (
      {stage1_6[111]},
      {stage2_6[49]}
   );
   gpc1_1 gpc485 (
      {stage1_7[47]},
      {stage2_7[33]}
   );
   gpc1_1 gpc486 (
      {stage1_8[60]},
      {stage2_8[29]}
   );
   gpc1_1 gpc487 (
      {stage1_8[61]},
      {stage2_8[30]}
   );
   gpc1_1 gpc488 (
      {stage1_8[62]},
      {stage2_8[31]}
   );
   gpc1_1 gpc489 (
      {stage1_8[63]},
      {stage2_8[32]}
   );
   gpc1_1 gpc490 (
      {stage1_8[64]},
      {stage2_8[33]}
   );
   gpc1_1 gpc491 (
      {stage1_8[65]},
      {stage2_8[34]}
   );
   gpc1_1 gpc492 (
      {stage1_8[66]},
      {stage2_8[35]}
   );
   gpc1_1 gpc493 (
      {stage1_8[67]},
      {stage2_8[36]}
   );
   gpc1_1 gpc494 (
      {stage1_8[68]},
      {stage2_8[37]}
   );
   gpc1_1 gpc495 (
      {stage1_8[69]},
      {stage2_8[38]}
   );
   gpc1_1 gpc496 (
      {stage1_8[70]},
      {stage2_8[39]}
   );
   gpc1_1 gpc497 (
      {stage1_8[71]},
      {stage2_8[40]}
   );
   gpc1_1 gpc498 (
      {stage1_8[72]},
      {stage2_8[41]}
   );
   gpc1_1 gpc499 (
      {stage1_9[72]},
      {stage2_9[23]}
   );
   gpc1_1 gpc500 (
      {stage1_9[73]},
      {stage2_9[24]}
   );
   gpc1_1 gpc501 (
      {stage1_9[74]},
      {stage2_9[25]}
   );
   gpc1_1 gpc502 (
      {stage1_9[75]},
      {stage2_9[26]}
   );
   gpc1_1 gpc503 (
      {stage1_9[76]},
      {stage2_9[27]}
   );
   gpc1_1 gpc504 (
      {stage1_9[77]},
      {stage2_9[28]}
   );
   gpc1_1 gpc505 (
      {stage1_9[78]},
      {stage2_9[29]}
   );
   gpc1_1 gpc506 (
      {stage1_10[56]},
      {stage2_10[27]}
   );
   gpc1_1 gpc507 (
      {stage1_10[57]},
      {stage2_10[28]}
   );
   gpc1_1 gpc508 (
      {stage1_10[58]},
      {stage2_10[29]}
   );
   gpc1_1 gpc509 (
      {stage1_12[44]},
      {stage2_12[19]}
   );
   gpc1_1 gpc510 (
      {stage1_12[45]},
      {stage2_12[20]}
   );
   gpc1_1 gpc511 (
      {stage1_12[46]},
      {stage2_12[21]}
   );
   gpc1_1 gpc512 (
      {stage1_12[47]},
      {stage2_12[22]}
   );
   gpc1_1 gpc513 (
      {stage1_12[48]},
      {stage2_12[23]}
   );
   gpc1_1 gpc514 (
      {stage1_12[49]},
      {stage2_12[24]}
   );
   gpc1_1 gpc515 (
      {stage1_12[50]},
      {stage2_12[25]}
   );
   gpc1_1 gpc516 (
      {stage1_12[51]},
      {stage2_12[26]}
   );
   gpc1_1 gpc517 (
      {stage1_12[52]},
      {stage2_12[27]}
   );
   gpc1_1 gpc518 (
      {stage1_13[13]},
      {stage2_13[15]}
   );
   gpc1_1 gpc519 (
      {stage1_13[14]},
      {stage2_13[16]}
   );
   gpc1_1 gpc520 (
      {stage1_13[15]},
      {stage2_13[17]}
   );
   gpc1_1 gpc521 (
      {stage1_13[16]},
      {stage2_13[18]}
   );
   gpc1_1 gpc522 (
      {stage1_13[17]},
      {stage2_13[19]}
   );
   gpc1_1 gpc523 (
      {stage1_13[18]},
      {stage2_13[20]}
   );
   gpc1_1 gpc524 (
      {stage1_13[19]},
      {stage2_13[21]}
   );
   gpc1_1 gpc525 (
      {stage1_13[20]},
      {stage2_13[22]}
   );
   gpc1_1 gpc526 (
      {stage1_13[21]},
      {stage2_13[23]}
   );
   gpc1_1 gpc527 (
      {stage1_13[22]},
      {stage2_13[24]}
   );
   gpc1_1 gpc528 (
      {stage1_13[23]},
      {stage2_13[25]}
   );
   gpc1_1 gpc529 (
      {stage1_13[24]},
      {stage2_13[26]}
   );
   gpc1_1 gpc530 (
      {stage1_13[25]},
      {stage2_13[27]}
   );
   gpc1_1 gpc531 (
      {stage1_13[26]},
      {stage2_13[28]}
   );
   gpc1163_5 gpc532 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc533 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1406_5 gpc534 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc615_5 gpc535 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_3[5]},
      {stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc536 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc537 (
      {stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage2_4[8]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc538 (
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20]},
      {stage2_4[9]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc615_5 gpc539 (
      {stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25]},
      {stage2_4[10]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[7],stage3_3[7]}
   );
   gpc606_5 gpc540 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc541 (
      {stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc542 (
      {stage2_4[23], stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[6],stage3_6[7],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc543 (
      {stage2_4[29], stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33]},
      {stage2_5[24]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[7],stage3_6[8],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc544 (
      {stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37], stage2_4[38]},
      {stage2_5[25]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[8],stage3_6[9],stage3_5[10],stage3_4[12]}
   );
   gpc606_5 gpc545 (
      {stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29], stage2_5[30], stage2_5[31]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[5],stage3_7[9],stage3_6[10],stage3_5[11]}
   );
   gpc606_5 gpc546 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[6],stage3_7[10],stage3_6[11]}
   );
   gpc615_5 gpc547 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[6]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[7],stage3_7[11],stage3_6[12]}
   );
   gpc615_5 gpc548 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[7]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[3],stage3_8[8],stage3_7[12],stage3_6[13]}
   );
   gpc1343_5 gpc549 (
      {stage2_7[8], stage2_7[9], stage2_7[10]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[0]},
      {stage3_11[0],stage3_10[3],stage3_9[4],stage3_8[9],stage3_7[13]}
   );
   gpc1343_5 gpc550 (
      {stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[1]},
      {stage3_11[1],stage3_10[4],stage3_9[5],stage3_8[10],stage3_7[14]}
   );
   gpc615_5 gpc551 (
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_8[26]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[2],stage3_10[5],stage3_9[6],stage3_8[11],stage3_7[15]}
   );
   gpc615_5 gpc552 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[27]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[3],stage3_10[6],stage3_9[7],stage3_8[12],stage3_7[16]}
   );
   gpc615_5 gpc553 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[28]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[4],stage3_10[7],stage3_9[8],stage3_8[13],stage3_7[17]}
   );
   gpc615_5 gpc554 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[29]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[5],stage3_10[8],stage3_9[9],stage3_8[14],stage3_7[18]}
   );
   gpc606_5 gpc555 (
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6], stage2_10[7]},
      {stage3_12[0],stage3_11[6],stage3_10[9],stage3_9[10],stage3_8[15]}
   );
   gpc606_5 gpc556 (
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12], stage2_10[13]},
      {stage3_12[1],stage3_11[7],stage3_10[10],stage3_9[11],stage3_8[16]}
   );
   gpc606_5 gpc557 (
      {stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[8],stage3_10[11]}
   );
   gpc615_5 gpc558 (
      {stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24]},
      {stage2_11[0]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[9],stage3_10[12]}
   );
   gpc615_5 gpc559 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_11[1]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[10],stage3_10[13]}
   );
   gpc615_5 gpc560 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_12[18]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[11]}
   );
   gpc615_5 gpc561 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[19]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[12]}
   );
   gpc615_5 gpc562 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[20]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[5],stage3_12[7],stage3_11[13]}
   );
   gpc615_5 gpc563 (
      {stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage2_12[21]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[6],stage3_12[8],stage3_11[14]}
   );
   gpc606_5 gpc564 (
      {stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[4],stage3_14[7],stage3_13[7],stage3_12[9]}
   );
   gpc1_1 gpc565 (
      {stage2_0[9]},
      {stage3_0[2]}
   );
   gpc1_1 gpc566 (
      {stage2_0[10]},
      {stage3_0[3]}
   );
   gpc1_1 gpc567 (
      {stage2_0[11]},
      {stage3_0[4]}
   );
   gpc1_1 gpc568 (
      {stage2_0[12]},
      {stage3_0[5]}
   );
   gpc1_1 gpc569 (
      {stage2_0[13]},
      {stage3_0[6]}
   );
   gpc1_1 gpc570 (
      {stage2_0[14]},
      {stage3_0[7]}
   );
   gpc1_1 gpc571 (
      {stage2_0[15]},
      {stage3_0[8]}
   );
   gpc1_1 gpc572 (
      {stage2_0[16]},
      {stage3_0[9]}
   );
   gpc1_1 gpc573 (
      {stage2_0[17]},
      {stage3_0[10]}
   );
   gpc1_1 gpc574 (
      {stage2_0[18]},
      {stage3_0[11]}
   );
   gpc1_1 gpc575 (
      {stage2_1[12]},
      {stage3_1[3]}
   );
   gpc1_1 gpc576 (
      {stage2_1[13]},
      {stage3_1[4]}
   );
   gpc1_1 gpc577 (
      {stage2_1[14]},
      {stage3_1[5]}
   );
   gpc1_1 gpc578 (
      {stage2_1[15]},
      {stage3_1[6]}
   );
   gpc1_1 gpc579 (
      {stage2_1[16]},
      {stage3_1[7]}
   );
   gpc1_1 gpc580 (
      {stage2_1[17]},
      {stage3_1[8]}
   );
   gpc1_1 gpc581 (
      {stage2_1[18]},
      {stage3_1[9]}
   );
   gpc1_1 gpc582 (
      {stage2_1[19]},
      {stage3_1[10]}
   );
   gpc1_1 gpc583 (
      {stage2_1[20]},
      {stage3_1[11]}
   );
   gpc1_1 gpc584 (
      {stage2_1[21]},
      {stage3_1[12]}
   );
   gpc1_1 gpc585 (
      {stage2_1[22]},
      {stage3_1[13]}
   );
   gpc1_1 gpc586 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc587 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc588 (
      {stage2_2[14]},
      {stage3_2[6]}
   );
   gpc1_1 gpc589 (
      {stage2_2[15]},
      {stage3_2[7]}
   );
   gpc1_1 gpc590 (
      {stage2_2[16]},
      {stage3_2[8]}
   );
   gpc1_1 gpc591 (
      {stage2_2[17]},
      {stage3_2[9]}
   );
   gpc1_1 gpc592 (
      {stage2_2[18]},
      {stage3_2[10]}
   );
   gpc1_1 gpc593 (
      {stage2_2[19]},
      {stage3_2[11]}
   );
   gpc1_1 gpc594 (
      {stage2_2[20]},
      {stage3_2[12]}
   );
   gpc1_1 gpc595 (
      {stage2_2[21]},
      {stage3_2[13]}
   );
   gpc1_1 gpc596 (
      {stage2_2[22]},
      {stage3_2[14]}
   );
   gpc1_1 gpc597 (
      {stage2_2[23]},
      {stage3_2[15]}
   );
   gpc1_1 gpc598 (
      {stage2_2[24]},
      {stage3_2[16]}
   );
   gpc1_1 gpc599 (
      {stage2_2[25]},
      {stage3_2[17]}
   );
   gpc1_1 gpc600 (
      {stage2_2[26]},
      {stage3_2[18]}
   );
   gpc1_1 gpc601 (
      {stage2_3[26]},
      {stage3_3[8]}
   );
   gpc1_1 gpc602 (
      {stage2_3[27]},
      {stage3_3[9]}
   );
   gpc1_1 gpc603 (
      {stage2_3[28]},
      {stage3_3[10]}
   );
   gpc1_1 gpc604 (
      {stage2_3[29]},
      {stage3_3[11]}
   );
   gpc1_1 gpc605 (
      {stage2_3[30]},
      {stage3_3[12]}
   );
   gpc1_1 gpc606 (
      {stage2_3[31]},
      {stage3_3[13]}
   );
   gpc1_1 gpc607 (
      {stage2_3[32]},
      {stage3_3[14]}
   );
   gpc1_1 gpc608 (
      {stage2_4[39]},
      {stage3_4[13]}
   );
   gpc1_1 gpc609 (
      {stage2_4[40]},
      {stage3_4[14]}
   );
   gpc1_1 gpc610 (
      {stage2_4[41]},
      {stage3_4[15]}
   );
   gpc1_1 gpc611 (
      {stage2_4[42]},
      {stage3_4[16]}
   );
   gpc1_1 gpc612 (
      {stage2_4[43]},
      {stage3_4[17]}
   );
   gpc1_1 gpc613 (
      {stage2_4[44]},
      {stage3_4[18]}
   );
   gpc1_1 gpc614 (
      {stage2_5[32]},
      {stage3_5[12]}
   );
   gpc1_1 gpc615 (
      {stage2_5[33]},
      {stage3_5[13]}
   );
   gpc1_1 gpc616 (
      {stage2_5[34]},
      {stage3_5[14]}
   );
   gpc1_1 gpc617 (
      {stage2_5[35]},
      {stage3_5[15]}
   );
   gpc1_1 gpc618 (
      {stage2_5[36]},
      {stage3_5[16]}
   );
   gpc1_1 gpc619 (
      {stage2_5[37]},
      {stage3_5[17]}
   );
   gpc1_1 gpc620 (
      {stage2_6[46]},
      {stage3_6[14]}
   );
   gpc1_1 gpc621 (
      {stage2_6[47]},
      {stage3_6[15]}
   );
   gpc1_1 gpc622 (
      {stage2_6[48]},
      {stage3_6[16]}
   );
   gpc1_1 gpc623 (
      {stage2_6[49]},
      {stage3_6[17]}
   );
   gpc1_1 gpc624 (
      {stage2_11[22]},
      {stage3_11[15]}
   );
   gpc1_1 gpc625 (
      {stage2_11[23]},
      {stage3_11[16]}
   );
   gpc1_1 gpc626 (
      {stage2_11[24]},
      {stage3_11[17]}
   );
   gpc1_1 gpc627 (
      {stage2_13[24]},
      {stage3_13[8]}
   );
   gpc1_1 gpc628 (
      {stage2_13[25]},
      {stage3_13[9]}
   );
   gpc1_1 gpc629 (
      {stage2_13[26]},
      {stage3_13[10]}
   );
   gpc1_1 gpc630 (
      {stage2_13[27]},
      {stage3_13[11]}
   );
   gpc1_1 gpc631 (
      {stage2_13[28]},
      {stage3_13[12]}
   );
   gpc1_1 gpc632 (
      {stage2_14[6]},
      {stage3_14[8]}
   );
   gpc1_1 gpc633 (
      {stage2_14[7]},
      {stage3_14[9]}
   );
   gpc1_1 gpc634 (
      {stage2_14[8]},
      {stage3_14[10]}
   );
   gpc1_1 gpc635 (
      {stage2_15[0]},
      {stage3_15[5]}
   );
   gpc1_1 gpc636 (
      {stage2_15[1]},
      {stage3_15[6]}
   );
   gpc1_1 gpc637 (
      {stage2_15[2]},
      {stage3_15[7]}
   );
   gpc606_5 gpc638 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc639 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc640 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc641 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc642 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[3],stage4_4[4]}
   );
   gpc606_5 gpc643 (
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[4],stage4_4[5]}
   );
   gpc606_5 gpc644 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[3],stage4_7[3],stage4_6[3],stage4_5[5]}
   );
   gpc606_5 gpc645 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[4],stage4_7[4],stage4_6[4],stage4_5[6]}
   );
   gpc606_5 gpc646 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[5],stage4_7[5],stage4_6[5],stage4_5[7]}
   );
   gpc2135_5 gpc647 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[3],stage4_8[6]}
   );
   gpc2135_5 gpc648 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[1]},
      {stage3_11[2], stage3_11[3]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[4],stage4_8[7]}
   );
   gpc606_5 gpc649 (
      {stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[5],stage4_8[8]}
   );
   gpc606_5 gpc650 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage3_11[4], stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9]},
      {stage4_13[0],stage4_12[3],stage4_11[3],stage4_10[3],stage4_9[6]}
   );
   gpc1325_5 gpc651 (
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12]},
      {stage3_11[10], stage3_11[11]},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[1],stage4_12[4],stage4_11[4],stage4_10[4]}
   );
   gpc606_5 gpc652 (
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6]},
      {stage4_15[0],stage4_14[1],stage4_13[2],stage4_12[5],stage4_11[5]}
   );
   gpc615_5 gpc653 (
      {stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7]},
      {stage3_13[7]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[2],stage4_13[3],stage4_12[6]}
   );
   gpc606_5 gpc654 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], 1'b0},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[3],stage4_13[4]}
   );
   gpc1_1 gpc655 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc656 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc657 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc658 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc659 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc660 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc661 (
      {stage3_1[12]},
      {stage4_1[3]}
   );
   gpc1_1 gpc662 (
      {stage3_1[13]},
      {stage4_1[4]}
   );
   gpc1_1 gpc663 (
      {stage3_2[6]},
      {stage4_2[3]}
   );
   gpc1_1 gpc664 (
      {stage3_2[7]},
      {stage4_2[4]}
   );
   gpc1_1 gpc665 (
      {stage3_2[8]},
      {stage4_2[5]}
   );
   gpc1_1 gpc666 (
      {stage3_2[9]},
      {stage4_2[6]}
   );
   gpc1_1 gpc667 (
      {stage3_2[10]},
      {stage4_2[7]}
   );
   gpc1_1 gpc668 (
      {stage3_2[11]},
      {stage4_2[8]}
   );
   gpc1_1 gpc669 (
      {stage3_2[12]},
      {stage4_2[9]}
   );
   gpc1_1 gpc670 (
      {stage3_2[13]},
      {stage4_2[10]}
   );
   gpc1_1 gpc671 (
      {stage3_2[14]},
      {stage4_2[11]}
   );
   gpc1_1 gpc672 (
      {stage3_2[15]},
      {stage4_2[12]}
   );
   gpc1_1 gpc673 (
      {stage3_2[16]},
      {stage4_2[13]}
   );
   gpc1_1 gpc674 (
      {stage3_2[17]},
      {stage4_2[14]}
   );
   gpc1_1 gpc675 (
      {stage3_2[18]},
      {stage4_2[15]}
   );
   gpc1_1 gpc676 (
      {stage3_3[12]},
      {stage4_3[3]}
   );
   gpc1_1 gpc677 (
      {stage3_3[13]},
      {stage4_3[4]}
   );
   gpc1_1 gpc678 (
      {stage3_3[14]},
      {stage4_3[5]}
   );
   gpc1_1 gpc679 (
      {stage3_4[18]},
      {stage4_4[6]}
   );
   gpc1_1 gpc680 (
      {stage3_7[18]},
      {stage4_7[6]}
   );
   gpc1_1 gpc681 (
      {stage3_8[16]},
      {stage4_8[9]}
   );
   gpc1_1 gpc682 (
      {stage3_10[13]},
      {stage4_10[5]}
   );
   gpc1_1 gpc683 (
      {stage3_12[8]},
      {stage4_12[7]}
   );
   gpc1_1 gpc684 (
      {stage3_12[9]},
      {stage4_12[8]}
   );
   gpc1_1 gpc685 (
      {stage3_14[6]},
      {stage4_14[4]}
   );
   gpc1_1 gpc686 (
      {stage3_14[7]},
      {stage4_14[5]}
   );
   gpc1_1 gpc687 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc688 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc689 (
      {stage3_14[10]},
      {stage4_14[8]}
   );
   gpc1_1 gpc690 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc691 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc1_1 gpc692 (
      {stage3_16[0]},
      {stage4_16[2]}
   );
   gpc606_5 gpc693 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc1325_5 gpc694 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6], stage4_2[7]},
      {stage4_3[0], stage4_3[1], stage4_3[2]},
      {stage4_4[0]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc695 (
      {stage4_2[8], stage4_2[9], stage4_2[10], stage4_2[11], stage4_2[12], stage4_2[13]},
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6]},
      {stage5_6[0],stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2]}
   );
   gpc615_5 gpc696 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[2]}
   );
   gpc615_5 gpc697 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[2]}
   );
   gpc606_5 gpc698 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[2]}
   );
   gpc1406_5 gpc699 (
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[2]}
   );
   gpc2135_5 gpc700 (
      {stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8]},
      {stage4_13[1], stage4_13[2], stage4_13[3]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1]},
      {stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[2],stage5_12[2]}
   );
   gpc1406_5 gpc701 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5], stage4_14[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], 1'b0},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[2]}
   );
   gpc1_1 gpc702 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc703 (
      {stage4_2[14]},
      {stage5_2[3]}
   );
   gpc1_1 gpc704 (
      {stage4_2[15]},
      {stage5_2[4]}
   );
   gpc1_1 gpc705 (
      {stage4_3[3]},
      {stage5_3[3]}
   );
   gpc1_1 gpc706 (
      {stage4_3[4]},
      {stage5_3[4]}
   );
   gpc1_1 gpc707 (
      {stage4_3[5]},
      {stage5_3[5]}
   );
   gpc1_1 gpc708 (
      {stage4_5[5]},
      {stage5_5[3]}
   );
   gpc1_1 gpc709 (
      {stage4_5[6]},
      {stage5_5[4]}
   );
   gpc1_1 gpc710 (
      {stage4_5[7]},
      {stage5_5[5]}
   );
   gpc1_1 gpc711 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc712 (
      {stage4_8[7]},
      {stage5_8[3]}
   );
   gpc1_1 gpc713 (
      {stage4_8[8]},
      {stage5_8[4]}
   );
   gpc1_1 gpc714 (
      {stage4_8[9]},
      {stage5_8[5]}
   );
   gpc1_1 gpc715 (
      {stage4_9[6]},
      {stage5_9[3]}
   );
   gpc1_1 gpc716 (
      {stage4_13[4]},
      {stage5_13[3]}
   );
   gpc1_1 gpc717 (
      {stage4_14[7]},
      {stage5_14[3]}
   );
   gpc1_1 gpc718 (
      {stage4_14[8]},
      {stage5_14[4]}
   );
   gpc1_1 gpc719 (
      {stage4_15[2]},
      {stage5_15[2]}
   );
   gpc1_1 gpc720 (
      {stage4_15[3]},
      {stage5_15[3]}
   );
   gpc1_1 gpc721 (
      {stage4_15[4]},
      {stage5_15[4]}
   );
   gpc215_4 gpc722 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc615_5 gpc723 (
      {stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc623_5 gpc724 (
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0], stage5_7[1]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc2135_5 gpc725 (
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], 1'b0},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage5_12[0], stage5_12[1]},
      {stage6_13[0],stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1]}
   );
   gpc615_5 gpc726 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], 1'b0},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], 1'b0},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[1]}
   );
   gpc1325_5 gpc727 (
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], 1'b0},
      {1'b0, 1'b0},
      {stage5_16[0], stage5_16[1], 1'b0},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1],stage6_14[1]}
   );
   gpc1_1 gpc728 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc729 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc730 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc731 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc732 (
      {stage5_11[1]},
      {stage6_11[1]}
   );
   gpc1_1 gpc733 (
      {stage5_12[2]},
      {stage6_12[1]}
   );
   gpc1_1 gpc734 (
      {stage5_18[0]},
      {stage6_18[1]}
   );
endmodule
module rowadder2_1_19(input [18:0] src0, input [18:0] src1, output [19:0] dst0);
    wire [18:0] gene;
    wire [18:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({1'h0, gene[18:16]}),
        .S({1'h0, prop[18:16]})
    );
    assign dst0 = {carryout[18], out[18:0]};
endmodule


module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor2_1_162_12 compressor2_1_162_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2e82f9807b32db4ec99f59299d768d071a339c346c4277a7cbc7e8be89ea339eb5795b8ecf03f94c107cb7c38c6c17537bb4a18535536049f9bcede185b8f40cf3366e969f92a7ec18a8194303614aef3e4ee9c6f1cf9951eeeea7e411345eb4956c1e4677e7b255e477ea25962b0fb214c9a1cae70159a295d0d41efad0d38be292550d92592ef71abca29b3256711307fbee39e4128181695b9edfba251a9445132b85ce4a305d559c15ead269e2d7af7350cbb748fddcabef5525da5c5e3a639c042281af77e07e5fa3c64036c6e86db7dc18a248eb0c1e6f6f769248c1ae4c74e5dc0e70a4589f8097c233c8b9db5f2565;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfc1e7fcc5a46d5b3b55eba5909e0e02b8b4b475d5ca8f91d0e22ad5b94905a7395da3889459db192c434183adf567ef9e3436f994e6872a21e2145f45855eae81d30a2f3eb55ce1764a0d43293c4bf1e33c48e509210b4648e3dec80a67796e96e3ecce6df2ed7a6039f62bbc29be95f052175b045d2d02fa1e7c4ba038de5e5e98665d7a144edad1adaf9dc1b2b59489cd8fc57a2d361def57e008c306f234fe78aa7b6514701806642169d5dc0996ba94a5c039be4c3395eae4d8e656e968e524082569359320a709772d0ae22090bfb5ec9a5699f76e8572d96173d910ed5e2cc07ed83aeab120691066458e83e72912da6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hae069acde2dadb0ce7a288bc73fc5ee16d3cd31114d643a37c8f9aff8ff8d5af29caac4b32e60ed61f43b005747c2236d09c3395d6d291823d57ff710beea31937abc6adacb5e6f69d4aa68ad62924c86606c9bcb986de98343c03b304fa272fcdac529cfa6757c534757752e5bf6fce64e453c9888dff9066c137fbd7775739e7eaea502cc0178987ce985b19e38f3168b5ca0ef4345580c87ea912cbe589b2f761ce7ad666b74aa7423e85f0e7ec3a6eb8bb2ba023e2733d87a3cab622f832690c580da77e021155b3fab48189fcabd8d0a0c6c01bc387fa0aa12919a1f0b7cdda97e2ac3802dc98f09a46644475b6dde58c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2b12550f8123e91e711d694dca972b6999bd9b89da3f14b1cf876ac9041df563225e3fd7182d1697ce9818e0add4d36f875e50ff00c3df379a96ee9c18608d1b5983fbe71d342c82f27c846171736a03caa3151f342d44cc1ccf43e40b32680d3fc006a99d8ba63554720f973fb6fc3643f7dbcdf3f7dbbe7840231ed4367da489946a7512adccd7e95ea14caf73d7f0a70f1792a624c165b430730720101c6b109d40d14db1307ef53707383630331b67366a7ac605022707c9f7a5c423e0bd25b1b87f61365456cf54d7593dd45b8a1fea61e91d0bc33552d40d770565f3e55656e0b255f370f2bce886cc3b47cd2b33a099;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h6b34463db299f77cc9a730eb5f45d203f5c25fce1680076af86303d117068e97ddaf520d48e3237e755c09ff74fa337e54cbeb8773eded7c4b06c96f1446b6ab229402fb69223cb918b7fb7fbe72477befde448e55c844f5d875ce7e9de7736f90a6d53390fb1de9843f5c0b737bb095ef008f12c12b9de5fa1b755daed86ee64350188f7a4baeab66ca6ea03ca8c0f2332e0fa56c1894a59d55d5bfa6c0e711e0279ce133d686c48d99c8b5e73093d8c20d321fcff6371d29ca6d780b95c781240468800cef6e6a825d3c8d1aef4e9d6a85c8d4d8c2d9eab15471ef370f7c15f055a06683881ec2ad238902e0ae360bb2c8e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4b49b200a7bf0a45738e21fea836523258c9dfbd02069ab80c4011c4d72c6e7a2f8b927d919884cfc1ae2931649d59e90e3cc62bf1399791ca4db56006fc707239134813540b9862ef9198eb15f407a5bd5c768d1ed4518ba4ccf57b17c46ded97f5b47f4e4f12564b75e9d068dc4c82fdc1585114674643d87cecac21caedd79cc27c8b3c798c448fdf461dcbdf76f70862ee2f98c011a0eb8e7f8e623e43835bcf73665b1a6211260c014116a9354f313a5a1112cc906dc5cada9147e342c9a237b5a9669640bfd015aa300d7c093ecf491cb04004fcaa7899681c62bfc6527c3cbbe66ec139519206c64d5f18add4dca72a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5464f4cfbb01bfa69987037075faa18688866a76fec731ccc3528e3a2a8b329c926218483399d1ee7d7e5afe694a0388be8fc9b531e32444c150e63d48937886694b051ecb56c0acf7c4d6505dd41f5c414dfbe370bf00f03b078337b06c255f6ad2e7fff43a3984500683c902cbe2f6a6e156e9954caf108b77aecf907f4a0d73a0a93e8266aabe55bf2311f0e929ee6e292037272d364346ff688e7b851e6d388c4700936109e63c806d5ee7a5718dc04d09104cef91bfe040d4f47850a400e1d272de64ab7afc3fce4f982f9b9e4bf619dc66951a00ad4aa778e1b4b8372a553abba698ccd429da81d8fda7cccc25bb018a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5ce1d5343288a94fbd02ff22b9da305346c96a3387f04a65259e18b2f341b55d0846d17476e9554c171bc7a4f2cf4f27885fc71bc5a1f762f8355048c0dfad818a0549eb4b45d3bb3daa3d7ea00cfc6f7439017f08448c7262dceba567fdf2739c5b6b8b74cafdf836bfa310d5722fe044687d6c51d3e0a0b0f4b1e7c4dee37ae2e7de9fc070b509e0beca459ac9d70170c2786324135042368f66777775c6560c08bf941c5672da57b427ed94b51e38fe17954990d9196a56edd723ab71043d41bd0925a8fbd95e0d2cf771aaac2d9dbaa2ae3b328246d341bcca6ea4bb76c95d0dcb2962d1b5a7bda35c5d5a8cb022a288d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h996484bcaeb1a05e614256535073dcaa8aa4e57672b332000e17ca5af2b21e4e0c928faca0d2defc971f9b17d101ee609beee2c42282859049aa651f8fdba9fffd7676e7ae4895f346375abcd269d9b2a594b0447fdfc6670f678ecfeb33da904d76bb6c52c2e7e3909484b824d236bf9e605d4d0ee839dcead1882a3a80a2f1973fc3b3068d1086545d252974b8195733a18dee55d3758b766444a4b015fc495eebbe1a208bf9ec1f970e5f40540bf89fb54e53d5bd2cc6f68c8e0a103cea945479ce74f0bae21bde1b54fe75a6abfcbb52b0469ceb044ea1dcbadfcbd9b4a6dadc05dd45c559afd71ce72913aeeba9a5c32b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hce4f470decb83b542febce569eddb081a31d4bac3ce392c03bfb48e8b7263d8fb007a919dfd698230f5c1bebf8e201766b5c69246a375238a6ce402cbd5a8faa098acc48afa5112d91d97d5171d2bb7ad37877d908ca3794354445b8cc2315327bce05f26226d086773b23c3327c6b65d61b2b03c70fec94f0d896fa382e948a2110a086ab6dfc833121d9c7904ffdb0cc3df572076272cb9ebcbd4116297f7713867e0e364f3d93537e2a837d5245deb28d103b167f2d52e9e44033a1ab5039f8b8a356d6174679db121367f0df6cd145d21c488aa26d811c58d398860e5c1e549b766448dd3eae610e52b0229b58c23ded7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hbfafd5e528b5ba79a18f8a2f0d9f343ff4f1f44ccf5030e565bbbfd2b2223efd9ce568c91ce9ebb27802b618343a0525bfa431814c078dba09dd6e02db7742d06488f28f5b70c7a91be3ea76d57fdd212d74bcb8bb077a62b83fc7ec761adff493c8b3aa3802bdd0b874eff3f0ff3650e302422cc49fac4adfed2afdd19573a1f3c4c4380529d3db4baeebab42a12fac86a1a5fb873244de64d1b0100aceb3c41eebc9c433916bd7bd983e7b02ec4b23e61dab979aa5dcdf79b4a416b69b44a8c53d87de89a28c7857de14d80ed5a8f31b6fbd2b28845ccd8701dd31c8e5ab9b6f28a1d9f58c6264388b0fae6ff4605d8ffc29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h283ca915e410e67a07cd542ed43103bbc2f439abcadfe519a5aab918e6efaac0df53c1ac445c8fdf952c80cf35844b16a1e0d1b779ddb52e3e662f3106a703dba57b7d61af3c45803557c4f4f366a0dab3885d1e0bef6e0aee1fe6523caa1092e2934abfd8e0bb060f45e04b7627120c09eed65fbf85c20c2278a7a0f517edd26800ef3c81ed517eec3088b59098d5c0f45328fffe5b38876cf67686f4e86d58dd13bc3c235d41d98be596da51d5abf5ece40128ad9f3de4cc101b7649aef88d1a830e9b8bbfb7ba73cafa77b0f59bd8ce40360c53ac99993b5e97a0e085eb3b7f409afae0c8e65ca8091cd998162dfe4aed12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h75cc126adab2a4e38397cf4be66b32b4834020d25edf4d4735136f71ec85e44d3aebd58ce51f65402c41c4fe18d2b0e52f0b34d5fc4611a6a6a28130f92260ccbcefdc14a0bdc872168bacc02f863c4f37c2a627849cdd37f537a5a14c1a03e54b26a9237d394cb251fa0ee0e31f0462585345c4891c4e7c66b2e9beb286f109dbb1cb7ef6883e90729c769a76e55e1ad882d28da71565692ef35f74983080d6817790665cc6e78e3d8c113ded765fc79ede23d3075d216d64314716393a47424808481661db2006ab803cca784655f64bf79c8ef9489c60bc981596011d772acd81773e0020c5124671a0279b38de1815124f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h451d967d2005e9640e3e88ad0bc94caf4f824ab7ee40fbd087922148ee8324bf7faf90d163f8ef41c44fbb39225ef2fb8ff7bafaccd14c7b1f95d5f05d87e64478b915a35edfa317a5083359d231ce1c83cef84499e0da8f20f78d5dd3de3dc17a16caf293d5e7e03502b82562fcdea5a3a4faebf0435e548badda31b93da4872329c6303415450eac93a1c53aa3dbe2d2efcc492e86e23e9dacab03eda49f2fbf3b7fb66c981cd91e9194ee29293894f742c2bb611d5e113bdfea004fc3edd0f1a270fc4c1f79107b1de43a0eacc296ecd1d12a0ff3128af7d6db40d29032d1d73453fce3e544a1f861852067037759207254;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf496e858fe7e3f32678ff2a40409710a188a577c6e41495a5373bc183da3e45b4ada5e12aabed0a5771a6c3d57c75193bc9628ff807beb6ff6f8833940d7cb0229551626ab05cb00ce6b4871413a0fd5d0191899699139bee06592a6198d263fec93dff1348f842b3d593a7a91d06d1fb80ca5107d6586ca66f2d7f2adb0ff6c3c4eea5738d476c2a3fb621e50d425ba3fa4a4f19a6a09496cc7041b5ca9e16f4f01012c528f81cf8014de1755306af00f8f708efc5031360c867fec8484b00265eb5ba459e0d384e9d3815eb9787f343944c09f7f62fa3044c2ee2a1c1913db3557ac550c53a5636ad8bef7ba593d304a2350;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'haba02c749c64eed1408af74a1b47e04926e02fd24110895dbf6511c6d332d56db6dea10441e68744458b4580b3ffe109a4ba2488dea5a1acb3319d562b2f3e71349e325aa7d131a62ac65986ec5370fbe7f92932d007f698bb14186fa6b49cb5bab676ff9011720b5454f9bcf8cd9c6101ab5027b410a5f11b1d2701c1cad4deb149c9c559abc15256282bbed1eb5538bc7eb914b601433a9e87a0eb0b4ed2a4b93272c8db5eade1b88e75596294b455245ec22bca225634a1a331c47c2703916aa6ff905ee4c884ceffbe6ec8a86144917e17d1508a483d59b512fa94ddc1e6606eddd0e20768b7aad4f46d86d1478efb10e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd9b6d17549300c74fa46aa23717487ba735ec9067b23ff34a8e2161ef17e1cfbbfba575f08fc40388a4f1b81b91483906d86d53154050b9ea779a3d4b9d21767b303b17338343b5d4615afe185f3ff0bb263a19cd65c3782ab655cce399aafb69fd9743e3e26bd67c909cc87e6d6ee3f93c4354e58e1381c298430c57e6536dd82cba7ff89ed7bd76a4cb1ce397d22fec871a4e3ca0f8638737aeef5fbb572a083e874280daf9124b05df1e33ae073779088390f8299a26bd73d7a4210eae449aa11d6e1c971dc3169e5243d8f7ff009716a765ea5d3f2089e409bad3dd3c943fb5d489315313352b3c25fbee8a1722ce5c906;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3c3959bbff5f5b8f636a70d00be0a4be5585e6846bd501ee6839ca11e871967d003a7d779f7e08088a817cd26721db5fc221b4d8eb6b0cecd1279497f9adbca5b410299e96fea8df4b9bbe8b12a7b7428534deea2e120062dce657f5aaf6a2be02457f2098a7711dcea9e203f14dcca280c433b785651de09e140e17591189e016ecbbbf414e19cd2cc7ad70e08ca38547151d2e09fb82b88cc165dfc9dd6dacf048928913fd7354dea2066c26577ddc9d9739dc28a91c67933f267f97d8b2d317c53bb83ce1ac83ae5df9252127101923a8dd8537b42d6b5eaed0bfc1caa60cde607a010044dd2f8b7b85add46341d7be5be5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5982594c27dc51e180eff1d10b540c74f0589b681cb217c9d6bd5fff5978c70c7a82f1ed66d95eed7dc0c154de28f4f37212b761c29e3091ec390024a5a04f971975ec090a794e1a9d7dfc25017bc241c18cabdaca6f749e92b0dc635ba587c3efc0df8b3e51215f2c246a34b88c9c2b2c834a0a14d5df0a3cfbde22d6e0f53daed83099ee7d02b98e28c655dc741c6cdb669d51b3e8952b87e46280da31883c2a0baec2058e9947afd737727eaa97c8ad22953c8a1c5b6e007c193c9d285fc2d1000dccdde685b3d0d6d43b980866cdffb1e4cad9e21b26dcaba58d185cf1e74da07686bfa388e9c36a15e8e18c0025c3edaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h83506185e463e663e4bdd91287593156e07274c6ed8e886214d2699c6b12b5f89e5193d4517863b5a3b7b5f776166603b6441b9b79fce521d8d55276b2e24dd43dedcff1eac080897a7a7942bfefdf2837812391fd92ac583dd67e366df19e4e818ac7df0916cd43768819fb1109889ba3ca9db3ed26f938337c08a9ff362c5d0ae106d8c1a4c0df06eab4f3ef3e8c61457c8fb6f09a6eb803daae216ddeea81887206c788e6671d687d3e8ebe142846eb95fa87aec42319f5cba93359b712c7faa19f066cfdb682e2de1bea00a7204472d4f32b28566d1cfebe1958a8f77be27b225e2c12d27b17116531324b9fd510e8e1fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'heb50e6e42ab3bde603bfa1d8eeba1a497136ac8616fada91d50ebe91bf0787df67344ddac3ff731075fc11d9afc14bab2132c1afab25dbab8ad7d7aeaa9ed46bf152d19639862b5f10d70efb52d3addb966c3cda61239253cd4d43b2eaa272e3414dd925273cc69d4debff67605238d0860e3bce88aec39b3d29440450041a8496908264d450725be5119f0a28493d8cb7159ef10092d924eadd5e24804b5cef64d221dde1a3ce473ed9b7393223d9680d418b43e5bc0a5dec5dfbb53cd7e43bf531c5f509910ca0b344e2856b3414137569b858be8c1dedbf7083a3c2550de3271d01b7fe6685a462f5ad5a54ac1a6be7b3f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h8d3856db7c71e63628ebabbe44a9650c5cc05df87119c3b6cda8cedf5fa1bbb021fe24e9ff64f95e00f43f651850bbabe6373dd215f3f145b35a4a89e6360853c67133e0c7734768c456b9b6ae34cd1d845a2a7d6bfdacf473850d8a2ac22f67f72e054867a7a21dd77ae1be76c5c29e8ffcab068930cf851c0ce1acc00ce6a030580dcea28e3ee0747d6f168da6a05be34e7758d9177d4e0e8f21954d6c4f74a4bb2000175c00aa8f113edc73c557773fa0c18c0ab7acd875a2d6d7132ee34c94b4c60453599560decd09dd951c253fe4695e5f2d92678801436646517da441ceea1c091e3dd64165b3ea757511663a098424;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hff13a0052bd7dcc4d4d80c01df7bffd76798b4597d5cce10f51f3f536b6532fcd7302f65ad8648197992fef9d59dd29402d7185a21388c14288efcf9a7b4d37740e198c1c78221fa85d4cb7d4bef49f995eba43e72186e2f9ca259e1fbac3032bceed77913233af6277aa1f12500eb9d719fe8fa6e252fdf4e6660898c09346c3e4b27fcdcc151a844ed7effdb2b3c381822cc611e33023572a990a8cf629255c2a0f9e9a6b3bbf5473fe84376075735d0dc07e6ded4f55bc62502cab3080d4c30665b4746755803697d672e50660b5b2193adb82dcda9137440f029c58bdaf9961066989d04b11aaa7ce714581eaced1c5edd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h1d95ee8a05b2fbd280e46d16ef91ea00accac2b2bdd342cf125983712de60f330e02a71c27b83ae8aec2c1a20a9ae8664d82d265040a9ce3e0d5db6518b95da9e2e42f02999f5cb1c4876c6ddd295b05610e1fcdc212f4a085b0ac01d0d2cf32410903731a8e111e61e5902a11b82227e26d73c6a05f75c3a2b6ebcc35e24d83e164f81e108b637787c03251d6c83c69adcb76bd078fcbebc8b961cb8d956e3e729818287d4b50e82ded86cf7cbb31e05d6fc3bd1f8e71922d93dd3ba31738771c6b9f0738739c146a329f9daaeb66d7025dc465996e87903922d1af4e1999c20f9f8fc09afd8a4d411cb280776ac8a8edc41c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5eede761fbfe7a10093ac50bdea1862ec4633d5b6f4bcece239462cad6a31d7a82275624e6817cecfcc3db101dd8a97dbd64fc4a036b43b678675be1a01c819213173ed91270d7cb1679ea291bf1506c6943d5ff28a2da02f54d24de5744ea49a15ccbe4809b78a21b8567bde11a49f83c0b84688cec8380d66256a264421525295427bc32c6a6a636571e8f450d83baf9ccf2870c182dd005370d60e9fee2b71192e16b51821ced721d9280fea8987022e32f123652c74f051ce2cf408f30b31fd5680815988a1774bcdb553724db2cf164b59e7c1b5ed9710a044d74ee03ba1681b3c5f7db159f1e911b0c99d00ed11ae98c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he0d5ea56828dcc8d42a27ee7a062592fa0858b18e7a7661f69b025682a8863ff7a9b21388954c21dbd78a27a09cb347667f1c1c849f13d2f0291840015321d762fc713017cb0857136acb0705338245f515717b0962a3847d43f6cabff9c7a44579098490a7b89ca144c28158437cc6b5d36328075dfc2b7f0ca1dfcc3fe8892ec189f6fade84f4b9544e66f8ffab8acd0772f93980371ca2d35901180420484ebcbeb80e52b72132d83ad6bb4cc7b7193ae072a10fa60af1d4fe7931199a42556297eb77be024f7fafd816e1667f31f5fbd6582f414186c96b5c5338a949320c1a45b057900f66eaf6f7fe62888a3d4f48ef3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h91ce2e05020f955a3e66e945f315bd4e70bcedb3714e4a749fbe6c1c997d95ca370dfcd34418b9db62936b5f500e900e694e4a05b6d1c273124d39fd598d8d9ba5d47bb1450129101524c2b5117c99adb5f583db9f3eff7972e68e3085ba22b84896c72c627e775a9904a1dcabd4acc3e3e9ba09709489240fcf3e2e9055d37ce91a541b1b2be94fe126b99c78b592cfbbfba471694ad49781e31c15ec19b9a7f8c718622cc71bf2fac132b687cb27ec1a9d0bc74200a63b32a4451229e9e98bbf521794b76e1cc0c2d82ed0264b76c3b632e3442833fb7c48203f35f77e8beb66a6f9798bb60e3a01db4288be2ef06bf0772b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hbae2fd505ddd7d3fec4fe24d0208f5dd4d61c65c92ee20214e8e44d1ac0d3de73a334c1f57e87d8d9bc72d22f51e7c099c12c2fb4ba31ba37436a1e9e535f2b17050f05c0db4254b9eafbe93bc963da9b6ce5208296831b69fe5986209c6f47807e48e46f458c073bc72e2253e765e80ec29a9545fd78be568610731f257aec34548ee966463d3884fece22f7d433151a65e50d71d22ea0df78d54c1bacc50df51d4d69f2d406ae2dfb624189142768a4fd511023a8ab2e60bdf7d8dcee0af247747ac93c99208fc2f30ab3e0ce0f993aab5fa0ede5e9959c68a3135877fc06b2cf429616644e331d8f96a0375d6158df3eade;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc501ca20ed0255834f290abb0604407a7882953abfc7f846a61df6d4697c0f790fe0c61d12e2eaa5f581167aa55dd5d714d968de5c7ef8f8c841a6d5133743360f53336c0ede866eb87efa894d510456cb7b75eee2f3221621060cd0a051e84a3a4f0ea0754cd9d68e526834070cc26bb6bbb1ab263bdead609ff05ffd69f3174f61679fd702699285f6900f4f071280f27547887dcc8e802affbaca6324a5562135e951e5b1a2f267674ce687b94c139c4865d0e5b78f9d14503383abdc04487a099174a0a35bf557bfaf966d5673a5c27f26725898c351aadc5b22699aea58871935b0d8b0000616f8a2cc77dee8bade451a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9a77be33538d1879dd3d35c1c60a30ed00718d18ef3f871e8c35b6f4d4f4b971ecade5dca4f2b464fc6de829415f615d6479e8abb04824d37d9ad6c655cf5d30fc9578a82b9e62e59357dabab17ede3de66d0b703ba908456cc928fae9bb144a850cf0111758521799859e6094725b91550d784ef9063bc6fd8a554396556128c49ecb6b35782f732971ebfcdf85d2b4959bb5103e297f36c876a504449778bb44d4ca37f3be7fa05700266e883e64b307aec51e3dd2abddb515ac447a542785c7aae313042c4e715f8fe737520ef0796a078c1fdbff5f974559b044159acbafabb8b3e89d1588dc2813c11ccc8f365f1ea88e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9c154a63f68ab636c5fa0e8477e6f596deb97ce8360ddea5f7068bb78e28ed9fad6ac370048a1f4e511adb45c4cf6c86480501df17f8b8216f00333e33dfcd6030b45b624e98c9ab41ecb5ea8fbd94bb52002176ffa67d19f2c7789484008f678ea290e4662678904facf993ea740ee4386c843806eeb46646331acc5a5a87ee36fe1a28c2707e914ba58b4ebf7cd659d31c2cba5cc9056f457b5d0d9b20258024a2ef956b296df4571832aa37959ad709487fe7b926ff8d89486092d78fe090530b143a41a5baab51bd70b06ede1984028b6894eaa2c8c6b17e381b473f93c81c2c087ef0ef377fdc02c2132fc335d901c74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd86a599cce03a9f4d60a8931bcbf964be74ce469ba55e23087760a02498a5afc09c2a3a18ab3116a8221123981093b00617c949149e805a116e580d4bf4e6268fdbb00de4c0525fcbe323feea00ff82386773b251d1d02e15350cc723df11e017d9fd88a39a114ce7dcc30f31fa938aafe5fa2fd9bcbe4e5b0c02695d3bfc569c370833a6a2dcd3e16e81469e04c13a15d371189fe1df2af78682af88ac2c1882d61fe6a546bb4416c3c342b1cb1034310926e5b3865c06c42eb08f14b7e96a999fa37629cd711bf336648ce2fc2759fc5efff1daffd6087f908c34dd68156d28212d45e19ba4435c1cdf308312b01f5d8f67b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h9c090dffc460122c0ced8eebac46746a19d3b18affe0e3cf9ab03ebf4706ef69478bda62b5cef58b8e9cc61efab1f0b72d19fa71fce1bfb1045cabf7291de9be9a0868d5cd5b8e5cedb254874e52ef6a9f390a33efda1d2dcd9111e302f69455f751f57bbd9c4f380f8372e464aeed6844f9719282a41742ddd0f2e5d9918627f22e7e04836cd9eaacc4ab59374f1deda6655e974f53bc67e3e3d2e8644033f5a483295bf9e940022f0ef41f3e691bbdd16592ae075b4599fbd2da7d78ac2f2ea65ed1aa4b279a11c8423050ab0960845daa08c02bf6427724034c6339d93ca46c48fbd1dc5212e689a643674e427283684972;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc4e64f411777b2a063ab682b621c52b89b5f4d21ebbca8698f4528128f744dec31efa833c4f80592c6e28aa8d5f969b087ea8a3810b659f3385042362e3722df1f004ebf64e08ec45bf85f5fd4c7935fe0910a0f57ff12ef8b2f2e0a362a902e6623f81c438a58ee8132bcc2b2cc8b98e918ecff89f90fa216ebf2f2d2c63cc620af7b6d50b6a74ba17436c796172754d28601a8d71937f699d8a6bf8592ad10d3123c8a1003dde202197f25f887b13571ddb7b861633067c8202068ad96f2527e0b565704ab703171efbb962119da2a7d1ab153bbaf6283962ccf926d97c42d72faff606734c504948302db032ca060da6f46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h382dfefe6f2f1cdbd9bb8cc73bf452776c2666e5efe3b1494e7909f1cc8229b21b105d97bb61fbc927b8b4de81f85ba6d4b9c0e9b1e5740035ece9220ca9c3ec8c6eb06a11e12fc74e996964ac6a01cc496607555eb0729df0204ecdd240033549b00553d7d349e33f056a53c54b0b5b2fea00b5c09275435d6a2919f150f8ed92dd7e5c255889a02e0e53be3b8986a218fb2b2d2b9b40b3f2c6cdce2a579a52819e26373ccc685d4225daffa18fb62add48dc23b09736a229076cae148bd7aeab891d4b46dc889f6385922d02c0d27a8fb5a67444a689fcd4dddf8cd5e055446f58a3c5d2d785f30f9c0d5235233d424a4050;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha478753d3ebb3493c9361a6d1199dff3849346d0a71e0f22bb6a32835b1e41b751846059df2a441cb995ea786a6d3a57fcbdd5c6b125a41625f98f4306303c9b9e3c47fd150e68402beda22a0d668c2d0c683fd2d997b21020d45f5c5fabaf1c5aec7dcaab2cda80e8c493c7f712198ee360604fff5c90240d1457a9647262eb171fbab872a972c16412af1facf732157872d4711a6bed55afb33099a33a139c322336134a494082d214f32c560e100401c2175cd325feaf514f2c2bfb1514187c6ffece71ec97d6599c8d573015f345ef7bf03c821edf85803840ab978e43ae886394d29e6704fe3815993baf0073dc1b1e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hb63c24707a733ba97f09a07637797e05cbdc8fa9220e26b6757ac3b399e844ba89a58fc3fc0ec35fbbb093ff3937f9f53e4727a48fd9c35f166814d22506761d186efd34b7e8090531c824f232acfce3c118d76a8f0d44b21b2ae8b25b854f6b49ac1de3f32475bca78a05e5dd0bd6d554cf53c54f68f20e5e487d6926aaa10f068070856087b69074043c4647c0fe6930a9beb7a4ab9c2458422b84181746f27506dda4c83e83e0e40efebef1ca6817de995d9538c48bb0401cacc8e0dd9947585666eecf80866c82a67511123a0dcee6d1650c16cc59fbc37b701247ea38a2ef79daea734ac2a0eeee390368f21b4130d4c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he9d5cc48576706a2767463b5bb374a4c66c1ffba82636bc182f18f25afc6986afa097c5cc40238bcbe1701078828b180d099fc80817078b54f92fefef658eb6d707925b58efcab68ff276f8c0bbdef4462c03a6cb2d817febdbf6feed44061d6483a56a3fb197932b79ba500d47763d4ad4a41d01801dae32742be53b3185aa126885a6389bcf5081a56b1fb8bff8939678bb24dcf55994330a9e53a7f7d24dd88fc3f2d134e7491cebda7cca9312428cc9c6dcf7e8bbec6b975f19fa982e0a5aa63780b1c0d4f43d70008e247743f5d11ebe3c44be308c3fb184be370a0c5321b2c7fc996375af9e699dd88cbad418da3fa52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hfab48211d241d0d60c202f08ee56241b25c7e6069b0cd97a8d1d98ce82a3f3ec65a3c7a21e4cade88d5ede768f90ac70b4da19133526c1d37a6c938a157be6a4dc650a86c877dead59d31f350044071cb3c32f0d1671abb72335e592581d959aae7588475ff0022e3a45a04a1032dc8a6d219b3658693c6567657889b4162aee4090b8e231fb1bd1dd31e333b452322113aabb9087a5e4fad4b7216d1018ef6ad6d1cb735d4f77f9791d0b13a69dc98f3bd81cd4421294851b4e78c0886ba87a020576ac5d6f8a96ab4bfdcf2b7e5116a1bc6fc6851b821dcaabd477a4856baca29be49ffd2c901259afe87012b65da4aaec66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc369cbd6cced3b976e49e1ff217e2936ab3acd66c99c65929ddee109a4891ac360c3984c6a7ece5d8e96c68efb0f19e6f82b26120126bff78a84c81632e9c2774643256b2b8daec8aeff8250c5876d9f0079e6030f924a0e37f85a62593f77dfb6abf6ad11011ae46807df0df339cc6e0c2729b458a61d0f82774b6a056730343fbaf88ad1d3a9910775482dc4ac9cfe1bf0900cc5ba48b9df03794ec35f43031e8502e638b1713c1442bf3ec4a4c7430346bfb5c993e8acc40fe28f01ed10ca9a086de9d8e66fba269f1895ebce2835d7daf11646860934416c7058b846a541ec4e9c47b025be38212bfa597aaae5fbbbc4df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h50b692c063306397b38580116467dd2b708b856be5af1d8d9bc6cffa526c153b790b69028a198d49eaf3b652c25bd5b2b7fc4eb74a8216bb704f77f9abfe522fae154a390aa60568a35d2dbe4720af1742838354f19ca4799060f93f5d30672ab534935a2be029080df6b166539f714120985f337f5fe04039267379dc306f71126b46aa3b9707c1c725dcd2b233562c384122fe2531b2d58e62a821ee2c3f22bd2c7ce188b7a6834839915b5be6bab0a2f689c1b4e8e0e52386166e792b29fdd1c946205e68403bf3b6c0717e583b055f980fd0c3718845e6cbe7093d9ae5ffaf41a0b6e70c68d1206d51cb069426dcde390e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h140f5cdc8541088c1c4f877fe74810c659af71f2f0838b9a43395848f031dac7b45d2e6936f4fb61973824da1298a2d6591d196148c06efb566862227f039e2a7728fbda793c82130c7292958f60586e55a6f10da1600de4dabc5d99faed279db549f0efc6937765bed690f7ada392e85c6e3a7e89979f107194d5820b44b9a944cce9bbbb6ef7f6696ca56eabb974c2d2d1229d72e1770c6f43290e73d2dd825c616ee719689d3cd42b25cb90b9a9625b8e2cd903febebd756b4c3be6a030e2eca3a05b162aa90614e9ee6fe0e448d3b620be6d43dff1453583521ecc352537b4edc8fbe7a92254c7e67944dff556295e515c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4928a492f035877563e0c4b7039acad1264b76d050c73fdbabad1914cf4fd16083594f1bdf55fd59d107dfe23cba83e6606815969e5d55d3d9537f63983a5dcd062dda636be32ebab0dd6e8bf9bdb54a731e5c50471bf8845a476242cec39c9fa6dc6ee925d330a7712ca1bbb0ad638e018509f047d2e3027c37118558a6c9936898e0608d6ced6b71f06ebc8337b6c637b97944a57c77e0337c0adfa77ee382668f78ce45b794d763ad4a2a3d421cbf1eccd24a37bac007aca619b4fc1255e0c1e8a96ab399c97eff33455d7b3f81bfa83f5bc3f03b0eb3ebc017b94c09bdf13ceddf22e60a6d90fb7f68f28813156ec61941;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hb171a4d95c2ca22bd90ad37b790db1fabf33e10cafc5199b439a1802bf5b53b3a0a5887ce284942046a3f04385e665d261ea96ee194ef61d675d7b023e84145d2d39abc3bfc86180eab0a7f67251c58833c93e12f46ec7ffeeda7b59f01600baad02d114bba278d95706ce4d5318dff7617ed838d9b479e614064a45be5fedcb4eb1c595ec816061bec45af67ab3f9e5c81db8f2253884f0263a1df169813f2e79e91374fc63b416807c4c0906eca4d98f17fadc31016e44a2a7a8ecbb3afb88ae3698cb520e04c99b3970037d1abd17d65e1145aaa039dba000c740a4ee42241401e7eb62249ed3f31406dff489f9763483fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h468a813381fbdea1d72c1b7320da2ed792b3e57008db0fe3437a216739f07646d183545cf9db0f343b25d8ae89bf044e444e95dc752779e4237de3f788b533a0fd46453f0077f23fbe389cb7b1c0f8a9c2591e8faf2f2b023ba60b685d800a1e9b21ff5e8e8c42f15e660075017d741af986fa2c6e4fee20b3da18b7f7337ead8ab7c8f103fb4c4f31f970b3dcb58b7809c2182af714c8eaa25cd78b67396d910aa7421b15f44e5329a5efded14344e38f0ba8ea6540d4a147cd38f12ab13996f117c4f4f8d38623b559b3792a3b18310b7f9c0c200dc1321db37b6357f07e59e8bec13ca254f19a50b7bcab971b9a9e7117f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha9303d58d0cc036fcc2271c48d94efb4cd0e535d4a244bc7188b5927e29e6e836348903bbd47fb0196a6cc33caa9c2d2ba52eef494e7d89bcc950985fe206f381348eb46c1fd54378401ec8e29036d91ac941220f86c7867139a6c367b5aeed53ef9893181e8d723e9a6ba42e0a0ecbdf1b1192b6840c36054110d799b591f414647e74326deca589bc150d8a86dc2027d2e67cf48bd2725734ca7e2e1cac21e06d855c4fff54cf8176924fc82dc8b7edad40e052d69c982a09d78ad0fe1441c275edccfbd29f451858ae7b41609807561a405c07e56b7558728869c8a184f887e6393037c74f16bb26df55c16f17afd46fcf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h425d91b632fa9d0e2e0afecec86c988d8774fa8ab7db9e09519915a87f78a4c7f237a78640c01eff1aa6ab07d5ae88fa2565a30f775b94196f98084c7843aa230bfcf374f744f6d14f7ddeb3cd294f41e7e7a7a40e180d606e64a4742c189a1697c190b8a0a6f45c59dfbace929df629a51fec5c75527dbb309c6672313121c1cf815de054d6fc14d2bb1a9133c96ce0e0f5f8393c8d477ca8f87681ee170a2cbe4a74623c248e85f9d52fbeb2782046a43cd2d057401b0194ff89f32e29d0196c3a66e252533b76c09588aa733ee6f0d00b7bbd9e8193cac849c20fb5b3a914aa9d9bff41377af3a16d59342202dc286d6e3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hbb63b7a6d4708dde7aff96d5edd033db80d0cee90082503a53d78bfdd2e95a9174a0702c9d660f4ac07e26df23f20a60919fe96844b5828a2214e08a632ccfb8da93d91fd85c78d60fe55360f3c00b184a2ff52df71fbc52ee4632fcc58695abe30e4c7c641f4873508fe10da8bf48e4d1a9ccd1462a8d73f8ffcc890c689ca220fb8de555636d3a0f82e284f46e29ed45c1ccbe72cd007ffabb4129b1f7680a92fe150c81208b0990cd4d1429f157e4e889cb45a0a810e9a4210bb4d2186c774549a6e726fd7f3835e9fa389f6f59e3acf96405152cb8074b81b5e9218de254d43db71c178fa910c53132711d42cf23817038;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h71ab549bf66d1f4e6525f6d38af7591789375bed965d372fc3c32353e96aae03983f15ce039fef013826093562401404537a53105097ef3b8084ecf79db6fdcf54df1b5e9d9bc31b0a554f0d348d1e6094baac0b3852dbeb76d73982c4879b1179884a40aebf72640644dd2d447d2db6b036979385b5b5fdd5a9f37d5ef5aa8697bb338c9cb4201fb498a04a34eebe847b50e426d3ce90ee553c5626f62793c45a93e68b5c141990b2428b41c6c28238d054c8d6132ff9913fa12541540fba2372128d0095653f95e831bc77411e0bd11acd5b5cff3a2d29f88093a26814f982c12cc45d5ff4f7076383987612e437d118af99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hadc5271679625b2d00f8abf98bde5e138f85244cf1c17eee4d58afbcf896be83316b93564b41f19e19ebff7b4234b182ef683e96ead83c07082c6e6b964a0b1b20de58b748e6241b4ec84d47a49d7403dd5daa8475920c71b265d355f7ae00cc30aeb7855d3410bce22c8fa0b323cb597a36eaf0f1e5529a810bb2f376f94e05fefd8bcad2cc1f97502b8022f9aff6bc1961401cf3f9543bd833af10788edefc63d10e94e43a4801320c981c113e912b905fdfb4cdba25ff66dc3045b5e0b48fbae089b24bafac6febbe1104135dbeef7b2a8944df0c50c39884c2c2bc5e7ef4272d9dfb1c27198d07b9ae0110427637c8bb4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hf5cba7045b256566b3cb72da54dcf1c946ad8ac9eb3f9693f354f7b403d097410d945642efbfb56bd69add6547d391ed7565349ca40f98ca199fe792d3d56855e268749887a271611c2e417a09fa519e2092693dde791be4b8b88eba73630b33284352cb76ca6fedc107f13efbc995fa80c5145148d5682b9e231a0a6ba6794f71437bb4e3c2f91b1d9abec911f7bf487ad6ccf735c41f7bee96c786620538d277883230b617fde5cd80429f9515428effba09b7c5062f0e95d50db1fde13aca39d08ca551c7c271f28f5ad790764579c117bc992bbbdfe4e301cd2f7758640312be418c2c12927f87f0274d8572e08850c86a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3e8a50e644a74aba044d988bffae2fd654fcc47f1ecd7286c77fc008cc81c3443d0b0e9beb3043c889ea87fdc2e91fdd5e45726e963812f577f4fdde751ccd607ce29ccb3a973ae482e462504d01f8e0492f69efa30b8ff1b114b7f7976656a70fd9916c4c618e6e6cdf678fab6b52dc76b72adabd9e146100ca4692744fcb140fc8a2d34316164c8c61db60d06ab49b3b36eaf6af0822d7be2a477790ac613f8bedb0ef3d19b966a4f0e2927571a310097b58d96a0d1c3377a4bca50969a9cae2693c7fbd40e4563afaed99d8b147a2118a8735ce83ebcb3dea977b97ccf6e73f44a9d76884a3dffec296048288d45d88707a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4ebc845ef703cc3b782729a09ce66b082260663f1f3a0068523a7a492c763e411bcd31f664dcfffe96088dc20e3bd481b16e9c6fc3617f0d7a7e72c4e5ccdf1fb31d81b52f552780a599872fe539bfbb839ac0e2d61e708874ccfc865c6dcd4720d2e7a89141daaca3053d3459a4b48643db3107c25455d31d1fc3bb14351b08c54b02ea2712fd463a635ab39732c4ab8c79678e13d7ba0e58c2a3e8eaaa5f921b731d2ec7877ae7364854195482a0aa65dcd4a45b6774c649a6b0b1441f82cd31bb5303b6dcbc19813943e16f5d9d624eab1d0db67f150857fc59d60352436ff6df03fb816717f9b0f027bb58de8da96f2192;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h81660a115faff2d5fbb58d02b568fd532ec20ca6d267f68adf654f64698abb5c1d183519b07571e98eb5debda26d4700624538bf31c787b7a786d99366c45c97e23b86fa132bff8bd1557f054caf747d876211159af5467eb14373ac5333de61e3b670c58243706446910abdf8477d5a230ed0ce65fa401a951bf647dbbbb3a0f24b6c696983e3c63f4cec966e2c4f6324fe83da790dba34479e7e0e6176de0eb8ae1d359f9e1a8a8b33fa7e2fdba918fd2c8ee19a78ee40783825527b476bc130a85e0af65f0eca2e55ab53b13c39ee504b4db500305feeae11ac85339a32c73235192b50a21cc2a1cd5dccc934955bd4b662;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h850c57e46dd9897aa50465712e501ecad66c827a71d84e24d9d0bcde7f50e940a754d8f165bdb8669904e1abb90ee1ea147beb464bd665632d1d55e917dac41828f497e50962cb60a997946cc1d1a29aaaba7de9d475439191391be997e9862612b0218bb79bb14f4bb940aad8351ca66bdbb00a9a1c87cb38c63a1cda043d0cb5c7b9b5ee898889acbe3a431547ab74bbdb9d26af3d7cb9d3f3b060791953ad1d544bf698a6fdb9614c9ebb0b99e9be39a214b746265d8755b68e6e593f24a46045b611f075d10c7d59c150cdae5953621253dad95176c5af51001a11d004cd4256f64fdf229b06c02b6b2b52f1936f1985df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he67c33d0641bd23a84ddf4f0be412dfadc6089d8ddbcf1adc4bb95945a15fc0dba80971747f69a22fa29008345dcc11a869d4341f8e5bc2b61b57516e1328fbb7b8c6ca8a392af93e9f100d7abdc7d2dcfd268e9b1814fa70b08e24d26ef9ff2b8f7d0b0deaddc2cef3a4da71adb60e91f4adaea126f34e3df9fd8c18a0b65a1e19eeb31360f04490fb2741a0a53f1fe9c7b7c8fd8ea1c85f1566c3e7e3ac2c2ffca344740e392653454341859f568569cad48a08cbec8aa7ce4127d840e36a8ca1202162afa21d040251916b77f783fec6fa7a22070451226eaf09836f404be446962a2164cb7d087498ab61e12200e71ff96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h612fbbc1e0626d1a61506b423549be49f78460a2dcb27274ac4089ddbd7a781efd758e0ef8319a620d4cb85a6a2cb3245354bce2e456ab03bba269149493b927969a28a24255433e32c40245f9ea54afe5e34acfd33506cc92642601c3c69aa39e61c2c07058fa18716c83e2bf52bbc979fccac65270d1aac1f0adf762a88cce189f2066743edaa1ef85b5a79cc7e74fd87294a7785bdfed42eca819567e0209b5aca265d49a1813326e5cdb9d8c8667785521d77c2f73f1b3cc4f8d4d498cd5c28646840350629a93c59330b772531522dc61ca69e471d1cfa7c0a5086c7a5144a33e0b4ac387a240ffc06db931cfc407da17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he1c9c37fa1347bd75ff0d5582f4e13b88005165e91b241da2caf13080b9a9a180b6b99f09187c53cd2247498050c19fe1be19e5bb39eb53612bebaa336d5e719f14e49203a4772985e672ef06fee86095f0497eb98342201c88273e0b488018ed85608517debaabe542e8a2ebce9ee7aa3daf00a8e53812250d07eecbd4d8c3998110000e0f810a3a3d0a5e10194249fbbc29126ff8f8c191a49dc02724f97877923915365c8f5b1b83c658c4af5ef54bbbb280d36e7d7f26b38c4fd2b375a8cd91e8836d1928dec771f6bfe5a84e638869ceecea1910151d5669396a9c596467dbd92dbdb1bafab5881d64a6122a9da2d91f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'habf6d0c49ac1f97e09086a4443675c711aad3e9e615b08d76c60420cd782c8e435a9708a6f93ef80ba20ae286413e44dacaa11cb0ccf9247febc9c2151bde86b251b9f18de8282c7eae00f43c310d523e3644039c3d70573cce9ba8eb4d581434487a964a200a5d669b76afd0475355ccdfddc465bd42e64a4232eaea3c8224ba5be5caf22e202ac6438413aec73f24082a482a177ffe3c531a0ec59ddf9772475f2e7a3abbc8b6c8c1bc19852104a1db81a7de5e7217b0ed2ca5ef53f83d5f1a569368f2ae74bb4398c41d5c12dcbea116f9eb1940be0555e158a6efd81b16c11b924c1ce48fde442dd5877a8d711496ed4b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3de245f86d28163bba9dd661246e5126c311903e56e65ddd6589ad7b27a14ad9a3d65c090dbf774eecfaf46aeb4aa807c1ab97c9c0d0b37bc77b4f0510982e4a0351373b21eba846d70b7bacc988b82e7312a29326613bd0374aecf34eeece7f9d2e344b6a2f1fa14516527267871608afdb0008bb05301087e4685e09890955cb10dd4d19d496457baf93632d8097a65c07c86becbd4190c42e38c2818377dc465f910a533c567e64c30e6b998ba37a979c9d4b230eca9e8807714bc44828b01fc3e374952c52f8b2fd1109f90c5f768a6fae1d4719300f0b3b7a1c6e55daf3b378d523e311db5556dbd234803053b839e00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h853bc3ddae3de14fe43f40aff56ce1402a16aa9c870c0daa5d544fbf2e06f6142567d9f575262a3e0d7d56ed5b79d6004966069cd4ad0457eb3d68bef18b0864d4b5ebcda45cced77caa54822c3b9ec83f8817dfb212e113b564b947e89f5101b65731e5767ee878f660fbd688be8008de2ba27c876c3852d0a04e760d0dc2b7d815351298004eaaee597a641ac5732de98db6f7052016eb414dc877fc75064f6c234de1cfca1e2abf92c97fd55f027e2cd074b402996b46eef3f7b01b8fde6925e763a95bfafb839a446612264206d8bbce6d53673c0834f4c213b4106095dde6c97797a1bc7113c0fd0c2470177de2672499;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h67f6b43a903a18e89ee87bd9f0bb926de216110aaa0e2586f13524ce280d9ef9612e87f447bf542254e6e716e35813f333c11be0c17bb07a2593f11b4d9987f12f7364138ba923a4d3aac6390a7fd787e11089eef8b45a4425c21bb2e21e693de1b52b2e30f7405a9fed05c9bafba70546238f575125d7e2804dc6f3bf86306a52ad39fd011a94e73e1e5420c0089680aa67125bc2a932d5dc35883d45d3b632751c5d695c1f68637f5649cd4a9e3bab3ff0f563028a6bf204110e83885260d9bd449ce1fb1fea7120392989db2c78e0ba5684ecec78ad64977f7f347ea0fcd61e2417d920224e0440dff4b3d79a06dec4971a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha7841e05c0c1e104f942d75f0d7cd5f2e67668ceb282947a195e328a14673ca919e1f7a92c3da06eb52c5544f1b880242a7acd2a4b13bbc0f8fc77cd7e283a0a832ee6da0d922beb912202289974f4da9f310490a8afa32ebc1bc7b09c5fbbfc09c6c51a9acfd5b3fa7887a04e8c88698483b2c936d699d7cf642a864f5a761c35ffa4fefee4f91f6dd2ec72b79e9e0fb2d649d8dfa854d60f7bd1dcb4f3211d0f5e216e835b00e00e99b549272a738608ef7c7d1a96aab78923ffc5cb3ff7e725495f102b8c5932addd0d99b65abbc2ef45c7a8f764f8391514214caf798a69b702173792d67e70acf91e381143ccfa4019be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd309be99986935795b4bc4eac44c421c58606fc8ac027530e2c1ea25e600e31162b8a80aa9209fab9f97df55019a24678b7f23768979430bca167ddb45c40736ce9f6f625bebf1b2cb31eaae6ed1d7a25477415e8652298de05e4e156c9b4b58c03fe319ed8b8a662ca391ca38bfca6540eda450aa7dc7a83c90ee1dc25f8026c43f0e05e5ced878ffc0e08ef078491b64a9729d461536df5b727fcd4c4c4901e370c4d086764f90ff2e82488f24d1d6164d48a40e09b51cc543ad6461b89767f289c27dbbb2f53277300b4e8cd357331bb7952d561d288bc7be5d29211bc91582897e907ab1daf6d23d6806949070278de90a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h26e1bdaf9ab0a0e251ea503186543e2ea96df211e4e23bcaf5958957db02b862e475fc9e8eb04233276c43d13adc2a3e47e7a6c2006b7683e07f8951c16183a0a2b9b2a19d321405d3fa4365b1be31ab3d51e41498ab70e10738ef0b7c8a35eb9f5a272314b50c5b767d74a15a928e6baf6fd43395c51cc3ad2f50ece05432528f17be508419f023cb0ec318b34b58c0503403ebb9eb6632b20e19df23520c77f61b6cd019af1652267caae2b1f88bf8fc161d0c54b2f404442223e91eab8404e00fde924071fcac3b095bb5c121def93be6878560e8955418b3143f383021714c549d4161703dc9bd350bd1aafdb286f2b43f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h15e9f2a8afd4fb43c9079f88f845b92153021b3d1aac4010b108396ef20ddfa3aa0d78c2aea348530fcdc45bdccc5460c56943ea317e76abadbeba6d7d303f3df9afefde4c0eeea312da09ae829f28574f94ee2117319a774dafc1c8d585b2564481851c254639f90627b1b03953a4541dfb3a8b4b9c0644dd891106469d83c3fdcf9abbd02a4ab4682dcdf0512483a9ac6c1bfc1000e03647c9c1305a12ab59acbb2344d37fbe88c0fecc54989579da6f414d4b67ea723a4de3c85bde4223f41cbbeee3b6ae71cb69a9a8b5d2464c41470609dd377f37ce536d889ae09144ea0c3396265b89ced720ea0bcf7d0ba178debe75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h85bb6e93d656af739cd5d5376bbd8fcda89786370b548d9d7035743efbdb17b0e4a279247b280e4e8b9dd917b94648d56280527357bd03f0ab048e696b72d0c7939e1a59eb89b61026d02352dcc51ee57e87e4bf4360327132a6e2d069d2e3117d3d506a0dfd0fc79470ce7bba1649ad03965225af2da5a28a4145206691e6ba28ffc3f4e24bd7931ec2bb6e72b8039a205bb91fab4db714a65975bc6c799411c4f614aef02d671019d5e0f9166f1c216bc9dd890ef899904c1e4ab23c6b1d6f4c7f92e5256bd7151eb26872cbdbbdba73f5019cf8b644469a5fde00a4703c15354792abd34913474bca102c6a037b4a195e97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h67d0a81901dbb1515b71497cb14e8d86aa69372d008a8de58ee7cd2ac87a5e61526a8ed4375e4612e9889c331814b1bfbcc2eb910bee30c29a525d6974ae66f9095796be5e186cfc06886a540c1fe7c7832e256e0845c10b4c2b26fb8033dd2189fc38d0668584ad8b717f11d71f5065236259daba0bbabc7bfc78e68cf9689e0ea79b9bd40e45380dd5810aad4657aa58bc7b0a2dd2b26d9fdcb60b4111171c5fd790ab9221f448b53d21f125eba49b1615805ddf9f0b1be83f9e75549c86e528f81b504374187539475c7e58dca849bf80d892d54d18de1d25c931903ea475693704bf3a8e9e1101302e64e1a449cff20a86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'ha4f3220e63412284e7dcc509dcac2315169d437c479357afd1d02b952da9d5648f277cd97913bb7d314b855fbdbd85e30d65b9dee11c74fe30d74f1a52770169df236f43cd1f5a0d5f26ebc886a00544de21bf98cbb9717ddc09da5b334bc6e9f7e2399f1715aa225b6947dbb6c4dd40da7589750efba86877384c186c322f3be4e280a79787396df8cbe0139d6f5d82d9a64f543d7720048362585ec5ca023edeb7e0e453ab0ba1971370c3dba7d68cc77b184b2cf40fe0f8cb8a5ea54114602351da0e008592e10a5686567982b1c5e3e0d43cd6f7c2a4eb9927e3f40addc5818c86f86fb115db9d75c386c3f5c8f81137f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h96a5ff33d89b4f9a24389aab1035066b3bbfe4b1be86bf7ff25f8407c828849dda11e440ddc6137488dfdffcfd3b3afe6352617073b0413a193a020edb79071ac6fedb2e112beede0a0654c60c7709e89d39d00c4e107d122b0d9edd335064bab5513b9341c2fe577770c7c2c9f7a58e1533a743f0fac3b4abb09015ffbb7eb6ca3f84f9de444470000ef1da840e0897106d3e1003606d22d75f3107d2114bde5ae4445e72ce81a35b2e6c24690a03eb2a68f6852a7b7708d3e9fb12f027d2955de1196fd3233f77f2153867fef26f6eeaa5c86ae3b310522605b835dbb58c663f2ff5ab1359ba1bb47b8b8b8f7e1be1fa204e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2f4ae59b503d7bd970fad2c93614a60f8c41c65e399d49c3676b88946d333f803da8a925eb0e4cacd1f2699cc1ec4a3a8c205c2460f6a198076549801896b3b55235c1a46c0c6fd9ff9b7208f6d87a405b18e942765f8eebf83dca4cc98d5a4be2a177e3ecf5ae3f0ab2011f905442f9e09653705a2fca90663d4ff4d0ce127e2e224dcdeafd97de9e50c22ef5f1edfc628db6b7ca05081c3d77100c2ce614471c4300378c494ae15588324797462617c7e31dd2e2f084282a6179069191efc7be5513b9e1e3d70d38c7fed4515d483b495c443e17fd3e350a5ea70fad6e2dcd111199fa809e86977880e0d920c23ebedcbdd4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h78774833b6542629c02cde5d0005c02facc082815434bd081b78879961371ad99c9b821ccee346d9bec039aff372f63fbdbe99c157010a424cbcb70884b9c193005e0afb457f747792232d83bcb7f82cb05ff69e6a0e481832905a1e4e586f3c9d2f2a0a6e6306a83852d73a70e38fb1ccf962971a742abafc43d32d801724739c5f007e7b913f377ceb03c6febb34ff60da51d274829d95d65ef0e30061c867a9e9ff17516a35e44d8a2f3603fa60009c11f26ad951d0d93f6a973afeea9d9ab8f48d106c9ad713cfb3d0e2d4e426ca37c536d83e1a30d3094bb9f3afb689857e5a4fe28aee35a2c6f1e9504a105767360238;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h539227655f684b4e6f35e4ba970c8a35fb7d87f9cb6e9f05bca6a6baec68f5b5118f5070b6bd45a79a779d314b2eeb5d39cdac692619cfadc28143faa6b80f59573146e27c78f4dda63f5afda5912e9549a4d93dd85792c508348f6413dde39a16cce90e871e9f05f326874c5a9432dfa1df0e43f5cbb0c34fbbb9e0ea1e92223b8d8eab0044fc718f0ca0ef59455e13572df69c0c86b22ebced70fb6c621312e13446ce4941d8317218cd374a0dc92ba0f9bdba87a17643f777a93d6fb8e23e318e8100965650296c7f7bc26a247f04d7781cbdf13d0745e87fddb58d0b315f3aaabbcf0290f950820a70173dac96fda1ee49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h13bf373734948d0f5f3bc253857a90de330ba8ad50305ebe5d37646e0dda8c55a1b414a428ba932f6d6e73bd78ec7b59849229bf6df5dc346f0e7d5abe3a9c5ddc4b16880b9ffc73e6d557ba76edea65a8ca399d30a8da075d99593a6e2bbae163e9a2dd31a46304bdf63ba035dfbc0d36abfb3476ceeaa9e86cbd699b9c430cfe2f5368eaf3ffc129db0ebe218d371ee4a1041ed05e1b1decd28cf0b3e6ad63c61770e60ccf3d9f311c7987701f8e6b871d978f78307582925d0007075f9b35d2408e168d3611d5cdf78a3bc59e903c6c6c143df6b61252658fb9ae0842a325752766d69877c7ee727805c931404f7c9e195a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5ed71ff63e1d4f3bd88f30628cb181003af3bd99d7bfd37f13555055983146701193c0293a7afcedd72a5105f9beef12d11f7bb12ddad3d20c746b9bf5bfc234b1febc7d621a8efd7cd5dd1d238ffc106332980e815126841ac845380433b8f2e2f9a5ed0d0d4de8abc27050b183c58283116e721bffd9ddecceb689a8aaea83271db8cff1acf7f1e9abad2ab1c9ecb477842a747684de0ae437692a329e54aa9fdcd6432cda7337af24d599a0cb3778002a78682dc9fd1cfa5947acdba74b8218d8a59a2f78ed864dfd5ef59bb56dca98b3e7b2e21c6057a87b275039c53175f232cc51a1aaef4b674ba47ca99b15099648ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd032301787b81c0629eeebe442d1d812587400fd48d91659bc1c2e7ab84a9e4ce91705e4e71d2202a195f1e10433350dbc03016a5987558a66fdaffaeb3a149a96e198635423199be695b07e68f65d593bbcafb8170719e7a7e3be7dbb1f604b1a8df6736377669eb364e33e8c776288793dbc8bd50960984519dad46f126348a43e44296ef21d48ad32ab89a6cd298f756c0f697529256cde5020a5c6f246db1a7a7a51737437bd9589fef7664d70426103164a200844b81f7f8c4c9355fb6fb323355a23b7392789b69095e88c1408de3842b8245f177d6feedb462d27b3012b7024d5c4240b57ac5971cb12118d313f1569;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h54b97ea3249c3bc161383044da7df97204ef78d85d86ff8658cc4b292ef72248b34734fbf3659cfb5f22e9a01077ec728bff7a4a527e878dbacce139e2657f7924a7c15f9fcaac9ab0e336703cf2aadce2e02ce46b55124e93632a08f3387fb21cf5131eddc0f5a9d698c18728084d1e079204f702c7fc3d1e02fecf66b9474dae3003d3628e314fc53b8b2699391333882b412e6ca60ae2becb078fd3467c6ddbd35282de951848b0e34119067a352790c79e88c5d9a94cfe97db19fa8e4272714a2a4158fff286bd956d9f13cf72f6cc64e63c36c752b88c5e953e4f73786a2bb19b375fccfdb2759a1b1ac08ccc122f0368;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h31179e2395e1c699f5b282934a9a819249b9e6ce846b8f3aa0eb7ce730fd2da368044cb728e097b94a7fb40637b0a345e39e1a7a2333d73186af2974fc393a0c8a15a9cedcdf14df139bde2361a31700a75b06aad5cedf69f05d2a8d8d67a4c909d90f303828e5fbe67be64edec0c0692354443fefb1c30580b9399cfd693608c7aa1a2b2858bd987aeeab7dac2ca0c801b7a14fbeb965bf9210e5ce43f1cdb73f1dfdc7d5a496d05550d18057a20cb9217a71d72f15c6096af09a8fb13d535e2e097eee013f2a1c8c519a25a84474f870a02916be2e029dab17b6456ebda23563026541e15470de784408d003dace92b081f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h7bad4e4909e5f6621138d751fa1d9e16956e07a2ed099cc1edbc540b17ab4e42875d30965a675fc92c0414fc45f410f1ae43b7cab3825348e5f6bea63a2f74c85abbf8040f57dbed7633cd93538c99736187ff84a37648c23b5e2e932bb2bf76f2b1cc160d832596bf88155483373269f268aee2e94555e20a582259e80c03abf5a02160aec290544065cfb728b90b8442b5d29dcf18ffb0d34839f9201894275811eaa0f6a20013bf7f3330dbfd1c118f57202b7ffc45c6864606582b70cc1883533468bc71da35e51af84ae83ce41f62adf8df63392ba2166d45cfa0b4392fc53dcc9b8b2ec7d2837f28af2cb8057cb1e5f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h44ffae9e5d4a0daa3e044297f6509616c85c63d7723dfa8b2cd978313638968f8d94dea384f4d300a4096e08a77cb4455f0dd0739e312f5c12087c53d594ac96d94e94738acd56aae48ed2f8189de55df1a3ee8695fd02050cf72810eb81062c2e8f6acf084d1554889750b6dec9f711f44e43519080d636b083f8659e16bc48c68a50e7fc23b68b051707c432dd792fd5ec256f0f6d6ba3348f7ca182536b3b7ad71918d9cdf4e847677b8476a5cb389689e9125a2d3e0791f348e8a4e2d6c7e92144080267d082696275061191f3b9a86a83b4ac60d93b298e2e3c7fbe22f5161a7bdf55c5cb338bc0502981667d270a9b9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h5109d9215c4856ccf23ccaae239c263b5ad1c30a748c9bd607fdcecf9ac9c8adca9ba44c99aa13deac65c3625f344c55d107a3cea7b651bc402ee245256587b8f5d5544292d14d92657c2f0b27cdab6a41099a78c6ff127f0b0efa262eed795c11f3d2a2862f835918eb4eb34e76c88e8b4ecb244a48173d5680cabe0161565bdf88920f298cc6782bdc368733750b6c3fdc7d5860e22afcad8dbeb2b898c5c087544dfdde1fe6df1d05d48b381a9b3e0b6adc12f1386480f8126e860ef2d3c77dc504029ef9d84b2b0b86e8672eef3b4fdede517d97294397b322054ed9416b4cd6c40dab3238619334136193aa0942e20283;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h438b1cea9a07daa5972877d5a3edbdf841b45a196ef8e03ad093df9df7f7dcd2c2db41b54f0d474a2802eed7e9690ee638ff2c569563b8ab1912ca7f0edee1c4b3f00bae28d39ee82fa6452c0633180e7eb62b16bab2b10bf734e243f88d65f150a35d358dd4977bf6762a9a1230f0fac36b5f18a983ecf4719c93b57dbaeff10d0a5bcc559ae8b9be1ee2660233b2dbb746548bcc61ac0b78ba33fd8b5bbf0ecd006350c1d5698b89b04d4c78bb52fd717510426d0f24d9ea58cc7d534c5ab1e087b345e065ca1f063562ed18e67adf6e2e718be8dfd26c656b8f5a186f095eff35c2a40faa6c31cc911a23e52f209177174c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3c4592487cb2a489c4deee3d762930e4cce8d44ff6a5985a4146c241065fd6f1dab03699a42a3632179f0f7cefba88d264222bf2551c7f8451291609fc7b5e9d0af5bd364fc7cb4db77918a98ed2a8823da719fcb4f4a8bdfe957c8f33f52bada3c72ce1eacde2835ef4c64b1367bf7e705d200ebf3ef9a2d09da9cf53e073c401143fe818fb550e3832bc20383efefe1ad4274d1ccccffdee74a50eb827e4f88d2b9b330e9ee2469cf0d703d9e19154c0bc2ad63887f5d641009d6427cbfae7535c751138868afcd964d3d5bb399d25dda6b855040d42b410e4228b059e8a5921a2e18f16ce17b1c19a6f91d3689975afbfa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h6c1709bcd6b79918fb73d2d45f4dc377c229a0a293f42002888c7e9693ae64cba0b5698e70f197667b2e7f37403c58e1aad224e7091e1401467398c8a7323345db592a2acad3661110929f3f734b0d0158ce0e5e63decd9e04e65ee618b3b70e508a21928bb009a9c02f26e8d78082e93129a7a68c0e05f8a06ccd59ed164aa59c4d893fc7692f90436ab58240baa2e04d82e21de21ba7d0eaf1a575a2dcd025b7d8dd60967e7419d4dfcbb3355376a862c85c2b2e5c7b29dbdaeec062ec7cdd31aec74cd6310e54330730a5035a07906a6a420668e7a81e4b3c4ab19169171fdc402a45a6b3019f07c08375e7934ee1955681;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h3c0b39e021c6cea0d28508ba0ff0c827bde88373c1fa9074b69c0430c30ce38a89329743c863a603eab865cdafd82c1a182f1f23b606e92ad01c6f8cc41ab9f2f7ebeca3a097902024b78ec8d0d8fcb0645753f9fc1c015a2ff9a3372d1fdffbdac31b4d47be757b074ce2c173382bf6235fb76fe5463fec79108640de1cccdc4756b7eda4bb559aaa65f31cc25bafd1ab80a013ce4a757fe7cfa0d6cf619f9a76d6cc8500dcffe2febc7d1a3125973e918918bc0ba2b0ce1376954c9c916153212f04673b78cb270948e01cd7d0436902707c34f69da649c986abf945246f9a01ca9d6b00009cececb0669673080d07a6c20a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h276dc62b2820c508ee5cafd70e2faf93f7bda3f5e64647f17201fd9d87053951e449a354746a88ced6c3ea70a3e621d2d0cac35dec80315fe3940fe8de54a7dd2bac30d70e2f7470ac73c1f4af52aad1434eb3627343f013258516d758db3e5b8561033f8f06892aaa687a2784ea09c654ff2e0bd69f0941966faa194407815c99a459e849831a5e87df0e922567078c5c7553bece219b4874aa26cec3f9fe0da861132be5f405738565f7554ebb3a1c9660d32f9519221569c7f9d9bead33cf9790fa1a613e8a91b85727802e886d0910631ea906c3f34e8085068028425d86a76eecb076b3fa28bbd43f34c0f4f2396aee25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h280c776a477414532973082a08c2791aebe470048fcc503719f2ed2a0d24ffe063608705a1c6907c3bc3c34c4b0f3fbc38d3e41f53a5e826957ae4c0b03a9bead9969d01880476ffc604f10aa5aa871b62a3d592203bfe23555043153ddb15c654ec4bda9b93fcc1b9e133aa358fd34e85f2250f07f8fb0b3669a6d848ebc2f7e1114452c071395bd2c5582f83d930ebaf801c2164932c1232acd309d525082f61c8f8204b3ba02d1d95644e90c1b2957ce761977cd9a09af11c0f30d20531bccbb39b29c56dc3133265e24c1db6b79a84a0e6b0793ba57ec7d96a532f8cd86a870d2da700dd8ac38e75a593e5b201bae0aea3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h4f73744e672cf66adc3f5ddcbbd0f63b0ae9ea309ecadef16b46c9ebcca64e1896331de8117d1db1e3952428b690477a8d80e5f889e11045891d0720ad242e1bb9eecf93aaea1f0e7fe99e23b53e352dc5a5655e05ea940ca875a48f59b4f8f879735ee230ab76317b6a7efb3854b8cce10a2c9462a32178970d16c0ec3af7e7edfe18945a065e34bc5a30b4ab8461b54a8de6d10c6a8350b29b30eb9813b0b8c41641437ae6edd38766f15ebaa105d7c35b4a67e2dac4ead5278c0ff6ad8bb6347d84f9ae5b7954e4f441e1cebf6fe7b46a542daa6040e507b51d65bd0121ac50da4db438be76e167e455ffaa7ed44546b0e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h82ced794b333092e986baaf41efb97b181449263a7be4e7fabf88d103950fb5228e16462b4823ff0b728483d54a151fd6f3d785a9a6409db8548e55fab28a045da3dedc027bb452ff657f1534d959f677d7864e7d1fc6d582f403caa6cd769ba6ee3ee3b7089ecf198f07ef2e8d91993c3688c0f5c40de50c844bc117e551868aabe19ad3fc5ca380db564c5e663b1bf151be9636fda5c238a7aac95d150bc5d5f428c5e99c0d8cef9c175a39dc89672a5e577b4b424807769bb11e7e9ee33821b57101a20c19f8e7db68c354018b2cf4c00276c20f8028478da3599ac1f17e3e0a767988d6d30e10ab62cb3aad37b9d65bea6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hc23ef4072cd81bba646a886d1398b1e132325f2c1f2caf6c4de25233187ea6c6bef47478dd3d7eefd5ce8066e9f2aae98227a2082e17e828c0c23182816a2c93e8d127a4b2cff133770d2634f32abce6f2c3200eaae2e4b7100181ace1a85e179141758321525f58a92c3a9253af4b9405ae930b2a791243737b3d54564dd002ebb2efe86b7c50eefc817dbc1b41a64e662024a685572094f7d514bd67e3c1979fa8186ee7fe80bfd4bca01898e325bebc5f418f628410796ef823b8e70a99aab6e62c80be4a8b8e260014f9da7593cac43966bbc5dc59818451824960772f8e1fa334016c2afe50a7ebc1eb821d6bfc4c3e23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hd1affb946d942b02d8506bc0a1b70a566615c0c7cb036247998fe013f9b320980bb20c510fc9212c89b8f12c4f056dc308545df4c0c7d282f4fe9fa461f9ef0ec4f09e069b9aadff5c991cff6da05cf2bd12440de13bf477db5cb31a8c79ede83206c29437e48350b916d55a399d8e65b8bff72a6487eaa17f4b9b41bc90ac557e75b8d2e1d0e1f8b7a54e98eaca732411e9f6690f28bb4682c6b75bc4d4bd3aa047b347d4113ccd8a9040afc30089fdebabdd19f2c50ff5c199d740102698cb9caf12eeb855561608114308ed01c762748ef38d7458cf6b9df7650b288c627e3e78dd11cc1e873aeb4ecf8df3c4f83d71a95d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h45f42c72a229e297874375d6ce9dbd687d2eb682450f1b77525051332fd7240608f956d9108cff497d0faf1c5516a01c346baf417f015f68d570c993725d31a85a67f1f019d6b1aa7602cf63d9f33c046c2205189d3bc3c98931e0c9a04a72c06957f6e8d325c47b64e9675e9463de64714f228800405ed73f0f827fddc3dd9de93c4d9777dc68d1a1d68e8f2350b0303d71ac91454e06909fce5f239d5dce155d41478667736635b0180e219166835882a365741c215fa429b20b9dec9a2da9503dc9a690923b4bceb677d643e7868792729ea74bf0b96538d9b12f0f26f5fd1e24015d4b23a4a4a5c0b914adf23b9117cfeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he033402ec12b41eb897c310a6d9451a9913af3a3f9cee1bb688280a24bc9429f52f3dc581193ed4e4ffd880ffde0ef35b790063c2d735a57da7b49a4719a8753f59b071a86ac1cf9d040e50b803c2a2e6e2b74ce0e330c661923371c1e8cf347e3439513edf11a65f02ae0639ed7ed9096df0217fc86b1c3fda696b4a04adc94276348c8da508095fe0effe7bb593156e3556604fd56c36a6449844d7ff5b059437b4ab31232eefb5e1790e9dc07035ac1f7157faeca51298a706d2b730dd5721e7e5c939db425b40205d95b02486f21f59f711eba1f96b380f8686391ee99c0504214fc47d7d51418e3f6bc1d580aa3e26471;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h2a0dddbc29d0a2c2d22506c8ddc879c5461989dd1bf8822a0727b192b2b460510b8efaf66d0a36031a233cf44c8189b0f81e7f050cb36c59a5a13ae7f1079391e013ac47f23f472378dcbb63be100395f4199efaf991117ee2945727623907d38bf06d3261238b7304321803111d0cf1047a2d606bd9b0b5e26fed65453d39fba1bed214b17f5ea70589cd9dfbd22162da8575b0bdf6c42648e7b11c676107dd38e70887da407dadd97c684868e9482da46aae93799de600000f411d0801d3e46dc347b479802b2614e618f06c7309d59687f80894e5ffb4a3d02ab8099b0d0753fd72441e1fa2ce7e4b0f7b917999f9c71663;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'hba8e1900883328b9255de300e7887cc7c6bbe644cbbb3b4ab7189e57ff4b74385fb14220581007f34ace931cb32d3c977e290e3b4a7f22ed300b0895dbcfb186c065955977d00f33805f0988bf6944a1e942f4487be71395ed7525b11a789ee34179564de75bee77d15002d2b07b357eaee932abd03b4d89f54a92c7b1215d956bc87eedeec541fc88adc70a5d2d8e93141b59f55403e8a192cd588f60450de3f97480319e5df1e3f6c8c3e7bb62578e438a73c69ac0d734bc149c8d5d9af6e2eb1eb3265de886628dbbd3ac1b5299e0eb6353f25efca2c2faef0644202ba2a2033674693f93f5724966378ec9007b6cc3fc28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h24b66e78ac361a056b8a5d5d7eeb2931a1901a7fb1bbad50dd086aa50deb5625329af6960fe53ba22598f1b5fd3e784ab6528099db64926d90f3db43c5d6c5daf45743261a58241e591a453841a4a98b1fd2e1e0229037b456545a8c610e9545a49af05d89133eafbbb902c0d8905bd42248c41368a55b749ea67eb07a961f465081ebd76900554d4503bc928ee97b07742345d7d841978f505fe96d1471dfddf46ddd62592aca5718af5c753be24baf03f8d8d9474a82dfdde7bc744812aa596f6881e4780844848f729310e2bdb9fa15d6a378f98473b55e25916a45feb67db52fbcfc473bc2fc474700bddf503242bb840b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he20c8305b5a41f2666b8bdffd956b1e4e64c2ff65d6a9035b30205759dd22907035d7045fa12f3180bd39c953109e5f01fedd3a2248b5cca4d470b673d288a4ab03a1661de09ee241ce46f6b0c045ad3184d72644d5c7cf1fc6049e9a199f1f74eb5d77eea8893bd77d3d1490882653885512a23fcf40865b244386052475d76d2cf6dffb06623c3c6f7dc135892107bc9d7a46025a6e510f43ce1de8912d419f32a691b219e0308ee2ffa2b90993b35670bc6e1e4e8a58ebea89c7e19fdd263eda56fd8c1ec6a2d987deabdc96a18d60fbf06d1bb34fa9dc23493c7832ca32d1f28b715addb1f544600fc4080ba69b143cd84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h465474bf2ec9ab37bc13afa24d193547b7889fc1a33d5bd520b0b36d9692df20b720b93599bc1988c5a6d5a346ccd6b3a38713858811ed1c7b04211f2aa09ad76e21d0a1dd0328b6ade8a244fc2a8602702c7512af9cac8abd65cc29794fa44d2d741be6975220e85412d61c30715e1a463716d9e02d7348889262309e3ea8b7f1e56f8cd2ef6a9e701f1606ed47bd56fdb7471c839c6cc08afc9a28cf6cd81728c31ce90c8bf08d1e54272bb35bdbcc63913f3b797b9285c33b3f27e162b95fbc6e67ed841366d28fecfae9f71416dbd5b3c8f4fc0fef0e4c04c5d395acc3a3a61be8131fa89506d6c8fb0473dbdb61610037;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'he1f4592dd8e4b9382dc6d12dc8809c8f29435035489fd85fc6a8533594f0d4330045e00091ca1b109e747a99fd4a3b1e62989c19638742ffce0f6661389fb30be65ae3270330e9ca859b3da6b4ffa7a0f1af84f0891cc0a95bc39651904fbbd95375e64b19c60aeabe62981aabccbb9daa5eb57db38d078f225998c7de999c3b7ace27cf4d8d7ccd14968fb7d8e95c2aa0b48b6de6e6e095f5fd085be27194d788e14c31179d53512bbf6205356b91179affc0ac9968b9399c5b1e5238dba9239dc4dd72f7fec0cd21410760d2b346a73b053679e2eb28e7d0d4722a4f12cb600581aa59e151a03125f0d91dae913532be136;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1944'h826a474ec92b5d89d9f872b83cd78219436b8bb76dbdd518f4c805ec7bfc3a169dd6b7e0e99741e46ec04589ef0f3bd5c9d7c693453d93f24f0a2c596094db0a0832b7fed324bd803e6e660fe96845da0f096b57abc8e7616207875ca6a79e047a8ad4538ffa604c75b3af0c8a57df3bf8b39e4679c3a806beafe27e46b122277f042670e0d0d6c750a41e736b8777bf138d195f0c2bbbf154b8d2575b7a6f37a9613fa3e6af031cdcb761c3aa9401d760006a1674791b9d1b27e63b5c4d85f14f7f8ccb8bb949ec842ac7d8f56575aa7cb003298bd3313346794f1ccef9ffa1942caa74aec3e1598f4a0c49aa48ed2190997b;
        #1
        $finish();
    end
endmodule
