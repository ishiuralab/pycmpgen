module testbench();
    reg [9:0] src0;
    reg [9:0] src1;
    reg [9:0] src2;
    reg [9:0] src3;
    reg [9:0] src4;
    reg [9:0] src5;
    reg [9:0] src6;
    reg [9:0] src7;
    reg [9:0] src8;
    reg [9:0] src9;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [13:0] srcsum;
    wire [13:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfffffffffffffffffffffffff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b989f08bc1c9df358c5bc039;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84ba04f95c7a1ac878cb54607;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he47aea3f6752317db104feb3e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78e3ed2549d72f04c73e70bcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h701bb565318ab7e385bff3239;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha202023ec5cc552232d39a050;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he92833eeca65be13484532b53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6f14130c4efa6d6e37492e0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafbfcef960869154867427fa1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf2a666b7202512273b90ac4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd9181d4e09a672cc426ac1f4c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5912215e807e506ff56b9df8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b4852d2f8e30e1cdb209bc99;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4768b511a027b30f86603d996;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68696f1d2404edd531fa0ca7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha905f462f72c024837eb9eb93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5d437ca3bf37a4f32808cbd1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca1b8dfc8da656950ebeb081;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4c783db7dcec33d1263311cae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbd7275282e233946cb5e5cb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac7de7604a97701a614934151;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd82a6d2acf8ebc51bd0713e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f802b7c1d40a7a570db66ede;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9daf20666577c3e02e4629a4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74aa35e7f2f5555a7bc516c17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf472a131ccc967764d08d15a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f5ef40e3f1eadf9de00c3132;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57cd33839bca794f2b3a38279;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd82c9cc51f53dcbdd087de7fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8939632bbb69f1d92f9710d85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h71de4e379787c4ad1b57f794b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf113fa60d14feb0a6eff755d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd372e7962532719f535e856e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7dcb0ec68d19848adf85bcb85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49e123f577832fa64a0a73f17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17fdb48447fd9c754aaabf034;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe46f236643877b2c03087836;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcac130ecd672876ff82b1c05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e8a1429de15083c3388dd7e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d8d25806687a9f3e75a37b21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86389e2478dc2ce645ad11364;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9ac0d27f1a7a1859baefec1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha987ae065dd84f4b2369dc5b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d94a9015c1607bb77ca114f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78b244279ab582a37faa0c0e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h861210685300feb87c80fa984;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h909368e35d980890a184d93af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29a54e3bce91231f4923c2286;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4fd52f39837ac605e1f53d3f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h574eb192b9810c788c248f51b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1c9139103ec624c4ab359b64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a1a7394ddf713718ced1d5bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5a14dc14c093f73ed2b0feca1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hecd42a44ecd4917d181417506;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b058ac3e4a996d6ea9a63591;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h960af49e3a0683eea9b4a0c46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf51e4578233b3fca6a50a2b9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfdb58be3a6636aa72d8325f19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80f15818c663f0a79627b49c5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha71b74b37912af82a37e017e3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h227e58117a4e6b1c81eeefe1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfad9a1f15b6274ce63ef59d20;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1b35da599e3871e7669a93f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96ea172bb4d8b118e63eb9366;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62dbd17ba3901984bb6a6565e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a2926c97b332c85bcf38aff1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1fa5a1b4da114d6c3791bc4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98f6d7bb6354ede992812b5a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90dc2538cdc6b20a5866784f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h314d9254f056e9da875354bae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h119a92cb4ace79da1648adc3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5747d16670d310239e2b405fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf7258273183a9442427b4df4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54d8105f65c677ba00e71c37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbc93a0dbc0e3726a9f8f03bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h79996568668350b2c5392ef6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84ec642bfc321ac869c1b436c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd135f5857689fa08f3d452417;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h624e81739538cd702c8732f31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48d4477c493b645cb1083a671;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h966d51be9e33cc01bbcf6b621;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4934872c37408081dc01c79db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h512d00d010c64dc20437f6960;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9d746844c6e398195bd31799;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fcd6d90052c1238035d52e54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec15a3b1b3a73ab4b68b67af7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h804a9f600e881811359dbc834;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56fb6ca90acb7c8634ee4d5c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca3ca15f8bcc08f72700c5679;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21a3296c834989d83ae24e358;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c9cd727bcee191de2a4c446c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff591d9925f31fa29986ed3e2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf408bacf267b6cb399b03a717;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h727e2433d9a4b4ec54b39bcaa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e29a6c1a09adfd5ff57f5cb0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h676c63d49325d869eb43b78c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4ce745e203e3a30ea31a5badb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h626f8980978b1842b3df692bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he66e679de0f69c94b9eb37433;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c8b15386f8f684c8041dea2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2001bb0a110ca1f3afbe13490;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fe2a775ef964500445b79416;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9e6959cc625067f2da8edaf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11c8e69e5893681859623e5a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddbc401393972be569ba1d61d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e2f987d10eec8caf891386a8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b6881a4b825b5cf1264c982f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hae66c83ab6c0cc7bc159f45f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb88e3be06190502edb88e4c54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68fde33c561aabb1fab137e85;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc027110dea8d910fc8320f1cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb85b9844db9c8c6950c0f23b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96badb0fe7e822633aef24761;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70bc769f0ff860a8a0b560e80;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he70d2f487d13b635366a99897;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc0f04e523a2aea7d45afaa20f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h51d7a08efcdbd5b366e1f5f8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h165d015dc07dd8a7e3a174e28;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4930ad3079494b96dde3a7573;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5778f8bce3205dcae90ade0ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd83f38da098881daa54d218fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddaed41d0a1a4f66188cc14e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1fc14228642d1b356760d5af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6820f63120dbe90bce88d83cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf14d28410e6502aa49520f1f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9bcc0d7857e7ca3e010136af2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5eb61c56209fa991df98ecdbc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d125060004ecc37629c8c314;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcf9c7d3825c0570391fcc72c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7dcfcbbfe66aa9c87011ab24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h725b808b7ffcbc80605a1a7d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c73d666e0543254f62056b82;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he82c0d00fb46125cfcfe71e86;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b88c3a5322c3b8111e2feaaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hee1dfb9ca25943fdc0f93f646;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24c0f37e8ca0c252d1583c570;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5cdf62fff5b538cd608263ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8ece078df4db98c7e4a97f23;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha086e9a86fee501e32c2694b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f2d6ec7f1f55d176f90b672a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b7d75e5e6969b065ff0912d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc6f73c35c058b5abff7cb620;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa8cbd4dcf5cb101230123649;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dfa41eb6c18f26bafdcd696d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc31ef556dd50385c44c8ce90e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66bc37c6eeaffd94dff9c1913;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91e38eb2ee7b343b0bb617a74;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hacd3d4988fda48be5a7b607a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7e27f257443e0bc0b8fa5531;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf980c42100246eaecaaad6ac4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h376e232ee544a509f3f641fc0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb5a1678888d24f602f04bb3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h514a000d476bf523e661fe11b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f9332316331e2b63237e1404;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbfdcec9b454537159f0eaea7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5490a608c59da7c2ee2aa33ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bbfdcfe249ad7bd52440c7f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52734c5f7d3aebc59d3b45ee2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbfa4449ccdcb1f10eaa25d710;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h355aaeec52294bc39d7ca1292;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2beea4d19c549283542a5b39;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9819c4c9c8c9d7bcee68da7ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e18ca5daf2f42b856d67b170;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdac40eea3c3f2feeeb22b049b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7dd0f4e86f876ea7a34d65af7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he54ecef032aa53059941cf077;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8caacac276cdcc1f984007f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46c9a52cf3371c56358b1d72b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95480ec834a2868b7a452e0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc08d1c8c52e7310533483f537;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha83f91c70ba28efc295f13bd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd90fe1678df9754976fc4c013;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb75c65c10d84b3f7a8d39eef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce8751ea18b22a363a5b08213;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19dcaaf8970dfc9d8aed0b0d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3240ac23c79f20be7e77d9f46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c224425d567ba39ac030bda2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha1d8a0d394d35106760c16db0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h280fd0fa66bac2b950ed3fd1b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4a0de15e412350be01d969e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h536309b273a8a31d1c09f021;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48c6c9b81f0b2befbaa20fd3b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a3d200af4635b96eb17e6c44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6c544c931050e1167868a0fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb56459b9954079513ea323af0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1eac17096fc4d7f805946dbea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cf33806840c4c8eb3409d169;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38a5c66100d57f93ec69e1dc3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43dd3ed7b61a564953bbb9f43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc899318fd590778affb65d4c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ebf2a37dc0fecf0d11920724;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f36a51e860e7d46d0fea7e25;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35d58df5e5ee7aa52b990f0fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb8b8a79b83ba9b9869c7f7ee2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdbd141eda8f9d7b8eed3831d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfca81283c557bacfd8b49662d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h98bbccac83e23397620c8471f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd41ca8791aa3c6d79e6779e00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f5562327ca07a13c591839f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d28c99688ecfcc80897a8b8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfda90ea42dbc6df2642054552;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2bed7a3a5c002fbb87df2d22e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcef4b7341828b876b3f6d6407;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfccab4b28ea25df8274ace61;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdd19bdec0f2985926726ffaa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h311d239f7fca2eee652f0ea22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbcd26abbe3d6aef365167ac1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h792ad946170abf8caed6ddb3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57489cc3f33422d8276401803;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fedea6e2e17d827b292ca966;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h626336ab3c723b22341b470cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2eab9725416c9e280284150d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9f940940cb2aa8ce4d779375;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb4c55e39ed6ac61cf49573f41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea8fa000b70bd873f6c454778;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff2ba8ad3034dfa5f54916c63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd38764fb36a0a797e27f402ca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9634ee4708c225fff49553c4c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ea713edd28fabe28c92c6086;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d883ce258948e0bcf4aca2df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31c0fb5df21cd9e7afaf4a03d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf72dd4ae858e77476d7e7b1fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h825935c389a19e075528d5bac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc435416af4dfc938f1e3b1cec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3b352180edff271dad32e7ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9cfc7f1d9b1c52565e4b18d15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h817ea36487c6322ae8152920d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fb45a2f7b00bdb86f7d9b4d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1dc4f4347cb5b4c5a6b801804;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0cd3ba4279e4ba51613bf95d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7d09df6911d5ad1264843be6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h612a0d490ffc5d382754fad15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc2be8f15c112b26a838ed0a0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hba4e7ce4be8f60bda73b02645;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dc0092ff97fb7b31b8b05e51;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h80aa1ede5092afc0825241bdf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75c87aecfc89776e948aad6ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had54e1b36c0aee81c479c2a63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde6c2f8d26e8f3e717a677e15;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3a219271f51b7c0118f4b0180;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1d39c76ddf5fcfd5d0fb31f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e452353d22bdb49ab3af764f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86b83b2ff8c5c99473078885d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3d4cc18bcb6a734c78389473;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d14cef87d7a85ed2449e7931;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haab87cb098c769bba37fa73e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd569acfbfeb7a366d9b3926b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb3246bb65e52519af2f9188d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf47a873ca1f700e9dcad56599;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69ca8e0593e14ea14f5b1a237;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34652767b4c2b442970854caa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1f7cf7cab46333234d7d4fe8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb5bb13ce9356df60db19e3ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb875e89265e4fad8d75eddab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5ef7e284b44b24228615cd985;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc353a272bb1873f419415a251;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h805853cc90cd8f5b65dff658b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4341dca9d040ad152dc5791c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39634a226115c1fd0ee93261e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h178a8388c50ec759bc10b1585;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4dfb8b6d01b0ddf78a4b231c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c454134fa67f7f5498b0d362;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc982213daad90b2968c865064;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48452013ffeaa7c040ff4c7fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5eba9f67e5a99bdb684fbcc70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26c77cc514500593d4e9693b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd8ace45544e4b0dcf6033d6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he12a36c1c359bc3d58eb55b2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3beba41e19cf4a59ce8a494f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2bd8d23563d05c4d299202fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf68f332543aa0d8924bf9692;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h590ad25df79856a1369191712;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17313c96c85a2a2e795992518;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h22c4774907f6dc94f2918a658;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9e59d0338fcc90065d4516bf5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4d399efc967695bababb9b8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa037fea82bfed3ba6e938147;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3538d9b584af20c900e65b5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12f36ddfd82d591e305e9c77d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf16e8957e70a8bba864a9429a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2fa8fd7dc2658cb195dfe26d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4a24b3f0274ff52a964da087;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbecb1509dfce2f3014ae4f91a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d8b9bd713f5e95a7c9ee678a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he367b8306ceb704ddc3987697;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h792ae572328800b6e18e0f30c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefb8408aedbcf55946766f392;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde49946465fe71ca083ab6189;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2007cc1df02bf0d484aed6227;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb64e4a844e85fd55c9acebaa5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdd0b4f614b1c9706e6d947ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6963430def2c17138ad5e337;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h524cf37b0652ed4f5307b25ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c66f0a5b2f0a5d54628b32e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f265e7f7d9f282dcd85f7853;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha82b9fdc42f6313951de289a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he1e5ca3294f66dca1d03ee58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e0552aa43955a4b6ce47d9b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha260905f238f5ac9da44926a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd22258538c709be7f5fe785c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c8bb0e9374f1f1dc146fbbbd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3924dfcf2a97f9beb04b19d13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5685c226206d7c08832fcc33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c0c29b9aa402df023d8e5e21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha183b622eae8de99d36c9fb6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5675556749ac3f54b1420c452;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc642e6982425542f87099cb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3719c71ee894965bebdac4c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f54c66cb7e2bc8dcb16938cf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2f9d4d5db1643d5aba97b289c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8aa73027bd20ae929432f21ef;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f5088f2b7ae1a705f39d1f08;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h78c078295e763d5a9fbcfe2ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf391cb0c56cd266c0d2cd272;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9635be50912bd12d36726a715;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d758f72652f65b10c79c585c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had395252f764fd708fdb6c487;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h226560b1dda097cabf1fac886;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h35d4cc24d55973c9013ea652b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9d10d2716902f93ccc8cb0a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc497de9ab8eadb3cd461d5ea3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdae12213279eacf804bb6ebed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd29238e14ef83c708b2ccf3d9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fab95771c13e22c8ffb07224;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc8f5b2602bbe0c5f29aada24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2e6c5b6d1ec12d3c357ae93e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b2b66b1405fb7d066e14b2e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49621535966dc47c3e044e699;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b51c486586cf4058778e23f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a37775ee569d2a9c4e28a090;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h370eda5c00666ff9e3296993f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84a97425fe37877c1e4e0518e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf827c0849ad2562ac8428219e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91d8e2a396d7e0c4acd43dad5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13f5e0cd6404ce661ffa0e1e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4613bb132d6ca81769bd58a27;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4653bb09e1d57004c6afee84;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h47e189bf87082246a8d48a8a2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h695f7d7a5611613c0a7bc1922;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h217e4cad1531cccad9f490ccb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6ce600319290d7102933a446a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cbcab9827d89818a371fbbc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea19fbc37d8fe43e10ad7afc5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c3655427dfda5d2c77d86f96;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbc4f563780cd57d907b642388;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa9840d0d1c260159fbee34b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf723d68a7bacf7bd0c0c54d4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8eb59af06ecde08be550b371;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9134d9a3b6b02136e7daff473;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41dfc44793d36a9dd2afefa41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b8556b325502a75008a66b8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hed29b1a37da431adb9dfbf4e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b7e41067bce47c227909b106;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he4c92da86b75f503d620f2167;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he84d3ca603e716296eb10a6d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9dba4c97c273cac640630b55f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he531699de41e9101663e46bb5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h874424e1ea5fdf051b6da617b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha14e9490d884aae8b08941a67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce3c929130ad591051bf19619;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5523171c68ab8154c69e00d05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcaf8bb336b9cdff102b1ca11e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haef75dc8a2174d742c5ac4543;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7cfd70a53bc772e96ed36b34d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf59c51deb7223d0d9a96c453e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ee10f7551e6a329ec49300ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b2d9778b1033583a60de580f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3f8f64bcd6d544402c895b7f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c5aa7e9a503fb8c0b1ee5a44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc2acf83267207a259593c0f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc092fdf54835a0cadef9e52d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h571feae3809ea92dbe2541595;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2b93865b0fcb8e6705b5f7d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he92e53a40023e987cfe566827;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73e804408aafd6f104c803ae5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7714d8ef57053021c45a06a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h523a14f28454c206a3f601952;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h336bd647d25ad60612982000f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99eb7c9e3bb6122af6e544455;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1aa9637863d602033e16e242;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8df8d5a936ba4ad3039e2eeb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h384ee8440793107770628f099;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd78e57efea1e4d5a020af800;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h12f52f6970c831bad07273725;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3899c90afcd4a16c3efabab36;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68df9c1c1a12ed184cf58ba1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9236f7da8d2bd6565b10039fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70c7c2906293372a0091da6dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75fae56a17fba28477998850f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cd8c9e7359a0569d0b346445;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ddb987e8144321a700d7893b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a96ca9ede533a9b6b73b5d29;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcc345a1ec688d41204aec986e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9947a35d024c89da6604efe12;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e7fef50d4671dc7b9a6cb352;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h29207bf6d4b0513c2e325b55c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48531b0be9919538af44176b0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha31d2664a3d4bbd93f44c7ff3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fb0d76ca70c026195e60418f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66ed580fe924ed1ad89138851;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h69e2d110fd193750204183f4b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9ba34748bf977219eaade0d3d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdfa233cf36b1696584e1755f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h262028dfbeada11d6656d3995;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4e64971d699d60333ce7ea12e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h41feedeb0ac777a5fce963f6b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3549524eae56ddb99ccef82de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb050f2abf5e557ad4e02a0dd6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda0f15a48bd67f655686f4672;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fa158dd1aa7614c1348e53c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4b15dd6560c302f72a457d5fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h785623c4b680910681a01272;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38ecdbdf75070e370b3c13ab5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ed7c5c503e86b1e88fecdcb1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h233006b520b799ddd0c361a6c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hde54ccc9eff47d877183f51d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb39c6953475ae0747965469c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h52cb20c60f0acec4a2947a65c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b8660170222e12b38a8ee5f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbef3fc3d06c5929e5a3b2d12f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha9126c58917154ae2f65ff824;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7829a1775cf4de4609e7d21ff;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd0e76f1f0cb11f5a6670cd37;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he53cb6a8b67fbac581182f86c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23a19286b03ddf218c5a9b505;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bf8bb0aadadbde1547a2ddc4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heba7ef8b3dc60f04a7e3c36db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89cd8bfb94174a19a320cb247;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h693acbd8e595bf11e48f2a8e8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3efcb949d6c0641b432122a41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d860463e475981544cac9d93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha5f893aca84afdb18930b5b58;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hefe411edc77f01c310b35499a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc24145f88af99ea60cc45c142;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdcf16102d8c7fe9492e3560b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3cb378de942ca3b0be8050cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he00f85c2dd5ae1d15ea071b72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ec1a2de81ac295a8fa225beb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc371f073531d27e9a33be72fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7405a998d43119798a1cc090b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a233454288992f5ef33e4e53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2079c4896cded0a82f104cdae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h695ef21ccf4675c2211cbefad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h133dd15ded49b81f3f1364cdf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce86988f6136002e318e546fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h55019fa84475efed7b5351639;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1a3c8e63209b51fa36768d234;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he964d575746cd7c518ebe34a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd87d965874b09f0265eb038eb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6972c24653c56036dcdd052d8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62bd9506392046726ab01c348;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h649589904b9de3d2ecf5eb089;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcff4256d8f8e4849328c9dbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd58391ffedd7f3fc5b82bd7a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf0b7230ab40644a05eacb436;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8be5acb8a3be2672a9e674dc1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h77e7af3422c829b67a366ed50;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e5a9bdd90e8fe95e11bd4f0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4aead917e5478147859c8c6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha79849bed71b8d489f3386133;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a00e27b02f74110636dad744;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40e64a3d37e8f1e2b098a7ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h810f052903d385327ecae06ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he47280454b5f7b6c6dd18624c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcdc56c8122ace27237cb5d9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40d89130169e0b962e000e030;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaa22e01de633c399d076cba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ef22188b60b99d6ca9b1e7b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he003015eb0c2115d7954ac01;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf437ed895246005e65fa3043f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h451103ef7d928ccf98bc4d0c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h19d56542c837528f6a7eb2871;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1c1fb97847642fa4a5ea1066;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37cc8dbe8999762889c2923f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dff37e83a140a904c8341e10;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32cdb05c731b5cb1a5b7e5b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6869d6dfa8d92bba879adfbf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf15ea9307b7371ac5afd7fbf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he108e4587302b528a30e248af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc1fd25638d070b695fe9fca24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h345c0373a4fd4086972a1a954;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b34a346943a0337ed02ba633;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8dc1c2f7c7316cae0f33a5e66;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h363cd1d577c44c29300c62d7b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfe4914691aac118508c6b566;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h700a50a4766f7bfc9ee91dc30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h893c9e936c1225ab9b77f6ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65b16e82d3aca8e09b5fc44f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3680fe07ae5ef5215fa261da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h995250338c995ea61fdb1b97c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h190239a8ff2517e51b4090b21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he88ffd3fd1c6814d40de0fdd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hffa9e3f8b61c1d40a04aa3aca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74937d1d6dcc83a775feb172d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h13a16a7f1c75eca72c48d0f1a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2e6cfba9af4d7ba56cc0d4dad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha383de19e19b8c8ce6ea0a7e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbcc694a748f59ec56418315aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea6ecb248cf288a392fcd652c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5046efe8f0c09800de53639c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8e26dc7055efe1e977d3df18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc57d2523799d155f1a74c8f5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he59f4f287780bb91abfe18a8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf85115e9bcb4cf502fd388a6a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8cd178ee3771cc4beb2295a05;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9239bf0e53752a817818e13;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73bc73158322b543861dc0454;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h130af6c94326418c435ff28e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6fd793b7bc4861ab6f5dbacf4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fcd996f46b7695539f5c3787;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40aad42610c154f76c3c5f68c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e0e199f61026b4df70e8a7dc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20b37520a846a5b61dab6f498;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h152a025e4caf3b7c750ab2bf0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c53d50eb8a927a76e4b706b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d3cf34447c880a1d6f3ba2e6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h27fe5fd75c6fd7574dd008259;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a786a6c1e6a0450b5f6a1383;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e2d890674494ce98c703e228;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7bfb20612bcab566695b1bc23;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h765a5502a85cbd9e6cbeb4848;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93d25eeb59da60b7fa1998d07;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1edb1ea2590c3b9adba89c13e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he464428c06108352dcf0d19d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9fe9a68a5457522350dcdfb00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h156df27270111b547df9dddb9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbfd4c3d2e4ce755e74d4939b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74b6e0565add7761813c75666;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd165c161fcfbb93544291b5f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5976f61802141388910c3d9e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd6081e78e18acefa944b9de5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf791b32abf86112449f9b7a3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h931f91632a286b13221ca9e7f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbeb15ad0ed41de67baa66e76c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb540b50a4de5c4d13cc595147;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17112096aaff444fd1663fd18;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddeb8211cca9f296fe9130b8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88ec636664d06211553bf969;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he132cd89e7c66d365a7245181;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4905d464a31869a16cd987f3c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h25e03141c58a2e7985061d988;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7aa0b76f94ba9d836cad7378a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a2b4738099ac8f72a0d14147;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab2500f0616b00901c32da415;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he042ee5d0ea0db2d969ac6a33;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb257b656379a6a0464d29ff35;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34c0751b6d18135839d3e79f4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8b8483f96bab8f66800f2748;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2598fb134367c110cd5d447df;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe8c5580e4d51ad63c59a58d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc33ea237314ed2387fc72f2cb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1ddc4430f16c651106608ec19;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h625e11ee993afe23cb4d67e46;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dfec90c0e57d0c2a54b9398c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34b80d780bb6403225a1a0adf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfccf429c3e8379e410d2500c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7b569cd683a26052c76fa603;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha58561488667868bcf2fb66f3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48a2df38331f38012473145e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f62efc7ad611e001c6889345;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf26045e491fe2eb2ecfae80f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66950d43ce2936c90db2382d3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9144faf1f3fe9fde20d5a5fd5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2d01fe487da1504af4bba41ae;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'had90fa8dbe2b6b679da1514a6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75e46d8b6dbebaada7c7a862f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd73e6070e19d4ac3d1d394d8f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f12c5fe1de16c39d79427f5c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfb1085a76785308e0817c5a6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf60a1525ab94671df0ab7c07a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha3babaa03701565d1b8369b0e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce2e410ba4c2384ae01711594;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cbd2ed6d057aaa5c8ac310d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8851d38f13982f0139629253e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd74dc91b315bd3493cb57ff22;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h696d1b9847f2f29acdd33007c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h518ae8f8e80cabf5a4629f3a7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2830eb5bd6723f0799c484f98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h166d7cb3f995c934baf9658bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb1cf038b3eff6f62ad53818fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha2f2e20c74f250901f75b1e2b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h46e6ee2d9779594535f9a6d5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h501671700f657e9f146f366f8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha791b4e0e671a6089b32bc1ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c2958906988777459b0c54a5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc369b9e866204c9fe72e1949e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64998b4a635ba78d43dce3f89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b2fac0690acd04ef02248d5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dae21eeb9257e2717008df3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h445f39ef210ef02cc5ac257b8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h324f397dc4a769c05cb056a92;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96cf302199773ef84390583f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h262f3822cd200f7b3d023297f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3fea105d8422dd9e5ad47fb4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcba8f01d3efae590def581aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33cc92143260406fe2161224c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3e798fdbb101afec478c235f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5e59e2bc5bcd85674e724a716;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8064428d6e68c8af0a5007ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfc45e52e700fd24c054b5770;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha90de667211bd79537fcbcb91;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ccab728a94325b43c393ea9e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8d50baf0da78ded17065ea984;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37389a52df82b824c24ab79c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda0be10a3b9c738db3a54f2cd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hce6eedb78d1cf769c0978a5c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb599ba8bd0d8e2edc33b833bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b36ed9a70b4ec8244c6c3f5a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h718de28b22cfb0501f44401c6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h352b501987b4322c629f89d64;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18824da8b36d1c6d9f529f0bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf379d436db2e68b0011159c2a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef770d3390bc87d284ce3058;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1496fee9d331372f951287fe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h614772ec904f13f41aa0333b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5839b3b9c83710aa926a21d4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7d02c3908828bc9098b042c03;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb377d896890fce8e781d06664;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h346d8b45d0ad82a14ab392107;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he78b11503e95dc285a435b2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda8770ae5e867e9ce3fe2355f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8aee85786682fc4ac611fb92b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40abdb82e8a947a02ae54bb2f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h57812377712c2635bdb3c95d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6f9117724e49ce09e41b229c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb129cf29f17383f106a560aec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h465287dc33e81d09807440153;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff4d1571776678b4c765973f2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6635eb94b8de0c55d40e6aa0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3e803c7c990b54f7e6ef9dadd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50d65d30499e9a1a61bbe0f5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0d93d20738aeef692cce1b09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a73d837e27cea4311f173439;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha45c0899aca37a0af7e7999ac;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb5e97661639e6751292462a8c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76291520e38c7db190c1f78db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1743463e6fd80d545828d96ce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf8223ad51abe7d87f33190ebe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h84f65d9fea7365e12fc9d0db4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab861a842c4226ea52ea30160;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd1aaa28525af40316a2081132;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9b3547880301248466b4a5251;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d876c298f5799a27427d8f7c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cba77e61e243c42bd2f599f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h592ff16d968880cd171027372;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddb185decfef8a4c652b643f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62543d95f3a3f87c8a73eb5c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2dd8423f32b08b7ad8a464e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h969d75db70c4270a6de19856f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h421ba6cab70ca0505ecd2b1b2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e5a95314d0c200147b4bbb2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h968bf2435cdb17d865915683a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd12c43359754232e111e4a5de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e3403637ee5a9c630ce86b4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he7d3bad1b0b897b8405d02767;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38c1252e2e049bba497c02af;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he227715e0fa3c09fb15f78ca3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdac15df3d0d832da3039111d2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd6e5db98a1ad35807205a0320;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4711dfef37731a99c4d1af9da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda8b6365ee8e14c935b341bf5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h277116ef4201fccd1b461eae3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha97caa6d476f537275f729587;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h49b4f5015a764c204524faf72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbd5300d0eae8092300fd8ad0c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95c33d566a9d1d3f2df06069f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf811b4ad875f461effeb1685;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haca75f1e2c591eb063fb75f3a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf870c83951c3077787c96eaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe7093cf4bfb3bc2027c680bb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23fdf60c1095715098f57acd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18ba529c55d4c29c991a21714;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6eb6344f4123d1f4b53dbb190;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heee9c89f631cffdbb2a6fed5e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h799a7bc61970ac2437df67ab2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d3fe7d1bdeac12b25e422647;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h920e163920328ad8fc1924d77;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf1cfb366f1f1601d255114e53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf29fd23968082946b999aff4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h864396124018ebc6ba0b96c9a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd8237b3fc70aa0e1b227665c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heeadf80eeca7f4c13599f45f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h454c3ffb98e75e6b39ab6e03e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h32e04ef5bad1879602586e72b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26183c912206da4c0256c53b5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h54a27c91fae650ed42108ffba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcb5b72e36766c5737a552aa63;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h890fb9fddb3389606a4db40da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3594e0ae19724d1960fc9092;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h596a2d22d7ec90f6fe394056f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcda7f775eee2ae3f19334cc7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b2ea9ae23598547c3b69a21f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haa08027778ae763193f354a0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2dcb8c0fefa2c76aa9a084bbe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8f6464ba98cc9ae9d49a97c41;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58a2d229cbff914014bae90f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h639d1aa940882816a17d4895b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h988111b547457ad08cb7dc9e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h949234572ccb45d3b1ea8974e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe930d5cf27d7ff8d86286215;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdcbc95d808b351a127d472402;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h770fbc20663233a0b24be498c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h63effff775c6387859b004009;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cdaa78989a7bd32af548899b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf08cca14c76a83f7fb08be76d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2551f54d20c9436180d9d18ad;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h18b0bf34beb3d471b06b534c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7e7b36772cd18d294247b699;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h304e6d16382576174e99cc386;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a0e73a23c8ed227c393c6263;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc8f6fee2ef55b83392b522b60;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2ab93066c50021f69f685c6d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a30bf33b68dc6975c3891dce;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb921a0c0dd9958d072d0dcb2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7302aff688f2e099658a633e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75d308443d1692bc42ccefcbd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5c92dcaf9cbef604f952242e0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb343580ab4e18eac2586500f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6a7ca2379ec5ffb8ab01829c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdaea2086d542197524efc5d0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h65c2ad9957888ecdf110d4b0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7df31acbb4753cd7849a9cd17;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h592e1d476692a8406be11c339;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf0d6823c86344ae220324b6d7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5cdcd465f94d0c3fb372ddd93;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h689ab16f17d41c9b30614b0a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37d1950a4d15afb0f15360cb4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h24fd5ffb6d8e2b40d699f5ab0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10f729fe54d2a9e36f03f6ced;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h91b317d0d9eef36ad587eecfc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70f386ff669c71860ce935eed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf3c3158a80e90636a95907f2c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha18983b19629204c1d0addaee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75af73a071ebc415e4b79989a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc931f25d8e5717172cefd7d4e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7408a9fb163a5c27dbdb676ec;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3df5c1ea0a1e610c95e47f470;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hca75b9a656e402b4289a5aa8b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h816bba202b86b08e22434627b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86d4eca18a500d31480aaf8b6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hafb9381533fd3c2cd0ab37852;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he002bc9529c0f109df443dc97;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf99afc205b06b707f29ebd98;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h20a57028ad80c788d2f8ab73f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d97daffc912f972708ad08ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h75d11a270b4ab4a374a90c0d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5465ab0278a5a55ec7dd5506b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h433589c2c5b515f15f6d31007;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48996ba616d1a2fc27e39e694;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb34c332f6477f93775814242d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hff8af7d921914b70dd3ab91e5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf7f816d83aa438e66cccd8878;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h621bd22cb704a03fc1113bdcf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf486b2b7b639475159e97253;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h21031d4e45fb1fbe02846b5fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h17dfa8381d21d9c7705c39b24;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7f652e8bcaae2f44cc57f227;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h40ceee7758b51048e82005d87;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7e2d749442c5b1eb9e77a3964;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcf2cdf67a385f097eeb900fd6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h23f1833a0b6222640da95b5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b5db979d37664c0efcc72ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c17891673794e43680c9e3db;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11281e28a75d835190a5ece45;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h342945996651b07681cfd4b8d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5497049615d9dd500de672502;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fd61aaa48be0ffccd6131ac6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h86a277fb174e3b17e2c685ece;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf9a4cb6cdbd6b737c20ba6069;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5124dbddfe654794af1e58d00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he417921e2377390f232bd6230;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa25c25019c5e4350dafddbb4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58569d00b4ff54b44d0fc274c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdc6f8ee37f458059ba90fd191;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5dd922c98721c0fdf31e26d7e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h58c0e4f0636e41e403113378a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c60de9e0e53369b6600ec23f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3cb65e892034eb217249d68de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4344a121d0a7de4675ad42c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha08ba6ebf60d1f52b5563359;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h754f33203f0c5ea4d7b5cdc69;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1278b27ddc1f2273b2dbc7ad0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1d689c20b1f4ad02430e4afc2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h64e44aee23e994d0baf2bdd11;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h74ba5ebc9533122592eb09c40;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h732dac66541b133d5fb1c41b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab4f415086d8320f280e8c81;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2076d42a9df0a2cbef5260dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h584af4a1fa67519ac7d5814f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9589318fcc0b4808fd4346654;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2704e10d01010ac658600dd6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h685769b67ccbfd9729d10bbf5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfdfbf800a7c3d063637b91c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5474ab56a5c4c0326ecb5f21a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7700fc0454d32e49a1351589;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h36017907119d21df56262240b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6cd86b6983fe1a00b18234f54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf2e11be6d7723ae297e1ffc38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he38b9273f5a158d99422ee4bf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5582e835aec3188b93f09e284;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf3b2d5b4f20660b6c3c0e625;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'haf7eaea49475e9fa1d1956e4a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h48c46e330b877190ee165fd38;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdbe9dfb45f46394312ce3a8da;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h76ae3ddfddd600bb32a2966c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe25ded1e3e82f255746927ea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2eafc4cc03f19b69ed40f0355;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hddb690e789e1b6c5022b1ed6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e3ea42d3c8e9ee44bf592e30;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2cc03cf958cc6bcc738917062;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3342767d05d44e33098a50639;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2c875e34978a067711a7cb29e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7c66fac0d66b346ce82af8572;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4f23fce08b383cba501221a74;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbed5b8fb74f41ba3b21de46de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66d7a4845cb75f1eeaff1bafe;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda55bad40134da60ea840be6e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1be379cc4a7af4ff18b639c8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb7e6801f53955deb01f752ae0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he66753f6d8129e78321bd6e31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbb630d9c3531b865d6809160d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfe1344d33a0de9631db023d5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h452cf35740753214d001a2a6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h97b3930cd96d29811b5421d31;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc59d71ea71300afd2f440a750;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hea6bbcf573d8ea40189f077;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3078c3fa013ab91053dd56996;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31f81eb25bf3545b230558a76;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5b348f83aa6de55b189bf6807;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb6c0a7ba366d3a745649431de;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbde2eb07cea7a8a1c9abae597;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h59c67cceff4cc1ab01af43a3f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbdc4dc54a5b7cd748661c3d02;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c64e5fcb6fbc81032d39f302;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3c9ed158e4670d97ead840d44;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h690b30a7ba5f5eefb8edc62a9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1e6410849af8fd65db9e5148;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb2a3831ce7a0c1c01af8b661a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb3182b0a8e4e7783aebce0fd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2bac5922fc687540b8ff4f4f5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd79efe537ab702e609788cc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95c81df55b2e3c164597070ba;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h89d7ec2602e98b34bbbb3bdb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4a3e916654ef4bf2334aceb89;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8a34f62e815528545d012aa1f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hf5a2379e4d09604f0f0f20795;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4c8f3351bcb367bef8b0bfab;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb9736863bd5a2ff04fa808857;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ffc7d746c9443a59db262f67;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7237476cd8277381e3e8aa002;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h528854a08d908341020f5492b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b372a35cebbef6469cc2e34a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd3c7dc5543e57f4b41cd6873d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h569b932363b070416b7554995;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6e7bcaa201c9a29d82810066d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d47dcf497f81ac05806b5513;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc9489174c8fed4abf9bb8e777;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h62270d94c23cd18291d601d5d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc4f4a0879c9407127e41bcbd8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h70bea339f7b117ee94ff9d99d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72d745dbaa026d36550d17534;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd2e6c7620859f3bce603e9b00;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h72746669ece69bcc12e4cd373;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h67e8d4fa55ce3af2df1a8699e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd29de702cdb54e252f19cdce8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c03c8a3318be7622c4d7a1d0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f79b26c192326c658833294;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1c2987aa2df0923c74a1d6a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha7d68b806d46b70a23e6272ed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he0f9d9a8efb865136f036e451;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha0b1347b3dc72d77448d4eb6f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h96010634f7ab471af3d0c63b3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hac27ed99e8cce8e47ff2e97f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h60ec6e4eb8cd002797f6d27c3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1b16af1608ad4672adcb1aec5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5d3a753f42c83a8d90193a4be;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfe3abe231d5f200fe7dc927d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd66f90d84589c9f304836e28f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f5e0c08ceb6d08944793c12f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6349346f94a370fdfe2883371;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h16c69367331c37a1eaf839cea;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha4692c9375933a435a04870fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h510801d885b2afc82d1e341fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd7b268a2fbdfead641fb80386;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hda8b7ef10b7127e2fdcdf7785;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he2e1ea07b506a4c9fcf54f93b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h195ea0da8ede47fe2ac9df1fa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3d625a1e125d5e6c93d0c1210;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heb5cf47c9217d1c6c34d4d10c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h10facba025e83bf40285d13f9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h39eea6a79882c6f1fec2eaf56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcde9a3402f8fe505a20b03cb7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h440ed96e1750e1b950b9a4037;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3075233f5c6f7a205be244dbb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68ffd54b6a899a747cfe50304;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbbe7ada7a3f9d656a4b7a7505;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcba5387c87843dfc7b6a14f56;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha8d63b6ed23d7d844fc54fe9d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he8e858a26ec7a238b8443205;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5bd2f10c27789509dbf22b6c0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6588490053f33878fac42e86b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h56109f8b08734639f5996b4f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1bd6796de0d3c00d8d3d80da2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc36c87d537ba40bb848450937;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4f01cdf52913483424f139b4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he529c782ed1f874c1ed44ea09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7212de11a6982d59c06c63f8a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b5451b6fc994e4cd7755f9e7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8ed0f9db2a3aeb3d006847bc5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he48eaa2aac3080d125df7596d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfcd5e6f2d0a441ab28102f05a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfbb1611b8cfeaebde8bb40bd9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'heebb19c5ea04ee9106e9184c7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe312f0ddb5d3f7035572414b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1f4b282a741ffc7f2cd305bed;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa1809a53afe43724ba0c7f2d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h654bf7af62878eb2782808127;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h38edf430ab38a7342a46f796a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h730145e0dcfad10e31859c3bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7b652510a5f6fd9c0467b7639;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e182811e4e90fc41c184f322;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c35c63d91e7cd84ea2253f0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h90b01812ac4ba15059be376dd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8e2bde70b2fda9e45794ae964;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2820ab4984094878b6bf4ea70;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h37e3a6ace2d84fcb9b4b873d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbab54c180fba04e894e62efca;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcfa0bacf7f9048bd8b1f2a29e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9f999290dd4415b046c72317;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3407af4be48438d10d38e766a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h88c29245522f68b70ce29df73;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdf72314412eb0ff5bff99c0fb;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hc7325eacca58c6b4c94286f09;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he757f9a15885132ff4fb9b663;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8aaa2be160b3a2319881f800d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h33968229a2f5c332d2a315aa0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b2d9a51820a3ee27c6699b06;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbf128a1114a4bde524985042f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7f11821aab7cf75c998bbb85b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hef4a9a0c94b2cf08299f5ca0f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfa4b3c4a34aae856924ea83b9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fc6763b10980d0a6ce0cf84a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h123e699abeba1f58ec8513ef5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h34633c1ba9dfa542611a6394e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99994f6150fedf3cd3c2bfb2e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h73badddf33336272a53fb0528;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h655a8c6cb85688757f7f016b7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d151daab141ed55ea4d819c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9d21f16b79100cd4c2d8edd5b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ae15b9cc2275e5c06db9b4aa;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6943e18ea720221a13e4539f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hb52e96514c59def863cee1c7b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he205b03738debfaf6a57cc844;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31c416057465b827dc33427bc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7a23095b515b17cbd58cd7cc6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8c7966d36f2fd199b8710caf8;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h411720fe758b0e1b405a7b5f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h43932f30df401fb6df3d22c72;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8770f0dc67cac1917c324e6f1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4cfcfa5426b7399bfa5201438;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6b4724c3b72b340dfe26c9367;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h858dd00a44e48d86be773b289;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3462f52246edd316c8520acaf;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9288a6ef3452772d84d9560fd;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9693da9d47dea26716964a21;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd4ed536cfe79263c3b1f69f47;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4caa6b76db1e9426d8c58e9b1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h788e6d2e16f725fe329c31aa5;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h532d4c01c0a689cb144742fa3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h93e251de3b71cc0cfa521e119;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hcd801464d679e11be87dbb708;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h783d995079009d4b5c63bb9c1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd89a6b4408770364462f7147f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5fa62090905d11df1a4733d8e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5744260193c414aa120c842a0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h529c16784d04af4c49c3f500;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hbe992143c912519c9b6fbe8ee;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7fa334b768bf9242e4fd0499;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd572a5d9be5ce13f4e5ff0e4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7ef6ad4adf9cbe1bf627c14fc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3ae74952ee15f0c3152a23ffc;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h961bd96f3879f49f7f9b101e9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6962af5543e7e36eb47d3d1f6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'ha6bdf83a514814a28daed6da7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hab78886fb589065642e571f62;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h50c3ae0f0aa2394a5c8dd950;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hec94f84dd9c1e87a6748000a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he5041870aeffbf98af513bd43;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h1804a1715da3c6e91a4c415d6;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he6f282a9002edcceeb68a39c9;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h66931efecd4f6a9ee451fbc95;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h44078cde7779437a7a95c9d54;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h95d29f95650f1bbc62fcaad1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd40c9543aeb9bd1e22e40bae3;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h143e6bea8fd33283b49f9316;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h100d0740baab7fa453286a1f0;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'he360b9f9b2b6d682efaf70ded;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h3b884f44713b6d902414f1a4;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hd06226ea7376edd9e74a74f4d;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdff65ae1a548a3ab30c36886f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h7510d0ba224e3c4ca471890f7;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h5531ed581ed638a7375347152;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hfd79fd4b558d802ba0c2b0b94;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h68309b44b95a3514b68fa9095;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9a40c8f83ec09084a5741175c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h99e24900161451886160d3201;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b5d8eebda02ef707ee310538;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2a05054d4cbe66693c626d914;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h11d76e6dda324c7eaceb3a5c2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h31b6228c7f5d0934148078e0b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4d19c4b5249dc3db23e9f540f;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hccc5ccd5f4285d6c7a3a29343;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h198e9ddc8d86618d0a11b90a1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2b2f1ad6bd0631dcfb3f57bd2;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h2fbed52fec29593dc9e0bb95b;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'hdeb3dedafaaea70b5ce2b17c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h114047d82c42d1216d8e1fb53;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h26e55129534ce4b44b767762a;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h4240b0b1aca28f1aa6580fb83;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8b4f1400b1665093765df114c;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h936c0b5315310720f8382997e;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h6c7cfc79b3b9d87a7e44a6901;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h8fdac6726a0e947e012ffa8e1;
        #1
        {src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 100'h9c196a977816a74116ce6cb3e;
        #1
        $finish();
    end
endmodule
