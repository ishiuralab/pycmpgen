module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77f91ca4df308a4c89cd45d20038fa0ea1050438d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dccd539e343ec40ed9b704bb4864c552c06410fbab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2cc24a39e7ee9960949970340916859c701b9e61c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7196a792409a982db4a84daa40742940aff5ae48a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb804b80a7a90a5d06b9be24b3162c29c62dae05628;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6900dfa3a62a84261d285f6ef5827ed4154c80a160;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha03f9362d9f6b7402d34a3d7af38d369887e5e4584;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb9aff290f529b653f73618fbc16dd1e60640fc5b79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1c21b929e77676d582774bb7baf93f241477d6876;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h28455385fdf5f22c5cfd39a9ee6467142ff2e7bea1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd83fc43f4854e9d0e57c58cc124c05091060bcb62e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143fc6559abaa9aabfbeb0ba5b16281967eef7cda02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d8a5fce19a07efcfd0b5ddd7af0d4ab0cd914b52b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h176f4dd9222294ad27d54a4a01340416142740f096a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba7ed9b39542d419bf515ea79ee6e63977b3f98025;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1357ff4059c6524ac2dd0873007f3e500edffef4d5a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc510bff9a27f546192eeb6b8da8296c40a216064b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf68c535677bce2db56dc41543ab87b2057dfab52c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8908da4a80e0bf4d31caeb18af5265c927a34ba386;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184728c8a9d5db0829f9b8fc8f1d6f77db573bd8dfb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c55da2774222e43f617388c5b82823e1233fecb597;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2a009e6b7dd1ebf21fa2dad12e6947d79f4362e95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ce8c7d702badf2e6f54eaeb8bcb243640d874a136;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6ab7b3873a424ebd4437b5e688daed19df25e8eab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193150c24a48289df4e93342c8fc027389038acf36d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7eaec9db39019efd4263c5ce0988049359093f639;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h160328bc7dfedc6b54a4a7397ea2102968d56bbf354;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167055552ec8f362b611d1c28670b2218263d4cbbe5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13061773c42359978af5f9de0b49137ce467121456c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdfe745d89ffeb7c19a0c5f278177e01d9ad3ed571d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe5fbb9a4038511259dd8c02d8d461734fe6679e02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h26d0c743581ea6c343f0c536b75afc78e3be777c15;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97caf7f84f16bbec443eafa01df6f7ac18b0c35041;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d3e244e91cc40605d515cced3e2ed9dd26e4e72c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h83ec132b74a31c1b2b41785f5af90e1c22e82896b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcfa2c531bce1be8d9636ad22cf0ceb3cf889b408;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h950cdc8e35859267239b44682e72ebc03d0d2b3867;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0b6aa3d04fe1ebe1575f6b639ed53288eff2f81e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140e4776a1cbef07c93cfc1c7e80310c901d8218590;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10cb150a1a032b191a200a90e6adc11a298aed2673e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18938a16ddacee3336ab2eb8861d18d2ae747348450;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h25c50942dd01c04dce16ebad528324ae753464b6f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h733e3b722fc49d84ecda903aa78a403d400e9eee16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5408a2b6e7d80bbf2a90614257ac3c084b381d0bf8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4032078f292d2b973342980e34af0b710a47a1cd4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1781c9ca9b4f3a1cbc04a4df984052f24c7ed319f76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bef55853e0efedf61d1dac60dc4339dd4e51dcb28b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h189919bea0084294b392a1420db5a4443a2cfd3f729;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23b22d87e0f3a60596f2987803a16f61e8f27f187c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h41193f690b32089d11d62417cb94d32fe71af5f9bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h266dcc854484048e1e355e0f6f56db4d5fca25ce7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77e299d1c838b59de7ea904d300fecbd31a01f427;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc4ebc92959ea15fc1a71c358f9bbce54481580111;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134b160d993e3cb146e37a677953dc7b32bb56cf88e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a509200a46ac512ca21bdcbd6a8c6541a062efe741;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4292f3766950411b169d34ea929cc80660aee7a05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9fd5cd75d569d532ba76e1d732638c4e7a8e24a99b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6da60045d863396cd999f3e17d63ba906c096584df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11759b1b7b5c339b8116b09972d68d4d7e7e2d42fae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77c00cd36d4d3e7db5b19c1b035b739172413549ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161292096be1408b3fc107f6984ec08ef0ad948580d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a02869476b34f0879d172d3b6ee8f56556f596ef1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9c6f8c8dedf17fc211a26eab730b933e426c4bf2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb5b2d8638fbee21427a0b13dbf41fa6f3f013a0c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31773c3a214cd56464cda21dd70e5ddb422df8ccbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h199e79b3a106b8273f6f9209126f132c80a46619b89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ccb34d8d534f3ef9d3d10f56498040a9d2bbdf720;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137db9a24ca8ed0f95905503475f3c23e58577bca1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de984d481eaa5671c77b1556912d8ea285f5f2b2b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7df13bec27b6799ca9d50d2a1d16e8dcb86ffdf0d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131e3e4fa6a1581fb4f8ae9b2fce3f1ac9f965a1f68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hada6956eab93546b2435f7b17bc65548d2cddfa893;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a0a1b166efba4182e4d84df68773581819a4f730c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb84410f2d6c5cf11a427f9c8bfecd361ffe329273f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafc22b36f7d7ad882e1b78f718b5b3bb99030e0908;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169d4ec979621cde4abc42cfba18ab0b75c355a6a21;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57f67ec653ef3a7cd0fd828cba2c37c388b9d74ec8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h633d87a71f41ac78194d03539ea11e2308d0492fb5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc429851f7860d11b82bdb35c5b907c223decb1cf4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1c0626bbc17e84fa0e0fb038b4d3748d52c43e2f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb02fd2ecc92b458f54924e4f941293d5642707b61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9a815a75b462066afb1421e28e712565402bb4400;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8b6662ac66802b9769c8eced7e75253fd3fa967d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118110fac6915f5549044e1aa2e89b02443774bb885;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19076092546c3d719194fff7ee23b96854f346503ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a9b136f66fa938f36c77a9805f1dda17e3b596e27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1943124e492152d414b1c6a438f7330141a4bf47910;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dde68f0c1c77e3daef2548cb23a22239c24aa66d9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ffc5d7ce97a081fa3ecb430ac595ac6dcb9c82362;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d326d89a1013fd627d6ee432601d025953e4e3912;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24518365f4ecd3903c15109827afda792a7dbca296;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b399abe8d00c189f0e3cad71c0d3688408b6cac94;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1becddeafedd78a8fff4a0d4ff79615e1b3ec05c2a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1326a4ba2155113de657b6ef78711f27821c216cbb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b596bc268dd1a31e7abff64f7db3bac6ea7ed7a595;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131a9e56179d3ab4c6c29f7606cb1ac85e6532c1363;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145e60d2bafea0834e6eee6701fab08668a9c9476dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c762d6d7f7a00f86778d16c763de068169e71a427e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ee8c781c4e7d2df49f6f7a594971cb58e4240413a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13dfa042e4f7f7c0599d466842e2907868fe15134f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107e5a5a971526bf5a71b0423d0b549a6c7efafea52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1414c772e846a0a6988689cbaef5f7093418fd50393;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfde72800ffabec41766e47d79d272558cb2b988de4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6329ec3d288a49990fbd61337a3252826b783b77d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d93daec954cc657b824d009cd2876c17bb153005b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122c73c5e380715fff593eea726b1ce5dfdc00a193f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1860198355ece3af50af2ba5620f7ccfde8ebf39f61;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3fd7cc113285bb3419eab9548b3a3c3b9fe2d3de46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c562923c5375909eb7026ffc9b2021f0d2149d0a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc94f83c7cb231a729082fa90d1e03dbbe50eddecfb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbf335b66ec296779863e8620bb409a88b737822d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffec83bfdcd5c27a92045581b6133f6e5333fd1463;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bf6dc143a7e07c33a9f4f50451af505e6cb9eed10;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137290d91d8edca5aa50bc6bf23db2f8f6008342441;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182596ac80edf6afcfb2b206d0ce470992031a2c1ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1098a787685601ab4e9f3545aae38442317824d56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23a41f9469dc86ae73c3a6833b67dd5d5fb686c883;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158d2d078b00e5704ff480a3df9819e7a52cce0dc5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha119760962ac5cc902fbff1395bfc42183e880898b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8b3d11b85295cd442c903884b6e2a4ccf59c7c420;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd75765be684fe61dd10cc0a6d1ef0a460f40e0f6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1035a5459e5065a78f480bd01c5603acaaf999882eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8a57630bbfb70d824a84de5315f7f30b249e7ebd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1462f2bb0e434c927567d522065a0c8f7489388f7ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1099fb86d81b848dc7f86c9d3bfb87119b7658da63f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b5acc0e52ac09363d8f1a16cc6ac55c26fd948805;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1220bc34546c2366df512135a524dd3f9d7765ef820;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8a52c263291536e55dadf17cf41cae6cb6c572be2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21f539d74d1f7713ab0bd678292597b3aeab4e31f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7827287869c94d0a8f2876f7acf0d140de407f3d5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b8906f1e64e2d6217e1b48ef73d527b7af291cebb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h41387f6e0e63e09b71c9ea7bc0a19694d38542c652;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17cefae66ece331b045b341e3decf255ded366d5a16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3b082f1c8055350193060ea2867f27e17cad85ded;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ab174f4a8e44faa2f126c53986fe74425f44d2a92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11db31361e0d63f749179b0cc42e5c38a81ad9eb43f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h41ce66a8391acd428dd81ed90e7b9fdfd9adda64a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd03212c52cd0c92d57647e46e53b0aa75f29117a12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h154ca91d4b41be5aa5f9a851aeda2856a40abba6426;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf38c028c2c0f0a34120ccef8a5c5f1d7856f7f9752;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a7649b2a651f68c125b46e9f89c3d5b9d1ee38d3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122baaffd2fe81a7da3c11ac3dbcaccda2cc1cc7c7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd9ee9a29b732eb52c4f7233bcc8c0de66dc8fbb8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142f0550477e026c392e32c730682e3c4b787e0da44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3030e9053133fd126f0a7c538f5875b01094b6390c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101bd3457ae5f8306809c315830c04f2f868bc0a5d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a83d4448c6db955c1e0b1a5915865fe83baed52adf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9a52847633fc5345c98610a2a55c2bedc4ac98a91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147d378b22479de7a29aa852f7b86d18a4c009fc46b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he215758bcfed86ba3b9b0ea628bf9073c5346c5592;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b5221324cf5ef6419f8c6b4c6c168cdf1c6832a06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1835569c7492293d83e994711603c4a24927a9d3ab3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea17e03621d3bf688ba85b92822f0ecfb45881f280;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1567e010fbd26cb2e63c5cce7b6d3b6f1c498e9b8c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1987fd9de38d66d7ceaa93c3236196432928118943a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1c061c7b8b648faa3042e0e04b0c5554fa4b5a72f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e21bbc63dd37d9851c785aa9e92068354907cdbab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8cebfe1dc2d64df84381b40b493ead8a6d7810cd0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b639d78a7ce1970b966cac242688615c420912fb7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd26e5bb6d4ac2d6cf722859793cba14ae5bfa07d43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd755ed1407f04994c3ebe6100cbb552bd8f900823;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1705ae839893ee08715e53ac43e8dc4ba229d670ec9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea6209cbbe4d8fb63e82a14480cdc14182950073da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f56819dab43c769c2cc778140a0ee86411b58d214;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16596f5d9499ef78c36ac5b18cb730d2c98c655b85c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc6c2cd9a5267263b055cf842e63405365ba3a0cc0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd23eed0cbc59df45db0b84c356dcbdfa0c81b7c2e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1beed12d4cc3e5c6f0d9adaf14783648c0fc39f577a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1659ee422a123df45a03de8121af8a98ae34157a4e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h236b248bfcb56d1fafc7bc8bd21683d55299e8a813;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e9f83d3c76921e227103f31ad843c84780c8b8315;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6043a32d9dc47abea6931c5f5f2d1f01a05fd1d9da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ed5eddb334ee385ae5f7b9c47e0a3414b1838c410;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b7e11a049a1970a0418a193eb6efdc997cb5b5344;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf3fbedf654372a7db7956f7dedfb3a1742dd0738b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1701eb44014a47f7abe417c12f7ce451b66938dd12f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b0d20decadc0851725afb8376379755c749822c63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a120c96a3d8bc4c312a4fc753d255427ecd09c1d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9502d8c124e97eca7fb31fa7f7191db3ae6890eeb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19daa3e5895535821705b4c56652511c276b93adccb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df2708d5893acd1b01b92db8a78b231f7e0c0abad3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha44db272f28b5e83b2378173b0ef7ceb1b71d34884;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11398cdff23452e18c404864eec2f02fd5e5a3ce307;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c6c49b871c57a5a675d0e9b9d7ee869a4cbfc4dee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ed19751abe6bedc3a4523f2278e9174401edcf065;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b062918839a21f915636500dfa1855ca45ae593f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9cef73ba967dc580ef715fd1690d53fc7e9b20f1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c8e14189620679532636bcd6cf9e100d4253e82ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12a6bbde9ad66eaf92528c5b9bb6448e0fd6dd152e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae1d60d0fa27b28de57a6c35243641ba1691432c8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae0b6d29b12113d71fea91982a1664dc35b533cbfd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he50dc3a3d39efc4e11e80f025865f6400440ccabfb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d9a7070ba97821a46ddf09dbb49cb38c8badd77c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3dfb93283583367d4d8e14b2280274896b617c2452;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93e470c7f4b6d03d21c30fe9e5a035023a9b19f639;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d11b4ed2f189627ec7398705927245299d510968d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13822dab3436178bed5428b42d472ed30d1542434fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae1f9c6cc64ad493f71e571cbe571aa97115de04a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19632fb2359a9882f53877de0486be802f7fff7c2da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d46b221944d2b6794f861e0353a6c834d85135353;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc76a7be97dfef234711a6bd4221658410afce8c1e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e34ae8370c8a6abb8186cdf27734403b9dfe0837d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9b680596359b50fd99094a6886cbff3bec9a46c4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc8fade6e509a7f4779db6c520a4e7ac1131acbab0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6edfd526f0b1a4de5f789753a1ff12674edc3e16f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ea0b00722c19d46adca6b34c2a75360dc8a455f49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61edf501bc824ff9c4e34860c0382ea57b7d8f8a62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19cd9bf7d25dc00a47c751cf626aba9d223468d7e4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12fa5f7522b4bd9c3592fb865b350318eabadd8de2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f490e8acbc6f67c33187f37358e37ff207c556a3b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h543de4f0f577552d3f7cc207a83b39633a5f0498c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b5c9ef0db8d13b343a19447a0c1ec692ab82f97f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90c8090e5b6ed3f11db592d2b5eb67ff241190fb43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa5a44dc3d92b8ef160e28003ac9aa254349545075;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb44e90c46d86b0b2c5db2eb36fa6a761ded22b8dc5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda907050e21ec708f400908c7ac7f3c9d44b3381d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75e79fabefd4a7c1793be30ad65712be09b344cb41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce6550afa2c9a453c2c0e145a63f0951cec37f37a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf02c43eac268cc406e78d114386e993c7df5b9da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfce81bfa0f87c4d4881a01c8ba931bd16689a49cc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2b34ada7b1fa738ae915505359e175bedeb1c152d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1532ffec99533c106146254ae779c297af8e9f50c36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha396b501ff5f4c8434d0b6365b9ba725c8ad2c07ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe62173a1afc39a1ef6063923f6fae6387ab3e9bba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c8bd92e181e9e9118bd2de09b64146d4f589c84ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177db94d827f70d809e21859d88fd72eda4bf83c18b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba00410c3e8a91366e50c1f1464f3e54c637741ec1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1256068714dfeb6465aae80f10dcaae683a9bfeb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h369b865e89552bb7f169be1cdf733de3062a10c5c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1225e1927d0a13502e0b7aabf3a4e753424b72c1543;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cd145f3703ae949c303d6f164a542e17860325ae9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb273b1397d95a4560b30cf9a6752ae9f78accc2f92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7a64a4babdc394669fbc0e25f204d6956e67f2e6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165347453903d29375a6b4355203024af0955e95233;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10eb8b2fad305768871bea25a98273eab549cc99c1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h574760a82c79cb5fffa63b2f453b536aca5cb2a611;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1236d8fb6a9aa793ebcc1577a9c83c7c0d95f72dc06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa111fa8fc41d8ee9df1256966dea6098ae0e58b2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90ffb8aaf41c1e88e784f16d67902d8230504b0b65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha14acc3a8851aca5614f9a8cb82ab6670544e0fe3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56e89cd39aef50509f67feb3dd586619be58566ed0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55913655212c452c1233b2280686e77bd02adeb3d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52bebd46e99f27ad190d46eebdb8b2a55766a0175b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf10c884dd9a9ada4ce94afc95988c1b4ebe16bc2f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bb0942bc624ba0653309b40ebfd0d3be2b10eaf5f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1275b209af1614059a662564321da6d63aeb3e0c117;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df6d9cb72d0f6e84af498a6e22b3bc8bd892a3ecfc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e57dc31c0ee93ed4740ab848ae08bb7d978874fe0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1adece9fd93d27ea15c79de5c910dbc7b45966c5f15;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8167721de207d9b4e64d228f7b2e41ec03156c1f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca241410c4f2dfdc623e8c0a004cd75f4807178625;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f07088cd6f5857c9b01dc84bc29911eeedef9bcd82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5b86de3485d93698c2822649fc9486c3fd7b00088;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h151852cf892dbee81ac9c59f8d044343e871f5d5f42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110cfaea2221a12fb1b4c1cef0eb824af2ff7b90f93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183ea362033825180dc9d65ed5d90364cbf113ce0a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb5323998eeba440273ee87846225252d5b8c8abb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb061f0380c3de29a46e51d96483ab13e73f332e0c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9c0f5b99d1a05fd8ae851ded7a95dd7f638605643;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d28d7baa7d3931b115fe9b7bdf3032b8aad9df1c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ada5a92a28b683ae00949c19036036952900b5ec8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c43e4bd7023560082d4819094053693e305e755bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h224af40955c22b2c857438a2b496ff70136781acb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h874af7de2f8f05fa0d0f89880f9e164a3b6e1c94d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he12cbbb21e203185dc87204a6641cb42cf93850200;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3801b414a9a974be748469f33c99810f7251ff0f30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha140ec3db066f170776cd0f2badd518582b24299b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1247ae6bbbe0c7e523d9ad1d05c28df837ac249f90a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4aa0cec81bffaff3af9cca15c347366e708cf6657;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad67638d9a053d634bb3faf86191862ffb30314f89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h88caec81a1aea8e57846b4e0ff5db89eaa214d19b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f2216490c763458dc9ff18e838eeac5223216085f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d34a3e4862518e4015f9a6a9fd0755b009379c748;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10be0f0526304cc87bcad7a2be043efc22d33bb4c3a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2b44c2a9a64af06f440dee97b27c418f953b4063b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c10cdf7d6ab32f6ca1967cbdf714b4ee95b4cdfd0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12aa433505a58024ce942169d709f7fb666697023f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e365fbae17fe3222a7be9d58327a96fb43d799af84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17108002e6ba634644be5205b8ed60f47bc97bcd213;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f0704410dc792c8379e9e395b74825fb7ea4085470;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b378ab83ce0648c3de92f6d1a5b93cf70a328fe1d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7af78d15a58106228f5ec3d4aaf1f0193ab05957d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19511c0f47258193d4f160293ddf0386794ec473a56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea87d6608342fce39db5aba3c58bd157911bd04199;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd4993fe00d700beff283839f6b95eda9572a0135a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10247e60c6216c3e9cd63a68469af889db9bd3032cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f5212aaef6303ff2c8fd7317c62e004e37b2ed50e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166cc7e69393338b99e099be61683115652aac69a6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1d88b4ea04e833da2a7b1e1134686a221078e08c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf7b0f179a14d2e76c0b27acda45b36006de46edc1c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198a4e1de19c4b67451c191380045bb4536b1dce713;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ab49a693ab4ebc72760191fdcf76b0bf0dd357891;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18dabae80998dcff22be70848f501ac83372e81d070;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1302f4497ed13d9f50409526d02089f98a9089d94a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171c1e701fd228e5c22be04aed129779f7d54106df4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3947a03a8f6283856af6e8e4c0f4da69b8457cb013;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171ab21b2cf00f5cdc1aa398429d5ec2faf9f8a3b74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c394f3c4aacda7cecaaec753ead1628ddc324f6900;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac20c942b37a7612daf60b7a49891ad4b07d38e4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192aa83f483978e3250453bbfabd48c167c5d2afa38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eb132c0d742cd7aa1f554430828ce83ebbabdf8135;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29b17b8b27e4b9508ca16fa181e3569b911b51a6a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he839b5db6a3a2623c4a9bcf131574519403d72c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3165458894354bb91f96b32114d49c76829663da4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc45a594933c8340499df19545d5719c71865cf206;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c204d59070ab1aebcb70cffd030c3cb081cd40de8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc01ac4a0c788b8676151059f93d3d9ff6635301f52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcf779cea96e92615d59a7b654c31230b643ec7eb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf472e4916633b0dd7869189a71de3f39911a7338ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12fb507b00bfc626d8081002effccdb5e7f1fb68459;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc86f181007b330bdf50740fa963c4ebd1e54a943dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c727335dadeba391ac1f8d7f47b259414540af6a50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h247559cb8204295b2405204c5e75785029a9e12372;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h196e63c39cb332e3a242cd91f67e047f8d3f2f3d3ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce031a0a394457451366de1eaba1f0b8fbd505e18b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc50d7a616171d324fe7b2866618233b3db98be8dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef3d02d2d9269f609cd25e161c945c7cf252115e49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73bcccf026db05f2969679d06ca804e5c29387c3ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cdc4e8dad292347b8fc44fea37286d952377fed83b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9cac976ba8f3b8dd9126d07871a16f5dfcfa11e87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1434c2c8a3cb0084cb6f26710923a2567c513124ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf37e3bad4f48e4cbfb7431652fc22d560a44a39da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd12da6ce0e9989e8dfce39ccf47554df53916bd76b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1129e82d6fc8c4ddc9df494d3e94da2390d0dd69154;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3887a975815e16d36f73649c74f2b9f53c3fed6c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1153097a6ecec874267bf13562ad7f4a3d63c8254d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a7a2ac1897944b83395bb36f0a930023ed8394603;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3befe2ea6efb58a506d942a8c8a036c440f9b5c2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9047c4facb55536bc5f63526aae53f82245f6850e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2bfcc923c77f15113a75001ad3033038275009887;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e26226d0a3f5575ababbabf821d086a180af7ca2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184db0de55c12eaa51e522120f20e39fc8104430c41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1ba58481fb64babaca2cc9733f722009ac35eebca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40982d4678c674492e989b41d5b2f0235a05b7c365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h484ad457cb2d805a51dbc39e4ab61964db3cdbf408;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h590ffa564437bdc276eebbbb53645ab15c56df724e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heea4893cbb16295f5049d7f4e2739863c333e7e0d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2ff56dd82d4f98f52ce0005046d8a65a443eda6ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172ceb64a85066013b4d5a94fcf0be03164a1b6e5b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1444f2eb7baa00ce778e9846bcbd63e00935f1fc37d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6c534fbb3c1fccbfdf8227054d506e81f5bf33e86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c2bb68d6c924c0f7ee09a0b72165b12e21a6e007a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he20ada689fd7d48927016222014e6d2268ce0d5a7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c6b18866c4713b8243b0275a53d8f7c7a8e73917f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1068510135c1b49bb56c03647ac398f48d6ff8c2f8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7af5710a82fb3c40d27e42745ac0cc01569430bc27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e86ad8ca212ca620cf551a7629dbfbd263c93ed7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafd7687d103565da2e768da5791c7d161d2c159e59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h76fdaa74a692d6afb6536308271689dd50dc6d5145;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16bc960866b32ea4c163d61d21dbacf90ba715761d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7be0a0cc42e0fb9531ec5b4e416f9dda9dd9c3765;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h433d185f1e39bd6ca53c758cec2f30c14241a0b822;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a22e9a7e2ba12d781355be39bc1e0f9087c0dbb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9e4f0579788e884041b7632fb97583a23e42ebd76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc675f3dfdc211beef93abf81e1f0b503c11ed2fdf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc8c955284bce39b6f7647195d27dca7c39849156;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174d44ca3d814f725376f6c20d533757560bb730779;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ed2203ba76855069ee8c2ba121c3c4daf10a1840b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h789125e8ab5b0d63f0221d9ee691474e0e2c7db3db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2a12e25d8316c073a74cdc4f231b907d82f677aed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1444dc5aff132c1733f76f31d09598239a932dad28a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bbb35c284ca25d882e83fa50b13dcb6683aa94b29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ca729a249c826357e69e8f5ad9b4c41067b43fc22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b0b9a7e6bcb57bb468f906ce99d4c6bd079e3ba70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124a4e650acdd436af21d0ba527a2c2971748a250fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h326a1a4d1399626c7019377aafa4c83b6dd21a69ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17be71b2d42c98cf2eb0dd83747f0e4ccb37a166425;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd6cf033f1d164e14a1bc7a9637409354d27d6032c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18621ce024e7200231d153772b03c34ecf968606ff5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa319e6703d3aae8f70070d186a9a4845e40f08f2f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af4a51919273ea82b5e2a0d206ed4b03e63d5e2b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1adc23220a50b99d071a726b594d3ceb8e3f17f1792;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1673bf5c95722d8c210716c537f6c4ebc0cec580641;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e19c0e70d172965708960daf84dec5ffb4583a350d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a48550f6bb6b1622676c533e48fe59af794d9ad1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e6ff23d9e601f972361d161cbf3174fb620a9b373;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1efddeab0b6ba4a70de439cf98864aa74d6ee0f0aa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc34f5f2e0589722d5f656aef15316aadad30cdf56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2428e47e7640c3a4f18ef3ae68c3306e5811c9ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9afcdc8a9a0e486c54baaabe09ee3a4a7d5d6568a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eb9fb62544f806a08001c1d92d14678167fc566180;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6442224f90da10a7c05712f4b24767a455176b2de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h391f671737181ab7b121053a2f670b1e8d5dbc4d8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6fa056a2baf5a3a24905658e19807bba2d500ac24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a594b07272fd8704d449e9b57b0e5b4b9cfee8d6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15329c10a366bc022c4194db7af10f9cdedd83ae982;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e9b7440f29d45cb21c45f155c96d4b8c118fc7aab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15500247aeaca65066c5d6c720411a2df9ec087d8cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12117b6bcb116e9a3f519d15283dcf88c77ce77d51d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea73bbb37039b18a20924f3669515cb192ed95556a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a76d3e43ec37e268e4f40c0dc6bac80ada261df737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1274f69b59dc3850721c9bcb93f257bbf562fdba499;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6396a426e87b5e07ff33570966fc30c05f9de7a6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4aea5d337213eaa3d2672d5b4a021bfd4ed802f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf91aa5ae05de86be269cd2d2ee8c744a4e298fe6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h615ab5738bb758857754601055f709def17548c2bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108d56853b848065001edb366baa7715cc29017b3e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6b74cad74f44ac74fa3884129d9d391e1ba9c9647;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138be72429bb7ad3cb894f3109cc48146820a3949c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a23ec5da5ee7f33181f2862f47e9ce1619e853c3ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a446c9a2645d24b6642596430d9c27e799e7be02cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14179fa68656f1adad49f1f9cc291aa4df866762838;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c95121f3c9b9391da7721a972386672906d60b356;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17fdf8399a713e683786e3365b32eabf61a49d69865;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18580ad4501a5ab4f5dd0c68cd0ae09534719492b10;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c58efd4293b07e86231c126c6251c67b18f08fd90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df9cd2b76d6f7fe54a46ebfa832a00e023e4a6f655;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc44f9649342d9c5fb4e5e4bb7ef3705c1696a94e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d388296d0bb2980abbaf6ba9e9225187efa9362b04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11fbf0350d35908d51fc3293929164be3c5ec6adb57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1239e55d0fbe345ea55bb52ca2c99a2f2f2113069;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hacaa11d2f105b419880afcca49ce3927eba9e34953;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12a16396723a35b5056a29b3c5cacfbaaf632855f55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10bf9db33ebafe6adab99bf406354a503d50f337202;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15c9dfb8b45e384e395198e6f48b549dda98068dfb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1abcf94593f9d1a9fa8e190913903e66c6f55f3e22f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6dfaed1278e6bea93e747e42d67ce03a6843ed698f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7d44593ee051eed403337a60b017497261af33368;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140700a44fe30fb9d384a0820eb5f2c5c8b058e5285;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe2b651f4c7054429c1b3d220d2250d26508696b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8912b1278f596ac16b14608af3afc4585886dbeda1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa659aa93f0d4014ec2894c6ea5f4f65a1720e9be8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0615983d482f117b37c9e150f6fed4a2398550aeb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4443c8401e743db884a08fc2bda5b38bb9773bc4d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13777f1b301df8dc86e26be653d4323ac2b7ae930bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d8d88913fd4904377e687d9d9072a17029911d87a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e3d2bcf66dbe25a3bc1fea8b080c9c96444bec60e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1737a0950bb99c5344d1dd2fd4bdcb75a0c8ac01e01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e65593b8a9982ea476eff24dffc4cd34fdc967c97b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12212c2b43de24a61edeae76c0d6e947e4fa2f9e54f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14981e69f9997ed73a127e01225fcae064201fbcbed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17c167e04546e9751dd8df36602db9d568cc9844eb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5af9ab6855391e8928b1fa6299aaa375f9c3fa415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd69a787078f6eeb23e7d36d01f638f763e46e150b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha34cf89747766e29a4ccfaa13a57c994d365649d81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1f53d7e4aa8115f5ddb347165594303d13bdc90ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1840fff92c2b297d66459e3db90d4b90fe1908d7e2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h34714dd653b348c5d9003b8413dacb846cfde75317;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd27814d7367dede21a419cb0880119d844be72fb4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113342dc88dfba7e67ed69b42525995fc115ad4f6bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f362755372354226e39a7581777c491588491e8e06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1d881e848d41b264b2281f07854952ad34221dba3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf3c77edd10744232b9668d905d7ab48daa1445927;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a7ab1e0619e160f7b629267010e3ac7c9d8daca4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b18647cb9bf3905c60f417d0921a08bc25c581aab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcabcb2ab9aa464301298c60218272c7a76b85e793e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1971adef2ef14f7da0380be5162a0f7e0e4abed0fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1267fdd4487edce12ce46ba0408a48cfa3455210197;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h618a7e5e340786625c4132cb2cd1eb30ffa828f15b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h236c934d80c1587a23d185157403b301cef66ce825;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1772f1ef5ac9ea513dbedc12d534c72dca0cdafc138;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53f7db364327ff16961d84d237adde5d49ea152d68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf803e1dc80b5dfbb188d0e46dac303f9e212a50a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13da097508a268bad1bb215ba1beeb0ffdcddddbfd3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ba532074387adb69bca35d1cb056765655ac23d35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f51364ab25cd7eade07b14163035533a6a6ab28d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h702416b8838d43134581c782e8e8dafa1b766bd72f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ca62c06796f08e231afb62d1d2e9cc6da55f8c787;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h513667fac111594b80ed292b8e25edc2f224c0844a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3e5b1a798362e131a9a08f6df16811c6a09f572597;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1b0c4370cfc0c2fc39323630cbb831f41ace66963;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ced44e5f0e2457514e50af2bb167503e0341ae0b49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6fb44a5a87ece1a92ff2ded2104e8f09a5b55efc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4c60329b525e127a0edab15b5de2b8d5bf3a78268;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d864eecc73125992f7cf39e6d587523c8ee6bc58a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h178fd30efb4fa9d7b6b8002f9703d68a7c170b609ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5376bd0ad0671a5ea176b0b1f70ee7dad124d3f45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198f542427b92246872d23f5a3b95abe9954826a596;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf50eb48d1cc9a2d4c765bcc470cc0fe02c6ce0885;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97b0982d0b4a5bddbb957e353a9f118df8ccf7e4a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14dccd05f551c3940d4175313eb8906f76968a0bbe3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1433ef0420dc70ae0f96c4a3ab697a1362973dc907a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1066b66da751cfa2e31c313d60859757ceda458c534;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8de31c4c694346a7e7f39eab8eb684b274dc9e056;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h440e8607bf8ad3c3ccfbca3472e47f7e25422d5e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c1b48b14a0d4d54a9952926feeaece416a7463840;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158a21ff1fa08f65682ec4bce7e50a1e4f232a7e894;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d79feaeb9e0e59d421aab44747b3e49d422ddc7eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbefd09beb1caf80f23827bc352abed774367d869d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h607470fc24fdc2842172f830182e25593c52ef554c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d7e3bbe97fd588cdccb7ffe8f1fe2987db4e22e9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f9a6e24a662784d0a2ed7220cd5b9c6683e71fabb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa616c4d3a81e67e19d0d6af8452d3a1f5c0cfba93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h274c2111914a24a3cd185922ec586e895ff993643e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd03cd035e9a03ee78b5b8db417ad91c3c1be013971;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6b94b93b3b86067fbcd89230da8f757ddbdbb3157;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9d99bc5436dcbfc62de06444909fd3d132553d8a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eaaf092beae9a318ffeb701369be10631e971c7025;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac713c50a8c9fe29c257b44cd71e0e6ace67837eef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ba3126862b24ca5f21568838c686c3e2327be3028;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63fed354e4369c484fe141bad2d8cd5e2038c8243b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4a9f8ad950c42f5220a6da56133d384f1892363b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e1acc07be0c350067d88d6502c064261f3f8105a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffd31b0dea5a83b3ab23fc0daba72a87a4df73d595;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1285a4c38c3427c46ed965eea46776263d017ca4353;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd8a6dff95a6f86f794ffd7da6a230bd3e5285e186;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e6e728e466bc66c56f443fab65834729135fe1d7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165e3bb352a27739d43843baacfe813b76212894102;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d941b4ac3d679b6b042e65ac18c7d6a3c0a519d4d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b2a148559f4cfb4334f2ec5c811e7e6fee6e1b3d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ad6eaa811d4a5f6565d57421df3359602c8634227;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c9166fc6c684307b3fb83924823c14c20415552d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2efaaa42575ae7ea295a8bdc2c9f8cbcf5f236d2b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125cc0a334ec84c777f023a3773bee1a89374475dc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b3753ad264a0915c83d4b48161b240b2d525bcbd7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a68fdae4af32b3ac1bc7e35b4f90c9d1aa956a367f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68870fd16ab670b988fc972666b0418a8a74dd97a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc44d4e529a278eff119bf85f8f1312e9956d255081;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf0b98cae3fc51ebc6b03879eef6015e180803d55c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137866dce5692efef549a25ca30ef495d0ce2041c8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12dd144e3f250861de02e0d251a5e47adc01a80301e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ab83fdf682af376e88ca913c857502c6b643490de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h793f5e41ba929caad5558881e7cfd26cb8c0402a54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h25bb4949b25417e46b839ec9aaf2ef43b80e9d0c96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc4d79a3eff04c1cce0ac40a4438f5dda1a4a04b8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4bfe0e33ee362daf9b12cb82a5dd1c2c804d3a5b0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h186c22a2b8436d72fbfe3a9cfa7ce0a906b9149741;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3cc7337a1b960ee3ae5fe9e700badf91762bc8eee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0b1f594d1911cf6564e72766828f7e2fd7d4c55f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1532e6339efd3aa61a9a3dd57048bf11e477c09f1fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b26368041cb2ad8faece2309ae855030d6885f488;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fee6f870e730603790480216db3b15d1218a725e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9381ecb5c45eff9a4800d4692f46fe1cc9cd44218e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha851f141858b1d41b0413035037c40f74addd36786;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e7c8fa38084be0b0573417522635f832a0f85b425;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ba86beb51d61b98272d0f1853aa2e108716a2fc5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38fb10230fc6a4ea61720bf27038906a69e4a85fa7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b914d2b1d50dc15621265d9f7182a3811cf8284ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8fed164a760e106907f132c3ec98b87a3b5ee9fb07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4bf3e1bdd6a71f9b86ccfb6a25ace0e5eb2a0f7f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150f67eac24a4e035a5daf58fffdf6da2c61403f0ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a185d97f238a75c0f1122cfc4708ce4583267b683f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1553b51d4d94349e6c282a8eecb6f609b8a2961c24f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h498e3e0bc53052bc164270718ad30ec86a2a68d2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146f9c38860ef3cfe2e17d34f45bceebcd321a74333;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155b4fc1e159d2791956bb5ff84544260a9c6113a2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13307c29329ef6d3eabf3292e99a0d2a679c784b991;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13173b2255d8044fc8b02a89d5357c1d4754b6c6a2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81127559c4b2039ae17992593f8138cb39a16dac99;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb925cdb2f8726e4a58d9ee0216339f3567b8715814;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138e85fdae93145dbaa5a48834ef7240beab3d9f8f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h778cb206c232264c53ed04218b08aea4d9a9646344;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6bf4d52e06ef6e3deb2309d3ad811a968847e88f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d1bee300ccd824e7b7b84ecfe04f3f2cc886fd4ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e274a35d4c17d90d4143e01a4a8b37754a2001a9fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38c2aee7a51b09ad10cc7a59338c34c044de5ef8e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d58db4f001f97a5fe27f6704c463874281d35a56d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171dfe17c951d2fc02669e8c6abb543794d24dee9f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h139a91e7c4c7b582376d819b3d31a854547b39f3736;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haffd5e6ba4528ad6c9860eb6a31fc19c3fc7930fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b0b17ffe23a0a59a5fe1fb9bad06c5058065fff50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h609bb0561d3c46ede482e79a9dbc389ddc5b6b4a04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4221e8c081a7d9b293295d99247f43026d306b5315;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb59c28cb212f22760181f585f121d8047b09193a56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4b971053dda428fec1ba587c94c6497329bdf77ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d5e6b64aaac55646638dd42a4669ca7d564c6f5d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14195485f61602c2eff490537748c03ca8a98c9d992;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1453db03ac4e8b8eeed46318fbad44d3ba15d72419d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f0ef9107869e2b6405f4d3617f75c203e5b30441cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169181fb5f68ec8b8cbbedcfa40b66b5cd394911418;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4edd851886e570a229446fdfaa1dbf1f1d2899d8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c429555e5903880ea28ad16b631d654b107cad640a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7fae2ffd0d590aa536ccdc8f63efca66769754816;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7821751e8b446b86036155969188e18f40c0a4ea5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac7ee8b4d8a5ca3d2c4737b250ed5b445c8ef02524;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e5bb0151ab2fa0ac31ef0aca6000cee0d4ece955;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c26eab4b25cffebab27d6f8104714d7ebe146ff6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd5e5f48455a079cb6cddaca1cfbb057777d9fe87f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1291ed3d637c949d46b97124ceac1f01bc559868ab7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ff9d8a25bc298fd592c3b307067af936c4beef56e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12da82360c005c1e780705f74f5ef8eaee2ebb80c83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d4c0d1ab481239634877df1ee0dfb94b505098db1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8caaedbba309ab4a0f604977d3b094a3115796996;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf223d26534dc8e2aaf25c61ca671ebe09ad4255397;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dae5740045340846fba74bb757ab9825582c543235;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafd6621b93d0cf9435291898224212af7d8b131391;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17493e1fc9e564bdac6384fc16a2c19768a569205db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5201c4c23717650425b8ba45f6c2f3201a3f5337ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h191caff1029903a3997379f502bebeb9ad888df4a1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c10e60d1067fb235fbca0c6b75e3d264ae31f6946;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a55f03a63b20f0ca8ca09a7fcd1a9cc852e6dc00d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f99d4ff9abfd9364b8701ab5bb8b8463b43a3abc26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h949912716db4312096cb4c025cb5120749e9cc9daa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc75bd159f1e77bc5710d36e3fc018b2e8902b9b0d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had082eb6038ed6d0106f8929adf562588a87b25027;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h358e9f3ab0fcb392372cd0c9d5fbe76a5e9f21f9b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fedc420bfebcbcf92ac03277e63e606a747f193448;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85ec24bb1c4938383cd127c0df5224a0c4f20048c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182de939d3d6dc542aa561d7367a55e6ccbf3536f09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd142719bbea477b252da8bc4c580a4da1fec05a40f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h103512108053ab3f6bcdac156cd47c5598b33ee48f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17116be1b6b52a170b271fec7e3c3f9ebf658f636f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d0440ae302fd8d934ed265e83f25646c50a29fd1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c291698ef8652847253f87c8d71ebe979966e05513;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffbe9766ecf9130145bd422983de447e5fefbd6ff1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5bb793104705aadc9940db24d34182c4c9f536ca91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14dd12f2c59720c06d6ea30dd52891775307a65e26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11733d8f8ee7197546c61cf1b0928736479edf27d8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha04550ea629ad082a96a58bf87592dabb88aedd1c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d7e772d6ff088dfd688aee059ef299640ca4f6bf2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9854494e94ced8ab25183251551eea9da9ed25ebb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db967dc09b86f6e2b859aa0bc190f470ec86407dcf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5e0c6d7630a98597376c9002ad9f2f544b2a241e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e806ca4691b009fdabb1de1fd6f59678f079e5d00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2bbb523c4652aafcd2dda6a0e56f269f4fb1fe1cbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ff34d0f513009b27e1fcd8362c41fd8ffcc3e0e4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h79b3e019d3a4b56f97abda99e6e2d4a22cdea7960c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb3c0d93581248158196bd33535899edabf832413b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef581efb65e12a93f729ef4b64071f7d3a91164348;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd327fe033baa1aff008663782b6d23e41857df1b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10958cc69d68f277962b779081f4266010c98e70e56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h33b6402ea22f4032ce20b58715a2a22101e680263e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he83c912faabf4f8420e08cad5c5693454a4d1b7f80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f9d4677a46ac54f3c8a50722622dc9419ce90ee67c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171e5549d6d9e64fcae1f95907e5d516aba9a924e0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c79f399d6bad9f8920070c5a6c1a4252f773cd74ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116d7d03eb336050933c7752bbdcf2e099817bc9b23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a784a34b9bb154775cbd26af30f254de7e59991591;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14146e9aee80b6a01936a48aaa34ef094fae62f7fb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3ea8de07494a18aa9d406f295d587fc0887b3f0282;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f523f0728463fb627d49efb5e78b2d19ec5d51415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h20d06c4c0cd1f48b7845046ac7e1b47ba2a40f001d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb22ad6d2c981d58d2c2138735a5677a6e635e09ba1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had38df3884ecb7f06e283dfdf3266ab51562913537;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h353bdfb216868b53356ccffd046070b5614083cb3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f6b87f4fb0154f3095704a7838feea9d31f870a74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h711ee7f28f0e7a8add28bf59d3220b533635268e15;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe917ec556c06c531a9f04c0dccc3aa345cff31a65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f598ed5849103f78f1733e3fdc4bedff1641eea97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a37fd7e83dc1b0aa49df571da9bd28650ad2e67f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11bb2685ea80c9ae34c94b2247027b1392d390745bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hccd15e37936bf3603ac10bc988afcc2480bba675f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf284b807043f76802cf09bda7641e9e98c5489016;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h100db02ae6ceff326fcf12c571eaa4be02b641fc60a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf9568a6c62e7b359e0740cb410292a3f299c2f7ceb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h775e18d7bacc7008bbad481a040ed08706eef0341f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130d07495bcd085d6086332167e552a80e7b9f91046;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff225629ac9ea4ce62ff143fbd59d05c26e236d42b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2b08816d19fdaaf626d9f5e82f894468ff9ff493b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b400a5b79e194907f6c813f765a7cdad2b18657b32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b8006aec9aa1b9fcc29839e75ea37c466945704a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123c1b204a98368fe93d7bb40599d25908a922f1753;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5945f4eeddb98778461cebbe20d4046f6b76ceb36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h154ff7eeefd2f769e5ff513b71263abf25fc3cc3719;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h798946b2789a4f7339922ce451da207cc6f2ede71c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6855d4f19d7fca0356b0bc4078e66a05e423ffc921;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h736ba049185ee45772565f57d896fa7ae8323fffee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f840408bdcd3a2d1dd2638e0177b5607ca7d06a11b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a31c4d76e5f6fb1fe0623940e268a4f9f3ef7bfb76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad3aeba97182b21d0a1df7cb3634e429746e02b977;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6fb1ce5c29149b1a08853030a67e500b01daba9dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1968e6a460c2dc3cba7e48970a8fe98d4766b180b34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e674a33e75d94106ac143c60ca7f96fa3dceaf9552;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb7be1d90b7043b134b4a8b2e69ede4c44c1fc8532;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11899b1b8a8f06e7e55ae890768c6e9ad5d3ca4d8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf3cdb46dde7df02fbf9ae4d11900585fb6e90d4da2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ee7934077a97efd31a4c12f7a7f8f57df47065ae0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1899295cacff25f57ee2131b7af9dfc1e5d23f5d774;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14cf08f4d0b59ab87d046d084d36e2223f27365de04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5afec17f8f1a918264be7a1fe624b774ec541ee910;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf3677cd21e6355537f1e323aa2baafcf8f33756d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4bad6f7c9596a07aa74116d620bd3bae1ea123c05c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db6397eb0e7cf2f4ab5e3d3d27eea18a6137b07318;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b61c6a9d6ad22ace05ed2264b5ddac30a17ad6afb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ffeaef267c08d02d76560cd29c3ba17461dbe05e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa17db0da9a1c32d48fd625756bdecc53a250aa88c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190b77a4e755564d8dd25dcc04923c66e075cac2814;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e224c9be3b0f6552d7075c3bf2f925057c237703d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a52827780d71d8960d0594455a026707e31d61057a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3de84d23ffae181269d8219037598345c3ebce793;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1c6e4b16c35f5383fa2121893d55460f3e8fbfdab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h28f3816c0955d9fa9c5d5b614c7d697428cdbe6337;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168f02471d027267f193dce5403926091a55cb4bd49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h48708a5514ea0bb890414cc60b9b21eb9becfe9ff6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16102d5337cee97a784c5abea016550e40db62c39b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d5464f842dc87b5566da85006eb84ca141ed7cb84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a063583419d8995a7b52b988af3f0ce68ede045dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f2e70fe320b5f8124a23ed3865444f1bd02a06ebf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a72cce5a7424b69841654fa851e8082662e503f18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156ec614e2fe8a38baaab7631c2e4f78b2c72654ff6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h99b1485fa64456d86f772291c1231d2d3e3c1ce8cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1447aeba8e8aa0cc18b9a85edb2cd8aaeb2d1ef5ec7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a9ed340223c9c2587d6793fdf47b0f777a494e38c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167604ca5470dbb70ce6343097555a19f64aa6af909;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd330e67180b7b303c6c0aedf7907afcf24f5547e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb37f4aaa64e5e896cfc3d41b31af239185c0ad315e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ff91c16ae6796992d3e9a7eb8151b7bcf362bcdac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h212156f84f7add37550005bfbdd30276153270b220;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146da01a66b8c0bef37dbbdb2abb06a2c44198ee4fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18491fe766a22256bdcbf5b398464d9a39d8cda986;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187d4184c1cad1f05bbf2090a38b8505ba44a05ace2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d17e9d0cd6633dee6789f0548028a8b91f25a1146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1241317e6717f1ea61a5b81df720a599ba0dcfb13a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b75f7864d60ab68907e17dbcd733590f96f21ed83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb1c4bedad88cbdf555120ae98e477b4bad83b9e50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h940013e725bb70d0cc266a99a621c4f8c3fc4cc1dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144f7502c25e15f0ffbc506beb4290c6afb224f710c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9fd5f823e36cffecdf4de73fe469acfca7a8ef00fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6d1c5182e78047b6b00526fb30d0f039638bf4bc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he398a0ef4476baa6e8079c1ea8e848d641c9cd0c20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165f8924f085dfa4a4bea19dad6d9dadad372ec2d8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d30a6e1ef1bc7125716b7323249e3ee217847cbadc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b2d1e97cf0ad42353224c6c62368289a7998bcad4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1806d7c961536efb4cf0510188842a73b2bdd5ca4b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c657472e37c5a395e7d6298849f4af614935aeafd5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35de62b343860de03ed548b9ce2d2ad754b0d2bd44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19735a0bfc3706127b6867744d4303e566aff339e18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95a8b35b2bb8e4fe7a6cf5faef4e6dfb3390cbfd84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3f1eebcd686cc3606dce6b83df9739d13ea841fe7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193f2e24079ffbb7dbdbfa2c2b406c37631a6ebe718;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c902379d6689a3bce71bdc55ce767b41b1bf32377;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8351e003abc1fe5f02492ade02820b8f748251982b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133c63f69d46bab6208d8dde1085e1ddc0697912f7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110d4c798c1c2ce8c67173c544dae176a9f501fe213;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68e99e33310266c98c24746a562d2368910fdbb776;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ecdfcf04af2742b6b86190b81942b18f70da8a8296;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbe42aa6d3a61c3373ecc2c17c87a1357bba5d72897;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4617cc2d73e0cc0c470f64943700868d4ba3e225c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5d3045eaeb375c755f63633b349ff905965e19625;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9570e2877bef5a0a7b27d0be42c194b1b90fe91528;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1970d861e8afe2e822e530b8c373ead45f95ad1974b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d20567bd6e013ac138f2b50484372c4e2b44bb0ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5cbae83fabb37adcea33ec0e9cea24d87833e7b982;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9464bc396ceda168975b2cfec4e1181d251bfdbfdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h293fd74d43b2b78b4223b79a6e6180cc1a00debda9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h88ccf35e259d9990b5e5a4e19c268a632c086dad52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8ff2f77a21e84ad50f18b0d27081901dcc48edc81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd988cb4e2ec0814995980b01dbf367157ad661275;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h860b7135df04cda7df7d5354dcb56776a4db29c8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda42635bf8375dac94468915ca66c615a4335a63ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b01231c37c1f4d2ce0f5cd70f830a92ef725b8b8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0f41f973843fba9cf1539d4f5941785226cfb74ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c3a924ea02f941e0b34ad2133f6fde0a03b9c86f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bcaa85504f852566777c39de2bce996bdcfe3c88a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5cb8c9cdb57ca698845303bab2e05f02576ea5998a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122016dbc0df55e2deab4a7c58d429fde95895d9352;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fda5b5f11fb4cac418d454a2c53c7d186660ef1b6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e35b67e48e6efa7910d2c54184dabd54db75f3c4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee5db3ab35d15ae88ce1c41b867d1b1102f977c79d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125b091b83ae74b897d7b16091e89e4d81898a13aa2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha309fac3085ac76c61968c6d5341ade3a0773148e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a0c25e27f26cc27e19f575759e0bdb6f65637b877;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ceb5400d703c5979e5ed9326c464c63377e1f8d10c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81d240dec93d7f59c91f47e153c7d4286fde03c48d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a08b87e4ceee9467b66d1e14f2dcf75736379f572c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2aead4d4aa7e8c512078744e4c537264b82b78336;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ec6856aa5fa0e5ed9ffed8e619567e4364995b33c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd21902f12732754704bb287d1e780e6d6e334161a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d14b3d22e66392cc691f007073c9c5fc22e8bdc87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1276218cc7a00bf961ddf7390ee219ec7775d7fb57a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11caf0a50cd96a68f6e7cd5c17869add832ad10ab2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h112bf3bffc699361056b60fb9ff04e19fa60f210693;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb63e2218337d18afb59c6593b87a92fccfd69de0df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16bd3f46c92870cf5c6c200d1882645210d07a3c101;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e67afdc80690ce7fc5c49e4a295b2e36d5554515d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155e74b12ad19cee4836982b741fe2384da608260eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfca4983c68a6039e0cf92671efd5c1801e3ec596ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110796e5ab7c3e461defe4861c836621b8a4858410e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he20872944df1a8719e340e19d6fad46100e066b04f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3315f6ba8cbbdf756191d960c2407031cb4280b91f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b6a3f0f2a9143367b46bf8dbb5163ae10f8683828;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ecf2415b03d5f08e08aa67bd80340036c906f3b515;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1677ce3b969e110735f9721a73068fc917d59055b19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bfc01626ad86d996937e698ab7a285d78ccc6acbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1282a871fe3614f34796b4b34c0e8a5a3e064653a42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6acaa8e7cd3c78b5ea9a8c6c91cdf260726047a29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d3ea521e61029545adc3624b7707f354f27614d97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc19b49dce5610ad4b859f648d501aaac25e929156;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e20da1386e968b28caf1ade7caf41e50c19d99116;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ddc0a5067fbf18a2a649826edb291df6e8253dc282;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df7b27bdefd25cc6010ad9eba7f730ed78e7aa191e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab30d83f5dc5a02c48d774b6d928be2ec8c42e50c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138daee66ab8a1542f816e5db0e1ed2d8d763fecea9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc8e2af23e20ff07a7a899c35b8f989493721c7d027;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5b34b91061812e8db2c813dd8a360a9ab3d882374;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc467f5e6669e6f6dc26672b635a72438ba6e3b8561;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7e60b93f98b605027c28e06fecebad7801af349ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f370e00d1e7070772e10505717905326faa7d1a9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b7fd977ad89e4b76095aa5062533a5e4aed1e9cdde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbabfe6bac86aa446c5ed01f815ee7fa405d1ffaf39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a4113abe44b245047697f7b8665dc213e74711028;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b3521d2059a4f4340f8a6cb2fb8b56a5cda9304fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h629c6412e0f32b6a51ecbde781a0de422805b7788f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50afbe4354e310150df5f37e757f61819126833af9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4b2226749737d7863618753d941a2e7fe0a2ef7c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha12184fd687fcc83af544e8a3ff6f93604e48bf8ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19776af1ce0308e514e00e4ace1abee7d69b86b20cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174eb1bdc9f712b0e466e579bbcdb84cebec0f6944b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da60c73d15032bd5416e80bc4811a850fd5271d465;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fa04b9affb0083efdcf1fc1b49b5921c7f9ec3dd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha105c4b1c5c495a26d7955d56396cde5b9b8e62635;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d1e4069b377e4d8b3f7b5cfef79949e7f67720b380;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e6faf2d2e4328f3f7bdd4c3811afdfc7d32a6c6b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f180df8a48e48c397bd6b6fca5cc5274b459f90d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11028b0006e349fa4eed627799b8ecddd46c4822fe8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h896702de79efca687cb866336f4370f56b4f0e27ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h224bb9a99f98e9fc4251471e23de5d99aea60c4559;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1df0b9ea05f5fba1f101d93f94af0430d6e2984a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fd39970aae91b66427358c0beac24badb771fee9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f0e05ccffe8da7555a399d63077349536678fd0f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bb6c68a81cdfaab7962eb8818a1e0df14b90b11077;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8bc46215e1cac5d4e1efb1df25c5685fa20ab26c6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1b785400a8c786b1c501e5ce4a97dfbd6c7fb93de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97fd97270572b50cdfba444d67e3b5555ebbd0eb1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e5dd7c8625df70e3b96acfd4c08cd2d5e0f0da25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117b3fe6ee4d732620ce423169f3225005dbb9cb75a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1628580ba1776c220701e1e08fb43fdc2a9c6ceee84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d94120569bc07bdf5594285a2d8da52cc447849f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb372b34b69ccba678a01d379263d433b5b4ae64bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e79d22e7ad524d9ad2a4d773b51bf6b12ab3a99e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141e45d57ef42dd20d89058286885485abad5077cfe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1752990640822b7a47713a7492d047bd29e075fece4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h588c4b1298765565987bb021bd86b317669afe8952;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8ec5e1c7e36560d4cfdbc5e7e0379a8d1dec30f9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174f6c0f8243f51ee998b2056457f47b0cae2fcb0b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c55bce74fc4eca324dec87ce13cabb35959b761e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de444f9ef589cce432b669bafaf02cc642b92e0714;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbefb146934754c3a6a6ef3a1ecab46d429fbbda95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d781821db49c2b88372830c62a41ec25df38bf689;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb64862029a23f99c5463e808cf89338834f5612ee9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h47546bcd345354a2eddc5860694528805b970e05cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa92e94537eb3b85311536da879e805618867336eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e261152159b75827864804ecf1536d495da2c197da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e3b502afadcd8860e0291a264b1119114f28cea82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5e868a49b95cc925eeffdefdb39599a7515842b45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce778365a7d7411c64a7748dc0c0ffbb72d8dd9ad9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15fd6c412e14b6b67aa503d3b91e2e5ea68cdd96bcd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ad90a2b920d5e060c03782f0f58c6165cb7b28e03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f531ac03c6ed800b2e61f5a6ae452331c3cf63461;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193913d632927a6868ae1397abfab3527dc2500c6d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc091e3ee78ff8e9279b42b3755275ca1475e4c859;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2fefccfacbf2d4c1b8f8bca1cde54df2fa2677b7f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6a2904e9663853702bb31306b6d7e3bf72e1e310a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b642d7abedc6e833e1289109fe6801a3c1fc382efd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c739b5ebf6f053087ce7b10f93031ae4676cf6841;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e40eb348878f47b40dcca49215e45aac04dc47768;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfb6cbbcb9c2717d4f74d32fac94a1c72be63bdd747;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd1b8f2ad4b507421b3a4854e7837cdb2eb6193b86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf42c7b82d3666dc67830873a9e495fdc2cc6c1c3a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f78fa46695e0268ec067519f342b1ba94efd76661;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f5a46a6f4e611e9ca8950f7ff5be3222867f6d0cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf369662a691c33eefedaef913fa05dd03eb7c6eeb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7365eed328688a255bd18672705f905a79f7de87c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f59ed464751d90301f091041b3a6fde562d2305c30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57319ec06205d642ef1807a7bf5cf8b927c2b5e6df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d7c8884ab772d11e89e380672e37b31b0d81d7c2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb9bbfcb157805549f3427c4cb35eb0b9e1316e25d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h448835eeac2a61e3ae03addcde0ea83b00fb001b98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h660116b153f72916b3f992d86ad9269d8fd7a94544;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf7153b3ec1815c6dd14bf9033fa8a9d32c039819a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca4d060e223b4d0df3d91b89b9a6344691d302b9da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h395fd387b977ae12a8ee235276bfbe40bb03d12417;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e111c85d330ea583869009053927cb6151aa541fe7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha7fb62e7051a8299da4b86595433afe9e40a8c5363;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdde036702afa416e8a364d37532162dc98d377ca9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea07dc48c9f9143a434e1ac187db50876f418d938c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d191a2643515490d1f53a22459aba7320d33c426;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91f6476a635ba26e4415723539e701ffbac067812a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195cc9fdce1cbb4f2b46935a05e953e797de7b3e9cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h104057cdd06e2196aa2430fefdee82dfcd7d580a8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbbdbac4f6183653cd51e1349396d9d373c7e527f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6641e188f251d6d023939d37fcce0b27727c55307;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2c02362a73df7353ac77d1625e381df9bf0cb6c39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2bec9f641286edab2792d964d3dcb1e7b48c2383f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170c716a7d1154c18f8cb98a0d004fc2353e450b0e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h279176f680accf970acc9a10225b88d6efae5999b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10808329f4524f2e1e02ac5520cbd8d7f5e9d252f83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a996897dbd7a718afa1fbd996183e57d57d589e842;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e76c9415e4c9d2050ec75390a33d7f7903ee451c48;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2635cac7aa61dca3bd66fdb5ae05890ec3cf74ed80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6877c1f1320ee5d9706d806bafbc3575e97b2d99e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11522c3d968f021bf07b74644abc91397e500d25410;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1577aa49e73ca12dc3c345e083e3ac9d6be051b4df2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c4396de4c6b61d61049a10882fe99b78510299c09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f7c90f3764a6695194bf2dbf337ae2a1a4ee45d2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a1bb4c2d476527cdd3a9cf02689b4456b256f2dd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40ca288e08a1878c09247b0d2192d758dcb5cf2011;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b2b70661eb0abd1958778b25db2643ea7190068f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19cfc4455da371d781dfab7b3bbad4a14d3018996b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd55efec06763f71021acd0ec42fa5cb450e99f126;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32cd4a6ef0aeff0b76e904fc5480630fc0fe567895;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf403718710e9ef62a5dccab2af749c8cfe5a92f81d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195ccc4af4c9dc832d2572b44e35c2e6d8be6571efd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164c16d495761075b35dbfcb8d8b35ea0e2fc14694d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b0c54b9f108426d11a856e6e42c7aace42898d026;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f8be1b5a47738a33794120ac2c0247fc111fa3bb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1854ddd3597faa9767ae6dd009956629869c5549efb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h65f5bd7c129bfe184534bc9a18c2ee8ff6c7e15f1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf90239cff27fb482d9d6c99a0ed531e976e2cebea9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h562676aaa596ace4a29b7d7697b8ed2ebb999a0899;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h903bf79bdd2dc94ec245ec17f800c47327235dc69b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a1086ea0e9a67ef7f381ebba2b89506c68e18f9ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187c4c130e8696dbb05bc49034186c2dd97443e112a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3c7908b0db291282992c4bf8c1d9ee7d0aa5ec487;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h488aacec8be37012e42672aca060e37577e6404ca8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda5abcdee9e4a5d65ab8826af2dc9bde865b63fdf3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3fd0e0df5563fc02e9383b1fa9d9aef498eb265159;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e5827e5029698ed8b10d0f9f42a34382062479b3f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194822557bcf617e6877a0b2666bbb57a8875c65122;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d84b942b9d3ff3170d1ffd25cb18995cfbe026163c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0c137e7c7bc046c839d4f3f333fa00a66f9a52e70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h76f15029bbc661827bdd3e351d5f1d3492cafe74a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1267110d74d8a00f47a441bfc2b27b6d5c383a124e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18632adad920e9ca957d57fba5f342eb459b08a098;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h409fd2736b606c780f697c6f372d35ff29390f23c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc38341d100e6fa1ce593cd64dfa79980675c3be05e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a7a4e09f6a853a051a1469094c140b21498f11f69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148e09cdeebc9acb687f0edf622d4e36e4725264534;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdef92df9a7885f81ba565452da4a5995f8eb17affa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187c9e7a29f24156e42523619a02ab6ff13e499c066;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9ad64a64ead7dcd1f84e735a23b618008eca7e7eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h28743c5d0fc39f8e63744f821f05ffa13260984e45;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d0b03866ae8205aa9e8c861d71e848e0dda4be6f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had5c4ce15d9a542157e7c54b92c6d86bb6ea9473fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h37391c03bdde7abb3b96966dbfe6e336587b693816;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2edcf5c4c0b86460a5633fe612b5d271982475d84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18cf5b1f70c73d25b4d2d90d9a19a15ab6e2ee70259;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e25df121fa7170273b1323f9e44b4c358da0dbb575;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca7e82ae56ee6fc9b43b71567a3c64413b00af5a25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a68dbd716f7661132b3b975454b796dda573d48675;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h895c3e2c87f9c300317d4d87e4ae3dee248755d279;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca8ed484d43373eaa5b1eb00c81c03a0af2d7fe397;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1247d0764b0d45cfae0b6a65d80ed1105e11bc1f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c54c950d9eb20a96fd1973e8a0fcf52ebb006308;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21936d0d25812a1c397369f68c941ca959b7cf50b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13974502b9a833b1d3e8bf6a65131d92f5ef5378d83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bfa2f3aed4e5c7206b4962846bbdd7787015d0c792;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ebcec3eaf0f0faf02fd3739fa64e77b651b728632;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b74a6d196b12f181febcc6d7f60713c7f9e33f7ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ae174231ab2a19af2ae24475ac59d86fe0c7d21f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c4914241935351a1efcb494c9ae319a101440798c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a65f5e1909c167f1ec0b12b7fa412ff87dc31572df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1ff4f9b2c6520d7a985b634706b8dfc2f41317593;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1addc3ea68b0fae43a16b39efc608bf170f77a74b0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h177e3e6ef37171b6ae24a4a2e0046ec4cc09667f1f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b24f595a7e87b32d66cec890329d78e0f69240053;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h20a0493f2ca39f663d8b7c898e55e81903a2aecb5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h234d4bc1aaa5a65d3bc2583a7bb8ce4f72d50151a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a581390ef34fc8590deb2c04b86c3d112a06fa5c9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d93fded612fd904b7b62a0c1a258a7d38e8d56cda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h949b6b9a638fdf920188d16dbea0f71504b25e88ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1809930df99a28500793e0099497a494bcdca83e5cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69821b6dc57d10802cc65c7da8a6621cbf3fe40566;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b976de72472a41a11b5a37c594dc337a57aab80605;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0df1bf5c0da2f660b1616fafc2dadbefe0d6fb0e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d61d3a327dbc6bae6d646b011188f7af06334b6f30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1946d7735ade36e1715bbace750a91534bd75725728;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13be691226b7130c06c74a3fd00510ad5195ae3acd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195792e17b923f7b58867e300e27965ec51ed42d09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee43334859499c27a8c6535e8f12020a16907dd3b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2f7c96629630d83e8953074c1e17ec4327dcb9a23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d3f76133bd66cd4731d2f053b0761c6b85feb3059;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb7acf5e9b88c2d15b8f3d3df1ea84be97d6d071f57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd04653f9afe81a91aad8de6201e1f39e68d3ac3340;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1599fc7df211b1f78593fa614c6354c5ea249bfaeee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6523818cb53bdd5d4cbb721ebfe9054d153a702b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123195e96c0c7cf2a749a14da3d86e886db52f762a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10692f0ca95d9ddf83c38da9eeb9af92416a2e990e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c3691ba060420cd04cc927259bb86feb13935f74f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1adc342b8746e16e863d286610c2690e9972443832f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d3ad7a485a9a1cb1805b8e117efda0a2f50cf7d62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d72bd6f88d5ffc89fcb39d904654bfa9e019328901;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h114a1175d6801413454b5364ba4ea169e38c59ca2d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4e3684dc78a8793a0ed4e050c31e52b1be9ed5167a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c34ce051470f3b785ffa227c24f4932108601a0190;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17aa0b2789eb7aeeed72ba3e776fbd72741bd94d34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b85c73caa64ad3c05610dbc14067eb6cbe7c0e3d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac84a67985e42b20a344583977d87a0e4e75c657ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e0a9fb1c9b963c609f89123826b9058a79a7408cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0d2cdcb9fac8ede2130cd064bd3d13c6450179976;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae9b479344e148f05e9cdccc85bbad1c4386928115;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d8c01f73651056c1313181d1c72d9e9402089b7441;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b0ac86820b4c6a960ecaf3360bc14feae7020af966;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcbdd038f1626a3f2f8fa82dad622b641c4b50e3b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ca7e36437ee0be154e920b1ba034b713a513a4588;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5640d21f3da97f0b0c97261130b37ac51f9719c3a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12206f0d6a1f9654d50ac48609c699942d51e7293c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfbb65226535f06720a766925eaa823e8632a3da7e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d52dc02fe87ab777280e4d18611cd32f27e5fbcc1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116b0cd4cde2c7b3250563efadb4598cc046784728;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5dde99340c39cf71d8633d395eec6555325ab49d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha3dc0ea85fbeac1667de456e89e702cc39dcd74a53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hacfc1bb90ea40ce2f8de538cba74f931114c761d51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc920c6212119db0c0ac393a4a87e54b4c2088554be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a1a734aa45203cb77e52003781ca14e21cec0ed1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heaccce8676e6fe8d08ea00533fb72a2d0bf004adda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17094ab7469300ed1e3b83422a376ed5de1539d1993;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecd3f61e9760d6f96579aa0be12da915b921a97dae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a366a2130c959ea73bedb2b612f6d1820e6ec3e7de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc9fd50d500e4b5ce3001065b7dae6cb1268439317;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1676adbf8ed5b64e598b3ccd77dca42ac060be84064;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126eaf1c41f3145b4fccecdd36d001abed8390ea436;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150e745d31470a35ac137014d70b9c77cd63a2538f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h21627bf74a7d1f7f81cb68897cb7fbb79ab87ce6e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1e8dc0085a8626a108f1fa42307a380dcef043829;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc127e6513f9a6d1e33f57738f6f8b2ce7daa940e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c4d4f41d80ad0351cd33d0408d35aa676f7e63142;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bdea57db53f1803808928e87cc6dcf934f6e9b6490;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195644f2907fb53606cbc74ac0adc98ef8fa5a6ea77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c596691cbd687218c6a02d4068e04d646949c15c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aeb0c0de6b182e5bb18fe32aace4e26d03022c7989;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cc597de3319d2870d3a848af1f8c796fbc247c9b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b83ebe8a5049545e3d700a0de047a111d1baa1bc56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc91f3cec5dd276008dab605706ce82159ca3350c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3fbc3ab3689caa00970aa62fd264105e997f5bf365;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1614a45201a1b56393a0ee4167ce3933cef8b1d050a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c362f112da5bbc95253541a39285cef3f888d49e08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89b4d5973c9eb192baac52abbf108e618ef15da304;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d80f98341792b388c1174b48137b5be140318208ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b50cc31f466f565256f40d6cf7695b42b120fbedb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h149d213087846de11e3926c03d7d930b9222f0874db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7fb850e5cb84b7303658db3b99df0019d918a65f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1272d980b605a1221b90f062fe68555bbf86ec40650;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c72b4cb1f10304d2127b37d9134818353eb6a366c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he389faa75c40eb77295990b7a5677c4eb14205789a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf59f6b90a6c4ecb784b43abebcd153043ee58d93c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h919e19f7b367886185295d1190e1d6321fc3f86e4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e8ef7988fe1951a1f6775374b6aea618fb042abd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1cf78cf17eeb15a7b63d64a0142f3db16ea3bea0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd222d180e3a9b704b854a3a450a517b25cb9325785;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2bea80c375e6be28e3e6a78543574a03e15ec7509;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5c5db76f66f3fb7b8377f5ee0bb1e537c73487957;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e493e9f1cba24ad3f6e60c90c5f98b122865631f02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dcf957208bf2edc9c4eb96ebfb24df00b3db2eb15;
        #1
        $finish();
    end
endmodule
