module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    compressor_CLA16_12 compressor_CLA16_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA16_12(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [0:0] comp_out13;
    wire [0:0] comp_out14;
    wire [0:0] comp_out15;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15)
    );
    LookAheadCarryUnit16 LCU16(
        .src0({comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [6:0] stage1_0;
   wire [5:0] stage1_1;
   wire [5:0] stage1_2;
   wire [7:0] stage1_3;
   wire [12:0] stage1_4;
   wire [5:0] stage1_5;
   wire [12:0] stage1_6;
   wire [6:0] stage1_7;
   wire [5:0] stage1_8;
   wire [8:0] stage1_9;
   wire [8:0] stage1_10;
   wire [7:0] stage1_11;
   wire [3:0] stage1_12;
   wire [1:0] stage1_13;
   wire [1:0] stage2_0;
   wire [6:0] stage2_1;
   wire [0:0] stage2_2;
   wire [8:0] stage2_3;
   wire [3:0] stage2_4;
   wire [2:0] stage2_5;
   wire [3:0] stage2_6;
   wire [3:0] stage2_7;
   wire [4:0] stage2_8;
   wire [4:0] stage2_9;
   wire [2:0] stage2_10;
   wire [2:0] stage2_11;
   wire [3:0] stage2_12;
   wire [2:0] stage2_13;
   wire [0:0] stage2_14;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [0:0] stage3_13;
   wire [0:0] stage3_14;
   wire [0:0] stage3_15;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1325_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_1[0], stage0_1[1]},
      {stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage0_3[0]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[4],stage1_3[4],stage1_2[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_6[0]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[5]}
   );
   gpc606_5 gpc6 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage1_9[0],stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[4]}
   );
   gpc615_5 gpc7 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], 1'b0},
      {stage0_6[1]},
      {stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12]},
      {stage1_9[1],stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc8 (
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[3],stage1_7[3],stage1_6[4]}
   );
   gpc615_5 gpc9 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[3],stage1_8[4]}
   );
   gpc615_5 gpc10 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[1]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[4],stage1_8[5]}
   );
   gpc606_5 gpc11 (
      {stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[5]}
   );
   gpc606_5 gpc12 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[6]}
   );
   gpc1_1 gpc13 (
      {stage0_0[11]},
      {stage1_0[2]}
   );
   gpc1_1 gpc14 (
      {stage0_0[12]},
      {stage1_0[3]}
   );
   gpc1_1 gpc15 (
      {stage0_0[13]},
      {stage1_0[4]}
   );
   gpc1_1 gpc16 (
      {stage0_0[14]},
      {stage1_0[5]}
   );
   gpc1_1 gpc17 (
      {stage0_0[15]},
      {stage1_0[6]}
   );
   gpc1_1 gpc18 (
      {stage0_1[14]},
      {stage1_1[4]}
   );
   gpc1_1 gpc19 (
      {stage0_1[15]},
      {stage1_1[5]}
   );
   gpc1_1 gpc20 (
      {stage0_2[15]},
      {stage1_2[5]}
   );
   gpc1_1 gpc21 (
      {stage0_3[13]},
      {stage1_3[5]}
   );
   gpc1_1 gpc22 (
      {stage0_3[14]},
      {stage1_3[6]}
   );
   gpc1_1 gpc23 (
      {stage0_3[15]},
      {stage1_3[7]}
   );
   gpc1_1 gpc24 (
      {stage0_4[9]},
      {stage1_4[6]}
   );
   gpc1_1 gpc25 (
      {stage0_4[10]},
      {stage1_4[7]}
   );
   gpc1_1 gpc26 (
      {stage0_4[11]},
      {stage1_4[8]}
   );
   gpc1_1 gpc27 (
      {stage0_4[12]},
      {stage1_4[9]}
   );
   gpc1_1 gpc28 (
      {stage0_4[13]},
      {stage1_4[10]}
   );
   gpc1_1 gpc29 (
      {stage0_4[14]},
      {stage1_4[11]}
   );
   gpc1_1 gpc30 (
      {stage0_4[15]},
      {stage1_4[12]}
   );
   gpc1_1 gpc31 (
      {stage0_6[8]},
      {stage1_6[5]}
   );
   gpc1_1 gpc32 (
      {stage0_6[9]},
      {stage1_6[6]}
   );
   gpc1_1 gpc33 (
      {stage0_6[10]},
      {stage1_6[7]}
   );
   gpc1_1 gpc34 (
      {stage0_6[11]},
      {stage1_6[8]}
   );
   gpc1_1 gpc35 (
      {stage0_6[12]},
      {stage1_6[9]}
   );
   gpc1_1 gpc36 (
      {stage0_6[13]},
      {stage1_6[10]}
   );
   gpc1_1 gpc37 (
      {stage0_6[14]},
      {stage1_6[11]}
   );
   gpc1_1 gpc38 (
      {stage0_6[15]},
      {stage1_6[12]}
   );
   gpc1_1 gpc39 (
      {stage0_7[13]},
      {stage1_7[4]}
   );
   gpc1_1 gpc40 (
      {stage0_7[14]},
      {stage1_7[5]}
   );
   gpc1_1 gpc41 (
      {stage0_7[15]},
      {stage1_7[6]}
   );
   gpc1_1 gpc42 (
      {stage0_9[14]},
      {stage1_9[7]}
   );
   gpc1_1 gpc43 (
      {stage0_9[15]},
      {stage1_9[8]}
   );
   gpc1_1 gpc44 (
      {stage0_10[12]},
      {stage1_10[5]}
   );
   gpc1_1 gpc45 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc46 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc47 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc48 (
      {stage0_11[12]},
      {stage1_11[4]}
   );
   gpc1_1 gpc49 (
      {stage0_11[13]},
      {stage1_11[5]}
   );
   gpc1_1 gpc50 (
      {stage0_11[14]},
      {stage1_11[6]}
   );
   gpc1_1 gpc51 (
      {stage0_11[15]},
      {stage1_11[7]}
   );
   gpc606_5 gpc52 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc53 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[1]}
   );
   gpc606_5 gpc54 (
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc55 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[2]}
   );
   gpc615_5 gpc56 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[3]}
   );
   gpc606_5 gpc57 (
      {stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[2]}
   );
   gpc1343_5 gpc58 (
      {stage1_10[6], stage1_10[7], stage1_10[8]},
      {stage1_11[6], stage1_11[7], 1'b0, 1'b0},
      {stage1_12[0], stage1_12[1], stage1_12[2]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[2],stage2_10[2]}
   );
   gpc1_1 gpc59 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc60 (
      {stage1_1[0]},
      {stage2_1[1]}
   );
   gpc1_1 gpc61 (
      {stage1_1[1]},
      {stage2_1[2]}
   );
   gpc1_1 gpc62 (
      {stage1_1[2]},
      {stage2_1[3]}
   );
   gpc1_1 gpc63 (
      {stage1_1[3]},
      {stage2_1[4]}
   );
   gpc1_1 gpc64 (
      {stage1_1[4]},
      {stage2_1[5]}
   );
   gpc1_1 gpc65 (
      {stage1_1[5]},
      {stage2_1[6]}
   );
   gpc1_1 gpc66 (
      {stage1_3[0]},
      {stage2_3[1]}
   );
   gpc1_1 gpc67 (
      {stage1_3[1]},
      {stage2_3[2]}
   );
   gpc1_1 gpc68 (
      {stage1_3[2]},
      {stage2_3[3]}
   );
   gpc1_1 gpc69 (
      {stage1_3[3]},
      {stage2_3[4]}
   );
   gpc1_1 gpc70 (
      {stage1_3[4]},
      {stage2_3[5]}
   );
   gpc1_1 gpc71 (
      {stage1_3[5]},
      {stage2_3[6]}
   );
   gpc1_1 gpc72 (
      {stage1_3[6]},
      {stage2_3[7]}
   );
   gpc1_1 gpc73 (
      {stage1_3[7]},
      {stage2_3[8]}
   );
   gpc1_1 gpc74 (
      {stage1_4[12]},
      {stage2_4[3]}
   );
   gpc1_1 gpc75 (
      {stage1_6[12]},
      {stage2_6[3]}
   );
   gpc1_1 gpc76 (
      {stage1_7[6]},
      {stage2_7[3]}
   );
   gpc1_1 gpc77 (
      {stage1_8[5]},
      {stage2_8[4]}
   );
   gpc1_1 gpc78 (
      {stage1_9[7]},
      {stage2_9[3]}
   );
   gpc1_1 gpc79 (
      {stage1_9[8]},
      {stage2_9[4]}
   );
   gpc1_1 gpc80 (
      {stage1_12[3]},
      {stage2_12[3]}
   );
   gpc1_1 gpc81 (
      {stage1_13[1]},
      {stage2_13[2]}
   );
   gpc606_5 gpc82 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc1343_5 gpc83 (
      {stage2_3[6], stage2_3[7], stage2_3[8]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc1343_5 gpc84 (
      {stage2_6[1], stage2_6[2], stage2_6[3]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3]},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[1],stage3_6[1]}
   );
   gpc1343_5 gpc85 (
      {stage2_8[3], stage2_8[4], 1'b0},
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[1],stage3_8[1]}
   );
   gpc1343_5 gpc86 (
      {stage2_11[1], stage2_11[2], 1'b0},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3]},
      {stage2_13[0], stage2_13[1], stage2_13[2]},
      {stage2_14[0]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[1]}
   );
   gpc1_1 gpc87 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc88 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc89 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc90 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor_CLA16_12 compressor_CLA16_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h60995df0e0f4f6fee930f473fed4f3fe8eea32400daef13f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcf1f63f678fc3598ed49badce48f927f1b6b319d188fa252;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9527ff7006222951f28241ed3edf93dbf78c5606a65b70ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7eaeca8a916de2acdd07a153aec2968d7b0a04d2de835072;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he3f15059c3bceb260a8587350839dbfe661a1fa84e5c4213;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h378f73bca49f2fb913c65d230cabbc26bc152a534850ef41;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha564e3b21bcedec97f53452395731f8bc68cc8c9961c2a16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h748c20c5882e3d809e1982fad0f70649743a1292587c04ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5b9c2920de101e153d8155041a9349e35d3be83ebb089164;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd166a60a2cef96d82a16e4c6815043b12b329e3f0a4b61c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2433dda3a6543b55413a92036ff8c2e5ba2f6fc6f6332c1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h43a10d57be28a0e2103c677b8e2a29f349f485eaad945766;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6b72aa98d35e98c1b89225a233d1157ef41241550245f7a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8be1020305b73cff75f79927c60e8ed2992d5100fe852b23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he70f4953a169864485286ee34e4a07ad1c1e43416a948f38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9f48bfaab409572cf874666fcdcc7e7d9b9931b3a43ca996;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7765c36d166690a9a4e2950a6e94881d9b2c0db2ee8a8b0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hbfc147b3f7256d6fe06f0e593cc137a7f067f8c46205d76c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h973cf38c7f88b8e9f22ce02f49bab073a42a2659a9a10e7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1ac806f3c17362889079a850a5516a57ebeb43cbf76093c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5f97fcd3404517764734dc9f02c442ab05ebbb0890ce68be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc4ffb7c6e269d9bc1e16fefb88f59e4549f578c6649167ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcd94543cacaa984a34d3f082363e78aa8e680806a43608c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h19a869fac5f740f8dcd968eda7e8b5b01895fc8652c46b48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h555a88f584698024bf556cf4bdbd855ed150bb4f160f2a73;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd4991b71114605098e18d9813c6f30ded20c45ed9901a802;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2a0d0486b58c72045771e34defd163368f455fa9a8ca2e09;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3c40325469d50130b21313b343782ea6998a66d819d6fa93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd316eb036f046c3d054e5ee1dd5e2c075adea03516bb4802;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4d8332649185fec0096afcec0d5536fa24ca7f7f81d829e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb743d7335495be6b32dfa67915243fdd994648c75d087602;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h76c2f24ab00d04036e5f2d3afcd15bc1d225d5d33e5a2716;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcd5987e16f916815ca1afef33f9165a0032407e82cb6c6e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h170ed8263af71ec8545a9ce2c10df47e5a0ee5eef7efb875;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb003f523276b2ff020181fb542497f2349692356983fd448;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h95bada8642dca298679bd82694fbc59a128f0af71814c4b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6f26898a59b0ca3740200547811c711f3fd9ad459e8f22de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h644592edf580b455498e812bee735d02b14dd1d92615c24c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd13e4410382e27d67ca00b8f883059d9204d2e0412d8e031;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h252162fb76440a4a6e51918016d68fbbfec9cb909a63c46b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd3cff36e2614df4c98f17b861ca123a42c96637a45050412;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4208b40504e099376b9e34f0f0266bba765e25e9406f2347;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he6ed569635a2546525674944a902a556308acfd45c0dd59e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he6fb30db0c5870f600e363c692001665395fddfd314ec78f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc8b9ced1553eef60a43e1e5ad11b35d3a884fe44725a0b68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h97cec261ca88bcac7e023be80667ee510c3443c395296c48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h576a4861757baa8cb1a3647498af5e8ae0f330728852206e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc8958e6236b13f828b49cf3201a49833665a3ce6bde94562;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h50a57de16a61f8daa41ad31913629ed83d405a51ed344b5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfa1bea49c1d5f2d43d679a3fa8e87ae7be21e07b2769fa66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3f7000bc328e231e8e46cd8ea1ed8ee5accd80dd9ea43d2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hae574872c533b3dbe21a83b78ef289c9c9cfa9d86c583dde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h67b3dff3f226b8459318eb97e9d12fd3e7d8f93c7afb0165;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hf27b491aa1a726eb32673877a8e0fa4f6e6a2c1ccb9319a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h549500ecd9a22f6feaf1246cb98749568dd3b60599a86516;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5fe63b5051aa215a6d881c4d5f1015e10a01e3f2739ce6ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hecc2f9cee292db7c8296d5d073963485128985c9e787f916;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8038d1341868538bdd4a5ef589fb0f2640479d8e4eba605a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1f3ef074b2d0b80b7e354dc54b98ea17bf9daec4fd918078;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3d17d33f1b0a7034efb358a5c89a640cad81b0a63fbeeb4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6604b7d633604bc96399e07486baa698a8ce60ad1b582d7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hbc1b1fc6fd3c9d7de84e86f18fac8fce1965a30a4f5ee0c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he7d42c8f9bc0d2b6f18217d4993551f51bdee79807414e86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfa434cf4f8b79697e45d0bfcc5934bb78a9706cd714646be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4b8c55f49ad248912f61e312889824a2c168fd4631585c7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5be865593d741c18b8930365c7aca752a8e72468ca03ebea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6a93dac47eee1447e56da16119b3f536c4db72c8eef0d8f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd1d6e774359b8ae8b10de688631938b9194389b4f3fe015f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3b6a0e3bc0e19e155505d64475bd02d809eb4011287bac50;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2c8f945448296765843ccd8a2979fda08ab881aa25d4c99f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9a8a7c8ad66b8567df6819b338e70cb9d68aa04d317353a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8cd5a2eaee0e589f54fb6092d5ddbd663f8aeb9a92a0cb9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h51e6fde667f86a8326bd0d81f3cba89689b824837b3386c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hef6b259c2975f6effc48db8b7d683a6ab6713dc4fc747597;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h79f70e76f7e12c75d7ad78817fef18470666b8b0426f1dbf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha5f20b69b55bc067a1e41cf8092992f4e47954ccfb13ab89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h46c72cab067294a0e36e3a16b47676a23c60c5ce69a7dd58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'haa6a81a35848bbfa2d834f512983594f7ab7cf4f023c36a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6ae5deb03cb8b0454161f080dab32bbf33a90b443ebaa4a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hf57dc4b3ec1e08e6374ed8d992414e9714251c27fbdc2e3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h14477646fb5fdb32f55298b9ccd98ffca3447926c6499148;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9ef03c1823d4475a1e46428ee9f65ccaebd8b2bd12df063c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb016141f6fb8d32a759fa06ac42de8cc3d6d7358f9ec102b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfc324960696cdcea1270851a3674e57076b6f61f036079d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7c0fd4a422f2d5bbf8b413c1da5ed614fe3266fb9214958b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'heaf4c889a31e41cb242d6c78ebf13ece29af7269e6bb2512;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9759c796facfe016e7b8e30c3b8dd6aa7bba64df5a16d876;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hf9a0e6d86df39729f2412be37511f9885555973ba61eb1c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8230312d023df60b15dd0a8bb7b1f8b67ed1b9a82452b916;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4f4e3458625ce7a4502c6c02f55de6ebc0f8b6f32ae74c97;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfe0cf4ec2b942c84ff4bdd82e6d8e36f27b278d52e3217c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hab8d71b57e06e668d40a5bc613f4331610550c241bac8271;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6baf423c71c58ed37f9b934c5a039dddda38b67b873d57ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h370e41011e9f95ad11029fd82bcf763e85ae167fc3acf53d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h47ab04583c9ec6cb1474cfbe38686f4f611799bb2493ee6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9c02537b1b74c4d046e60b894b05cad3373763552033382d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcada4b12ca82a5342a8dc6388ae616d89f4aa4db80c665c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc0074305086c893d58331d42e5122e7f0d790a1568519278;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7da8dc2cf3af907f862f9e34a8549682afb26412428ae2b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he45e4fa2406cf113d44678a9869adcf7dd72a0fce6b9eead;
        #1
        $finish();
    end
endmodule
