module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [29:0] src31;
    reg [28:0] src32;
    reg [27:0] src33;
    reg [26:0] src34;
    reg [25:0] src35;
    reg [24:0] src36;
    reg [23:0] src37;
    reg [22:0] src38;
    reg [21:0] src39;
    reg [20:0] src40;
    reg [19:0] src41;
    reg [18:0] src42;
    reg [17:0] src43;
    reg [16:0] src44;
    reg [15:0] src45;
    reg [14:0] src46;
    reg [13:0] src47;
    reg [12:0] src48;
    reg [11:0] src49;
    reg [10:0] src50;
    reg [9:0] src51;
    reg [8:0] src52;
    reg [7:0] src53;
    reg [6:0] src54;
    reg [5:0] src55;
    reg [4:0] src56;
    reg [3:0] src57;
    reg [2:0] src58;
    reg [1:0] src59;
    reg [0:0] src60;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [61:0] srcsum;
    wire [61:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3])<<57) + ((src58[0] + src58[1] + src58[2])<<58) + ((src59[0] + src59[1])<<59) + ((src60[0])<<60);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187f97c587d7f182685dfbd9299c7b2b290068ad76a1f78eaf0c753ccb2132956a31c83e6412ea8d7f7df503e5ab6e5e0625a6e6011b83375f0f78878cac174fbe18b40878ea1a0e298714fb3fea9e94882a0c809fc8f6231b0476754655de3992b51d1e71f48e97e8152560dbb5a8a4f9634964c64deb606;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c145f82efa3daa2fbc3f7759f6577331ce4f27a2f94fafbcf2ac972550420588201ac914cab9655a1c5972363ed54d8888e8fdfdfa7f181c25691484cac34e80fb9903361d6539a5107bae11ca9be29c45394d9bf92ab124228353f0e9bf1b2f86f271024cb270b090d64627ab27de38f9cd9c4a9b2a574;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfbe2fa9834c9d744d3ba128f6cf239e3f80b2313fe90b6f09637756cdba32b7ea20bbdcc8976b131f5b5ba2e6c28673e4ecec3f977883f10c7e179cb9309f9242628e22e2270391f2bcdbdc09afff8578027a70394ab639345edc020a7cc9583410403d79449d4b911810fd03513674665e8937d042be7d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1133544903ce014d5f1f415d5091602ce0472ae01e0c8ebb2a7d5cae3d49987da3316a15a89eec0bd7edd20ceee90e6facff234765e2526a24b548cd7e5b43d73c71a094b2b1988d70347f3a8bb9777deb21b4d2562bc453cfdff12314003ec12dd205a28140c800e0ad46f4c463fa83249e26497c3e2d601;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha307e9ac66db0bf7cfafa85a1dec3724c512563175fcfe5ddc8e92d248108314a1311baefb3b48db5f0d177383b13f4714350ae9bd3c84f7f96c9db56028c023b8a230c4aefb7f3e1c5c77d1994ad599ef19849f97c1ca58ecaed0e8f7da6c94690e7fb75a7fde8a08eecfd17b1d5003dff3e7091b5297b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h995119e8ecc0b138f3792ae3b1bd656ba5b8e1bb0bebf034a52d2ebee7f64230f7d3ab086f15f0832aa4dca5f96a218a52760bc66839a1eefbd2805e03d2065843da622c4682d782586107eb9c86f0f3269577bfb8dfa60a88bf6ecd296dfc03d72494fc046fd4a53442eaaddaaaf038917a860de155b6c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3124c9c11437fe10c227f69e1005b79b7dc91e92f893e07212f2cd999771426ba8d8212e7fd2918d86b2cd1f817a63fc6b1157c81567843303aaa2d20b0a5a4a88aa3c5fd72653e6dbf7441f5370216fdf3aae7f3ecaec17e6a6b0a1185a419002e4e31c9424aa0fcb5ef5738b4b211221685632d313904;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f14b0cc9c0bc7408be198edc31d7efdf07db72659339591e0b0e48e23235412f83348fcfcabdaccf8fc92001617229ff3b7ef02842df723d9bbcd1ee52953252ce4e711e8770935db6bb1f24a43c62a27db398e51f6595e1d1d02acb5221bb509808743d971b80fa5943b73b5401c7191cd6d63a18782099;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1399cc0fd2aab9e34e7200a8f8a115a2261b4dffc1ae9171aee61ab1655e73bc7647f0dfa259284135181410b6bd4c9da1e1dd45d0cd30952dac6cd1c6644c4053dd062bd86cfd0e21dc34202aa013fb36b46d2f577d1760d1aa724623780b580535199e470551d384eacb834fb51ebf0e12edf0c0a9e4274;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3e9720d2f4605844cc5201601564af4164e25dfdf4acc7d4f68854b938b22f59df022db95bc72169ff2fe6a3ac9fe9ce5715007268ac859a4cf2c2affe5ba773a936e111ccaa7d5f6cf1a4d57f8c6c1449a9831ef5eaeaa0feb9aa48a82b67d7352afce7d007195c3b23d5f87f6339f3829acd2ac8edc0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a29c55778208a705afa8d6ff57a4c03a6e43be47871b39bedfd54b5c9ce01ef155e82f142321b71aeb29ce9d575e51f6c80756ee9ca6c4b2fa70bad69f175e66c6e2151bda4bafab71433e2e8d7fcd5b3136cf687a0727dd0dd13fd4ae34ba692fc0072a1a228afa9329ea3d569ede6eaec4830ae64ae62;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88dcff170e42804ec7e848669cfc6b89100274979b79c034cc719152cd9bf16016967329305d7d4b87d5b9abc3bc10dce2ac7acf38558eb54d1d9944a41979ad298dcae85d9a87cc89322851b8ee314c9c3431c0e50ddf1c3b851cdf85e41be454607b512d69a4721969bed69a31cc4dab7ef1a28e89c2a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebf8f69c9e7f16fe13e3fbfd1a84d4c81537d4552ae4ae56477939680be00f4dfe899ef934188d8240c22de89fcc0cadc3d9be68d2c5ae671165b000337347fa44942302060e8dc699127f0c1fc301e1f4ac48985c62b41b158c6da74c031d6daf2ebe3482271d78826610786de4447d028c419307bd9166;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce9e9105d4158476aba4a55b20c6ee4e9c5b52b55a3c8ab722de3a04d50f50da3ebba7ae180caf1ac566bac7de14684f8ea162d7f73fb4bbd95f9e9b6ef5f0ddaa21112ce397294da987fe0a6bda4a6b8ba318a00ab5e8d0ff1a39e282a92dcb016dbd3d79ccd39c3e4e54236d77727efdfa47e93f761bac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfbbcf0e32e91af67d2f4d7c5eebd2478eb71b817685a148df346acc2e99dd9ca4c4a35adbda1afbccd90a55a5e624936ebeb2e810c78fb279eeccbc4c9230ce970ba67bbf2ce772a2e53ddbc43d492d1717dd012399c7915fb879755ef6a92efb089b2b28860e20a01702a57b122ddf9c2ea9b23d6bc0b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1767d1e941e9503e02f4c891e00c3eac407300cfdd32ad0fb2829755443489cdfa8f5eb82e4291ab68bdf3134e0c77cd41350343451b0d177f60eb5540c5fe5a66103a89d88d51052eeffd3fc9ee72d807720cf5946a6231fd7efd1ab37c50649f36e68e57ee7f1d27b7c331433ee106a93e80ed89cc3c36f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8c9c20473f92d6ab67d25a8cadde6ac419a3f291ac860717d1b88d118c5f28146b6fce8a988849c328fb9ac1d14ae2bda8a87639c076f8e0ada7e6a7a94d3cd37f21d667267129268c4ccced07984897e22039ae9484966f03512e074f53afaa575d727b0d150d0e6f6624f7fec1117531257718dac7af3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5d787b7aa24c329b6f79b07756ff8778a26a916f52fddfbe1b547f6a09c6e3671888dd5bf4e769c59a7da20f211023bd25135f6a22c86b0434264863274b6baecd70895362673118e9f9cb4266ecd43e5383ef22991dca55c30ba7de1df58d7a26812805e47022b640745545da3b8aae3def3d5a4d20e0f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ec803c186d7f830fbc8a3a2cbe0233a8a6183ddda9c8b17db4e37dfff852b5a4a6723252a5c67916b86fe18456238e3c413fcd88b0a214b4b3b2bdd351ce739aa86045e78a80c7a97349c8a847177dfc5574bf6e1a4459c2c0f47e0651d282bc1327aacfaae8805969073a11658c124823f8af9fa081c45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h817a0eb1bc7bfee977eb0ddb6a156a0ab4f409447af6f7f5b46c13ae524604c83933cae34be062588d2c84b63b90d149565b32060213bdbdc9480a139b1f8a3f6f28fcc80081a3733a024904a53eedb7a72b640a545c33f794ccde6ca50d33f7d39a67f81c7eee6c9539cb3350ccdf4866127f05136f6993;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef5698e82ed528a1e26ca89b1edb186dddca0b33f8cf5428647b1b8af19b53665078a0f04be417db7e5f6dfc74c45dbce313c4928e24f2a22505f7ced4714cc3e63348e2b5789d2f93e3372795dc1389d80d26892700ffb4519d731b5a357b39ffa5a7cb2bb9de1a9e4998c09d31e9578a42d6b03e8f8da4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4bfd55e920fb7ad45478a72f592ed33ef5a6900366fa742d92f5023aac7fe74727fad0c83181dc06c664199cd06b43d686fb18b80fbaf643918e4d61a128080d0c30d60fdbb986c66ed05e88d7c79b6664d9fae74330e6af41ccd09e926c4818b41553575e43cce6f0deb82262b6d7219821df4a4b3216;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59a2ff6ab1dad48380f490f8e00745e88b73ec11317fa1ee0e18d448fb7a688b7a62067961bcd4a1cc843212c1f726b2458c478ccd26dd2f68767c9eeec2d57f8df63547a900b9567667b3662c6b6c4068af38852c1d98478762c76a6ad61374e90e2299af63b3165ab39d64c10a375883034aca72c0cdfc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31dbc47c76b56bfce2afe75cf9e2a6800ff7469395e4cb3db8695a1e7af1c008ba28a7f7413bfeafca662719093097e3b3ffd21f2ae4a42a400b5a345bef89447bd08db336428a9b8f96b3e91606f6d9d3c7c2e8e5112ae3ea80934994d1e0cf2cb35756fc9ac998465bdd69dd736205cd7402ba1fbe8edf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1045a455dfa00ee0c1066f1310d6ebabdde223bf8d021ba941040943e35af06ba55dd756aff58d2b69f58e5da1e5d86a8c07c6b3c05cd09630292d9becd7446fbb1a895b3e3021dfe40d6b070e2b3af6eb6164e6ca97d28fbe081c278f4db39c4e98e5cb0c310b2ad5acd2f460e26950661b8525f438b0379;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacb92471ec9f370f4251cd50a597f35001a9795e9226bc55c4ede0a1e472b25401f04a85597bd6938acd67d13cf2abe0846f7a27e69bffd67ea3b183c5fb601d64239fd4e36a5bf7cf33800e937ee29f1c5b72a66e19b5c9364b6d9fd63927a8a0bd986a306a2309accb377c707bdeb32ca848425dd4d566;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2104c075c9556f084f34a93e43d0a84606c81cb8f3e4cb2f41b98e96ec086df283349f3ee3e58c2655622fbe335fd45c4acdd4029b62ea9f4ba4c2a415fa4924bd544292b7e9eef0f460200a1b74e83d8be86e69c86e38a4420eba4d33fe380aa85dbcc1064fa3c4148fe05ecc694b203214bb9506a67f63;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e5a4375851bc3e5345a9cb1f9ead6599052a34d774d5d92313b76883ca92b82250817dd27a85c4ba7fa9bfe0093e8a4f3b99b103c69aa967e29a803d9939d698c69bd22f2c7dbd774e4a1dded2a2012d805216158f207e0e77df2b26feea51f852650a1e8f3702acfb9ccf26085cf4ea0e54475ea2e53dad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141452d5209fb074091374da9c322627757053d774e75b720df5ec6085235199c416cfb845bf043526e762fa9605a4e104125cdb26c0ad6d2d6ed98d6598b1412ca144023ce2a44b6c0dac5adbdbe8684050557539b4bd81786b823a98c7680b89343ba9e9be829570f8865e850e0a43de5f279958da4eff5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94a38790c54878bc1a9814b41a964116516bbb957b64bdaa2a23547e5c2813f70251bfc62ecd58fd014ce94cd22a730a4e5ac441b1fccee5f2f681aa7de72e7c1d8e4182c338bf7db161d35added8e029117fc52e52594caf6e1694759ae0e21ef368cf4543f0f9efd56f6678b3dfdf5b8861f959d184c45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d5ec8a3f6819573f42b123694c2835984da0f12c88006aae0722bc5a902d46337a4898323039d4ee834e18edd4ad37451deb84498f1b41545ad906a46abc216cfe8af1ad368815b9cbde2b349a4ca4ebfa5e6c074ff87d249cf349e3cee78c1c72e160aa05cf4ee614dd08216ae220cabffe69e261b20ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0c161dfc374d2880cb8964987df217190410cca5183be7b22085e4ec9218ca1e4dba4b1eaf9473c5145f28f3181e4bb3775b2b045441fb2ea3c28aa2b40d90eae2137388c8dbb15c19dcadd9f895c9367cd6b989a342d50da639dd01b21c08432b0c94154168403f9bad0cc567ad7bef9b245a6800f30c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19614764d97e8c565a7b1e21fff3714f6cbdde3ca850c40592c08902a95bec9d3f7fafd0086e8aa6a05d8e04d00754f86470fa7224749231a442eceb4e506eccb013e6ad9f006920dcc3abede23ea7b271820953bbd07f0d5780e8c7645d94ddc004050013a80e0f2ab5f7c864049ee48568b7b55e9c2c430;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117ce61fbe9f7223d9d835d50cae00ce3234e25f13f2e2b0b85c741fe7e9b8f298e020d9f7b742569afffe4f48b936b071dde2692fc45a9d18cd535f33930b3120235aa4014b2a24b3aadc0005c1deeeb1f71552515a87ed496715e7cb8586c68026da287169f14a5bdb2eba08434a6204c8f273c457f606b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fee12c0ea0cea9453cb8f022c10651afb8910698264b4f26d6b1be968c75763318f3c4bb8befcb9c9edb262aeb0b1e6ab1c0204de33bd4f1836204b84014cb34a0d38440723c3ab3bcba748a34ecd4031300a8570c6df346a2a62c47f96ad0dc8518cda8a3000fbc9aa1df2f74d9add177150763e76de790;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110dc43d679a30c54c66ccf46b3712754fb008e5a7f4dc9dded650ff733f9e6ff6b836b3f260eca1fe4a85ec3e3a7faa844a0be99060a018d7d44556e966da8d9d17179709662b54c81e3fe5d316c19913f545f0fe2b6998924fadce7764ef77ab96ec952587e1911361c766fdd1d1887afbd353c7ea88409;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbd6546eb8b529cbd1691bd40487649d8c6af7edf47b56300d1db36c8167768476d83f98d0f8f783e5b4e93ed4ccc2a2d0527d59928101fd4076c64d99e17d73589548d090b681892b573655b7a3383b0db41d6573794f39ddf6acd93dcf2462cfcc0562803b3f07840f8550e33e05f0a40c0184429156cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h959549af3d970e87b949b5266d2a9bdbc8cad6f70504d09173235d709ecba5dce9e152722de51e52a8643304304c000f2822122254a4074c0ede82b6aba0e71be079daae6125d601ab25ebc2236db230f8c02bf69edd2c364fc30aa06d1d9bc85a1cab6937a89f9944f5d9902777d7edf635f47b3b144670;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdaf9bef37365b524522d1d3b5724c43a8f3918eb63dc238c50ea6c6c9c60d394293705497b3fc38eef543bfb82c921a0c5c15ed8785a809b7f809422a78d0eda7ad929bcd002c473f8c9adadbda22b85af9485aa11b8995b3e5ab359a06effb72fa2d9711d54c80578ab425d75cfa0ebad20a63a49c0a762;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157b55d793b51974ea1936037312f8ba0d770dfd300bfb27a4f5ea0b8e4e9d3eba99f5dbd483d1a7d40002d03152653438502685d9c91d44f55c68ab89766a1a4d91cb8530335f1b3ac160f1ad70feb1d7639545a379a50a75bc2134dfb3e14e10c389a461442f866a40a365764a49e4c626c96fe2c5eaed6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9de5d2acc37740c452101cf01d027847e8af3a36722a184f6d27fa6d37611b7dc752d30593cd5c6f21b834a526ddea6f24b362b6b4ccce1a503f390d6247555d42af83ebec3c648a66f1e2c75e67f5ff6ed9bd90173fdaa7d7a1a3f34183a99ae0066b974a9aca258837148ff87aa49542c8bace5c71e7f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1def511ed6eef1da12886131b9508efd8b5f11143790fac156f2591dc54a4d5178980f36d09337edc6083141100e972e30c13b0c33c8ecb89632a99258361caf738d30fcb5e32edafbb515a3c67706133dd0bc1aeb11e695664753268171e2e68e9d28d321d83280b1ab916397f804479978f59de9d5bebb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb919d735c302b40cbb133561b2e362e8fad0ee2803b57a2b6a24c922f98ad24c0b8572730da5c4b40d08046928ef6058d48656e2a81eed60609d49f102dffd0f607cfd8fa53464c5172c027382ed349a174b1ad9d1b954ec8d3e944d636a1cc68f7048e05ae78d8e325fb26799ee6c7f3f2f752370ec312a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15894e2b0c5ae304891e2e35488449a23dd22a854f16dc8d59211837494aadef5da70e16fb2c308ddfc7507817e7f0008b9e5be62b6bfea042f398928c0fa1aeb8786275892523c51663081f9971d215e0736d49d3e61fb0aa9f892667fd791ae87bea177feaa5531879705f3ec62d5883354d8bf118ba8d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea232365cf550f7b7690677fb21126e98d2790b80c8ef8612f628ad7089c569c8a5b15313b6bf9350ea8ffc38415c5cc64adb2f61829d42698550b4b64cd00866a9abf98d7127a778d783a5a59fc203d67aeefe72c4afd5fc749439c763c9784937e5b39dfce9b5526587bbe9cdac6813a6a4704ddd5fc26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4423b5d85e5d213f262a2f8fa86967a73d41e7f19ffa10aa99c590b46cf0d9f4889c4151c19fad7200210f62820ff95bc1b95980ce7c6ea57f1a99afedcfea0f68b24b71dcca12d825eadde957cfc2fa31c6727feaacb7affa798d44d69ddd1f331858e62ec3de948101916dcc286fccaf7a8c31d596420;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e26f22deed6dae63c07a696c846548c8e35d79596bc38c4b57ba8c4b9f85e0aeb61ff8ea6b3ae5401fc3afd1227db34fb7093e99e324c90d65d77faf840e7d290aae5f4511b77019e58598e723466d82e79594ca4e076cb7c0ae3036f9db15e98cabcbebd725dca3d9427e3e9c25365a606211fe024f94a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac0c19085a08abe7eb0b56ce00dee20009a8ebeb5c40f01be270c7f2477b80bb4dd561c129208e7e17f4e20ae97964ad7dd5bf61a33dc1e78eeb4db9db24375b64a2e317972d1116ce06c291e17c6572c288e8a54193a4e80d788f42c35750b4fcbd54aa26e963b89b88b9a63c19e839c3c541d0d6a26fb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18ea755ba89af45dbdd4044597688d6e21695dbe136f1cf7a917294bfdf0985e6c5167a9afb1503b2281495796d6f9da65cfe048d520e7f815604aa20136ad74e35dfbd1c7fe0c8725227a5a9e01e61a9fa91eedef60f52c26571d99e53f019675160d30672bdd1553be462cc74c24dd7cd6fa9921725fec6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146ceeb0ba8a0de87589718f02dfc0e41e09753b9338bcdf914f0803f51003a7937b1479b53e6bb74415d821ae243d546f254cb64e66fc456156dd8451d8f91845199693cd57ed82e68d6bc98b11baac99e500386fcf5df2dd43699637c3789a4ce736997af4eeb90ffbe13e2964d0598962a186cc3a20a47;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17116ac003430b4973c61d6a2898f95ae1dcdd3fe02415b626c1f5268da93fcbbc9e7af78fb047dd6fe856b443bcf7e8dc460cb308453e7159a07696de34235c3f7c26cbd95e8d091f40eef6e64ed4206614844ba1e8a90f48adfd7ff5887b9e3ddf48b3dd22f56c264f8d4b1ae556c6ee5efd22c6ea4051a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53ab49c19ef3f9cf1e0d4ac8fa6f0e47326b60262e86579ebd46388fda6028ebe943c1f7c2caa446086a4340dc522b344a738c8ea81b8fee2101b6b9f503255a02e7d6f68ffdc73b120343ed09926bcd2ce0da1c280f4b92abefc48311a9560b997559c627a9802343ffb7ab66719d4b3d94100061f676ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h815a5fbf7a924f441b6128965595b9e6927b13739f3ae6c7b2c3945c288c3c08c01d19a78606405606ea216b5fea6a6d7a195af9abbebfb59a3881856c242da16fe3a28e2b7a949e0fd2e1c4b53d2116479013b90069dc99db533817f3083141d55847df23ea97a7e72b5c6d19c65703b2e31ee50391ed14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bcd6c6a3a6cf6ba0f38f4e15a166c60545992b39897489960928a3d5d54db619fc6fe5f4e754af1c98e1c1d09d56fb85f13bc48bb9e77a5b8aabffc4dcd908c49952fb189dc7c5c38eb656474f8e55588a757f373c618b224564406a7d4f0feb79734dfccff8f3c7ce87a77b006669aed4525ddb90db77a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e7090d5c439a95ba6774a143119306498c8f4e315775a73b4c811860b5799b882bead3eec5ebd62846b299b74ca0441cd2085f37e7e77611a031fb140ce68a65280541bd9f88d0fe7fe14fee439a00aaef2f7cabacdd1f5882e92fdcaa2fd9d58387f1a4f4228062d15bdb85f15c4cc0a0d2bca7130dc74;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db634ba8bfc96fa6a74f9aeabde010d26171cfc4d22cde9c5648cab792a1df64ffcfdc176e38427124c51f3d00b4c54240159af81f3fa5fd5acccac5a2854be5add9c50286a4bf99e324a74669a9537636b1ba681bd94733d85e2f9a9a82c93e4ba19fddf4a2101592cb76107848465e039c6da5a722a94e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d92e4b76703e182ffc2e90f8bd69d25ab46d0210bacf67a62555e2372881fdb2bdab449ddecaf2e86c9afef9eb790c97e8017dcf6574180d6856460003f0a72ab0a56253edefdeaa708e4e9aa6c3ebc089ae7173733cb2a78ce53189dd03cf9f0641419528f02816cd71f142f4d1f57ced947c110ffc219;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a065c46aafb63227119a71453ec2bc6fdc0c8ade674142468b453fc9f68838bcb229dbc1822e26d8982b64ab06a306c293e3c9761c2f065a8790c6ec85d86d96b0468d4d44746656ea541aea34a4bcb83582da7067a36f757f8c32e341507bb67fba28dab72cbba1dc41b457cc30e70f3cb37a4c27e1366c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cd31d2096b9730946adaa51f977e1548247c6ee1dcea3d85f423ed812c9f9638bd19444ea735ffbb7de70c2c0f7c405c2d75c1cab848284b77f14a5ca4d0bd254fd33690e313d7ec275d50ae117fd393ca6f5ab4120e88a2ec5c54d46aeebc6020dce5c16ddc1415d2f9fa616851bf0cb292db29bb7d8eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1368f09583adf879c3a5902dafd9b9e042d239a46a8e95bce1f52ea31c8a5734680a59df48466402a0e1b25f715931d740026fa220db04107b35ff3abccb6a030053110fa3f5cd86eab7940824bbfab2431ce96b367b32abc7ec90bcbe760ade62c211ed689f6a0c709873ea659c5f5fe8282744845b96a9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c0b3ec00f92c0364e4185b6d11697915476bab24320b32c6fe587dafdaf7b2300defb1cfc52962004489a15f0a9a3e15729f1149c0c6297f8f67ac1fe202266dd266bc66ddeaa52501fc234bb1b42cfbe54013e785622cb344ab4bd550f905fc8348f3fd99fba6525e1cee14e36dbf8b325939bb3135f3f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14dc411c33db6ab7ef5f4556f8157492ed2e6ce9a16931a0fa61bfef7bd32d4f9cdb7d3a9752ad571ce2788390491fb2012580bc89959c748aaa3e7f2b466952aa6de32e1422372cdd2fb0961aab186d26058b5ed3c96a91b43213a0d285be6ce956c22d6175a05f01ac1e06ee8f2c2cbcf5577a171599cc1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac390e3c2163e4c5da3a5ba8278316ba12876cfed1219d08caaae4dda6056d56728d644bc2abf9119080bb7442afa119b966db3b8d384400a2e94e59c173a07467254ffc6ebb841dc56064a3959702c20ae5b9c42967e3ef0ee6f1ce3573e01971083ae415da05d054e95beee3b11a928f97d9217505b59d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf837bbd4310493f1bc03947ec2a59cac55bc7982ad8b4121b6437eb873efac8eb87394f0f1363f35fb103e1902c48c4ada32088f9658241d36be8efc264c1a9969ed7cd4d7c5c5ac1b1e55eabdd56007218782134db7a8d0dae39f16931186a8abfd85c6cbfc9c3b0a4ec72b5636c3453b5305cc0e90a5e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9007c8bf42b98d5d7b4a0edd6336c97803e864ff0d15419a8ffc4df5fbcaa5ce72ae3b33da317d0fbd23a67e089763e311d6ff43cae0819ec5fee066bf0faf59c48507076d2fe672b6e7c4ebb2b395d057548c8fa991a30cf80dbba133cd10ff4746a0d9f70f37c3e980c9e61c2345b1a20f5568bfda451;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f97af5873541aa9dffe6a7a4a27f312ad3141aeb124e9e6f01b75fc77dcf38ef7a57100dc8c964380638d33c5db6ac0d25095feb227f3146379adc2e6fb19c9f283b8ab8ed346b4f472892dd82f9f8ecba874105b229161918c366e4f29295889de51c2ed209d239f9c7d5af909762e128779bede43458d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9d1f2f8ee402243520607f420fc8962a06e2f478e3d64668ab70ae2ef2c2078fc44cfda28437a2a5ca270e343f01992343ec672dd4ff68bd65de7802228aba53941184fff376e08368259479e503ffa8b65befdad951ad9e57ca678b3b9c844d743b83bbcc613c34fa093ccdbe400eb6b24d99c191d7ad8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58f39c0535387a83b8dd8611e924cedd44ae744dd3f6912d5d8700da6d4fc7f1b5d167658e47bde64a2730e80027d21245d9f931077969f401650a722a8b5770a1c7f84b311da492329a3a3030fed4435614ff0b2cde85dfb3a5bbaac1b7dc9ad3b41691db8cedd4e8fe27f5ff8d182e1f98a19c9faea669;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb627356d35f3b1470623338c113cc638318e16f89e2d0d56d7ea1bd7c74caca1aec2303aa07f7a8d7c573790837da554b9ab6e18fac190f34cd84f3dc80190f8578b9fe5bdd71f6bb8b7053453cb717421a0a9bc80714404a980ea47be7132045b5d7dfb6d16cc8760126f871ca2c0e9c78f12f338b81d4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7b61df682fee2dfe459268b7860692bc1dcd1d98a0460eefc7f33390cf0d454a621a96dd53203761d0977a5aa7a4bd42450e1f765f1ee093309f0a3a3e0ad09e5527df89b6a02a3dcc75f8cda469aa1191d5e153efa32805c06bf51a63a9183392294e56a5089ce1405537d2d934ada26c3626828ce44eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf23f673e15a6a4a226a2b9be6f4f2bae8b7fe71f0a7710f1bb182e35b684f97b78fa5fb367000e07c9bb4f5734f94eaffb25d7b070873492f87efbdea8bb9996d18c2763c43f650013fb559e1c31df86f992bdaaf2efc31452ff662e049fd2ba728a5f403abdd99a4ca801f042345102af432e02a521525;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de21eb0e6544afb08a38f11e23d2f24efb4250cbde02da46adb14bc822d36c7366f47a227449d7dbd313c29dc39ca7e7437952badba158701eea8460b1cd00d79730e22f5c2ff51ff60781b4d47d9f7269ebbf07da922b39c2b30c47f4f0b4e95ff4d57ba7bb6942942fa6bc05c91b681d2ca88e9052e29d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b6e558fe6304ddd8ef8d43d353ecac9a1233e1473216ab62eada0475eb80b839d9bbcac9e5eead2370188c5c34b537c3e634abb1b5a9188b9036ec68f2e1b3d5affdf314a956afa501fac5deaa7f54e49b7a0384617a90c799487d11228810eb1efb42b89fa908731259ca5728bd950da713bffdd134fb4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haba9520641e10c9cb96149c3545a29b87f17bf46617fb2d5f23727c4b4ea137ce2ca2d718e2f45e341e5978542af5e7edc0699eb401baf13c7dab073bf7c96aa20c8aa462f1c71cb7c42f58beb5cb462a34381d08b1fd9ad3a6bc8b2df852ceb63a822df176b0473638274c34fd89eb29151360596db29aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a6728928b205200d19f283f482f3a14d285c5a2243c3ecefbc7cf941c2d17a9b89675401ce3203dfc6af5cc3f469ebbc15f13cdcb003018aca78ab6778b569c18a900c4b7648727ad0d2da8c1ac8a3ae4bd0258ec901925fb51737559062d6d4c308a11872d0beef2ac39b109a5112c23ea14b0078fcf6bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2361be3fe84132b1fa864e6a523e24b5a016298a77468ac1c16ba1b721c640e922d394e950a8638d30d75c4fba169e1b3f754d6449e18f6aa827f31c0c3115508f629403d6497bb7bc5a49d4a47e67c5ea3eec8375beaebba305367b7a74c7ef5fce017b91fcafa2887270b124d99c555892fc6435bb4dab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c4215334d06edca93d2c9c5630e8d71bd70fca549c1ce1b5c55fee0a89137882e854db2c9304739e298a3cf706dc353a654a48cbe64ee44037edfd686f5653ebe8ba245cc820b7264abcde7f5aeaa0e252fdf97d825ed535edd740c33e0e7288777dac8bf521b96a14ea2ec452e6b3178fe6aab5c3f3c97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61c025e30f56dbea1e625d5e31e37a66d83678084f19a33303159d411f764cd82dacc4a8fae35ab6c47635904ef82c2ab8b81d918b400dcfc14f6630b774fcb916ec3162eef08f81a1246e5141fd1af72df906fc3225c2a8af7f9478ae59a0c2ddff38a3037b9167be2c65bda531aa10bfdda821ea12b392;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b0892f5f9a1cdd633890644b38babc941280e0f670a5ee20705164693dbb91366960820d784862297a5bcfc603525111bdd48092c9f642da8ecccd3616178c6a30ab464945451fc473c990d3a9afb8742e5fef0dd310cc9303a310375064585284a2563c18ca700735db3ed201f1998d0357fd248da133f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a060216ad1cd69685d0371767344cfd1c4b8884afab22c18a3bfacaf213455cb0885c650d2472f64d16b144e2c00f4d7e9a248444e0129fc836daf7c6dba8aa420fc1120b4a7a929465537f3a1f2ddf2e4f31d6ad921ba5eab0c23f8f62b99a9e927653b0d50110eb0a79e84c144cb0a2cba272eabbb3b12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5a3aa30c0fea20cc8ee063fa92c353d9b4135ae204c053c1b33ed5b02206ff6a581d11e11f2a45d7c64398685b787fb920c0a3d28e7c17133d5eb6455b5f37b06a39dcd2e96358dd527c537ad1edae3f1806b0c6b46f8da61a2ef8c07db66211d8b790fe88bdc519d43e2b639cfb7878446f68347af2e1d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcaa5587f7ff1f8f5303fe67dac786236a1f5ae142ce7cc3f69edf361c8b0da7d275a7d50fef9b116e659041eb584a3511c3970276bcfa4cc593d76acda51b211a84ad1835b8f408eea42d84d95828145f091bafa237fde0cb93ce77719db22989cfaf2c6807529238593e118470923580be8c7e6bd29448;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96a2d2b6f5145cbc4367c44a6c4c8d996a22b279dba51a46bbe7f54db589dfe99a19d8b7580329df6824f5397fdec76b7c6c37dbd208c0af9d22f1d55c2e18b555b0ccbb5ebdd5d7aaac0fe6656e297dd0791bc7d551b78f57dd9114e6673588b643602839d90c892fd8b908abe576d3614c34a71a1adaf7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h622ddc8ae7fc4fe897fe2bcd7a6e2837b86bc72832a765d7d52c021a6271984a0658968b90cfba623a32e32a50b522edb0bc2f783b0df067e981ad424c7484e32eea844615cc280748a4b5c765b518c6234ad6efdcab0e0245475197f3084425ef8bff409404210da158b9ec0e83dcfb781c312bd10e2b13;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd0fed6a7e7b6a27c252ad6098686a1f1827b99973154ee887de73ee19eac4e182d1f44a04053eda7ff2e5d46b0ddf122d77e0715c2962ba385619f7e277fe1b768fef6368433b4dd5dcb9a04b40c02d0a48e8fff5ec4b076ee2ec66fd17ab91cade772339ae4208bce7a39e6ad22e2615d7ef7d32dd96f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9a24ba2e18aa10ab29fad7f638ac7ed65e28d81bbd5bf78365ab09139f501e0475383f8a88270a98444d36823653a88d30cd0b4454ff04851c4b415b8f29e1bd3539572f18d7f85b289f62d0d56d1e6eea86f728fd1759f6e6a521e64b63933da61cb2c7f1e5acfc6c7490a353be005c32f47141e4c339d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e0bd79af5339f1257dfe896c476adcd940d779639a876524d0291ec33ca3dc96a1cba7a0c7dad5431fd6b8d888d87e4768cff122eb890e575da829e64b77e23f6778ace45ddce948904745373c6f28b5831aa21f8adae5165b0a01e23cddc9d7516de6d93356e88418249a3df0058c92abd6550b84990f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a3e6738054ea9642d9fc10ca127cc543660b18184a20678543517d45ac0d55b9de465baa5a041564e6542767cd25a2ae0cd016753bc7315fde3b7b0aba384fe6d3414420701bb7c0f660b081f588f31e19831225b136ef296b29342112d3193905561fe8cf00ec7071dcf09f784aa9b796d68d85a7a88dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c25a1421b1ea8c379105da0110b67aebc9f73ff5e4dad52cdb96586503a8146068442207d36b6564c923f09230604c1d84ee31a460e6710c1e4c38080a2924baf202849c7316de4b1a781eef1655b03b51b622184086d35ad0ab4b7ab45f37d20568135a1c10b69b2820fb41fff3da42e07b6d8a798818d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115429e6b205314609175ecd41863e85b92a3ea0b093a29ad44cd87dc676ea29dd44796fb3f5ca1dd423f879347957318bcffc720691e02fc622e2bd99ee19ae2b46c6b79389fde58b9900724aac9bb9740e6276fb778333e8b7b7086b46e41034c3615afdf8e0f7d2f9798880f7ba549f84799a8bfa153fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151ddaf211a95c810e38c0a85f6c6ddf03ffbc07afbca0030463973b0186eb6d2f7f6a57c8e53fbd9bf083b44de580bef07a78e5c1ef3522aeef62dfe0167069a99e98310524534e67e90729de9e3ceb3f072f2487b1536eba1046f0ace0fc82ad3b0bf9bad00f92937fe744c3c4d39146b79646fd7504068;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1504f230191ee79b674929957cb160fb19c0bcbb6ebbbd8b6102331f0dc182a4a7982396525ab0786b4f7a2bb7b8f19acad209f0d9881d6a77eea3f83fd1d751d6af90a84f81163560850bd284b7ede755a0afb8f060923344db010083abd55f71e2ec7886ca201afeac207f4bd36934273b6770e119839b7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17bc0d8d03dc69bd0d45fd148973b2b92c7d14c69f803bd9878c228cad2355110cb88f73ae45789efb2b0d2e06409df6918384aa8b1af44b584caca6595036c0bcbb7e039b7d852c5993349cd26021646b2b1634a583cb07328817461331723115862e8363234e165b0e742daacee40fd4f453b63df60e53a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d611b0f22a02cff933b20cd480fa6972308d8988195d50cafe6f2c4f9a1b93522d560d7d8ebeecdb5d4efa4b8facaf5557f93ba6c7ecb75419ead74fb3df0a38cf5719c836a9c7cad823783a0e035770dd1aab9b7fbc24a68571ad6e5f3744bc0b169b4cf6f7130a32c6d61f6103522663224bb4daff436;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48e024f87b3adc5a8f54f4e64400f41d672d16fb14328ad19badf82755370e9b5b10f04c3f7cb40e0e4d28d68c6239a15f2ce1efeb1c9db09d381a91cf0f890b0a608cf45819fcb474fd69c48e67ea1fe0ed0102fbc19810bbd44c5b80227813de1ec29cb39257659c84fe60eb69940c21b4283fe454bd85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd772eb00edf2340bcc00e54367dc8e8ebd87d53a19b517eee7120a2cb0491a3365d51f7ef46c06c99c3a9985e78c8330c2408ae2623168c7e8f9157b6d1c96efc80de6fcac291ecda0e765072898600aa732f7b6c4f4e434270a0ccef9a6d013fccc38111931261d9f54b82a3362db03a08561791bddfda6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18529a700294ff9856b11ae9eaa14c7d5c2c79a1b4deb7738d3e178fdafe576008d5e607edb66b74a517aaa3f5e848dc2d2632631b92bb6c153ed606d028c094191cc5a6067b995cd8f68b9741590b032aae6ba2208470caa8a056428ec5d9c3d437f4f014fafafc384bff92c0f74c3a408ba344a06da217b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61a93012620e790aa22977d4e30b7b3c1061a1b243db3ad5466b7b13e8167cc84966784982a6f4ae212b2fb3e015d150fa4d5f7be301876ec705198323363a02d1be300c60c4d82c436b3010970c8620e6edd16c9cdf5d10e289d80953f852f3c6bb50c2a52cbe6efc6026e344ab0d3acf106a9168d1b5f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f30e31b5b2054caa3b25b2141ef44181f6cc23a3a8df0ef6da54f4bf533557ff3d117699430e346981cb214b5d6ee5d3f2adce0eaf6a5e76453f6258ae8e8ea73af6526462b7ecf0b119eeec51b67812295b2f91f3c37a27c80b75341034c959b087386ea5c37ad7ed2b0be25747449193d3a2e90995d8b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85e289ac7c4ee7c6606bb36671c4c39cf15fb215ac9c3fd7deb0e52ed34b1cc03995c7e48758013bc29c076671f4a1cb714cde9dc5e8c4cea985a8a2ac66e791feab431b047ec45d334a1f1ced5a8ef6dd5c80ff185fafca1490d9b27ba1abd4758c17802c2af9e127294a8ccbda87636ecf89109ec79677;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e9528e81ee17f20f5eb9851476b7195c76aea5074f100fae59fcf9c5ed0d29f4defdfee0de7c2a23ab5cb079c20b229ca3516decafa5c543c5e0517934b4c76735eb6219b16c152cd7a21f46f5e4f5228cb04af9598033509812b4931ec2ee6e64ea739d44d2e4597cf6f3afb98a275dd51d91c62d6aa4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha0cf56c514f6ecd0bdf5a1c020cb4be4a4f5710d835d293d3da9809723d224124e78036d0aceb423d3641d4e3953299d0a2fbc368be2d86ffa01f6fc3e9a93bc5f60b7779f852f858e1d66a55512eb6a12f5bdcf3c8964bf1481e7e92843149a0d3c070e33350aae4b10e646d363b653bfafc9a5bdd046b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4c7f84d8716f4f8ff48e445ce22d50883b98417adaae9895efb9334a33cc2084ff30236d24683e87478841b775a59d04c5ab281eb4bed3ca9cef5b9545acfcc8e460c81258f0e689e836a7a223f52cb8146bf78a0d4b68202903da5fdfd8cd13f2cf1d1b91fb3bb42d6b8fe0931d5c59220719b49852034;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hecfddc5ed753408949dec72d98e9eff96cd1f73d8bde3e1ef804a0f1e15bdd829253a9ac7149bb6643db9b1ca1ac6d0edbda5d75074c4177b92f474cc4584ec61b5e3c47c4b045dbe6a4249bee2ed60698210d0ba5a1efd480b69c76756703f8cf51f0e41b6c9d54eaada039b81f7bd047354781ee486ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133c5c2bf1bef799124033cf4337f9de024078460a0e22a260546b221a7d3fb5a32e49bf580abbd4f9450157806cf5420417d4563900705707af97b2d1aa7a95499b185a420e1f61c79deff18d32bcc352b9e0eab24a42b413e2a13a6fe866b2686b61ba7c90006b63698b1cbd61544d7855aecb69dd9feff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef26fb398cfdc1d71731c6a3e3caf5c7a2ac03fb559cedc922ad893d0c8d905db5672754f4bfb437980ca69337969cc2f0cd043dfab001d30235b2b264f1ccada16425b60baf586c88aeb7efc278d680ff6c546a4dda612c2f18cba54b01a9ea9f2ec91bc1283eef5060843a4835e4634440938d5910334b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e68901f20b341f0250c6bba3e9630c40cff11d6c43081c309f528dd4428ec96af2adad367aa04380681d1181ed4bf51ea1fbc2bcf8a969845ce7f974c7bc91d9d9708585e60113a32c4555f06c5f5844d8e1814df0f1bbe749b3bfcd2e41cab5c0b7ee2d587e7441f44fc8ee8bf54410b6928dd46d6f9c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13738a6e29e166c8703e84e2ee1a48353c66c96d18c296ae4dc449b506e8c32f6d3d4fbae1a9e7b742396427d5fb74f35d1579fa4f05eb5a7ff8e946d8ea6a2b6ca8a1adb04d7d677a1d3609f807416369d8a33ec8db243e6baf7e229aa05aed994f71f86e7cc2f92ffa244d52712e14f3c6bd0cf4c75073a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f0bf7936e2a4fe7d34547832aa60c722ec549c2eae817fe2b5916cd23032a7da5f35e5288b1311f0e0a47f934766e3acb17c47fa458afb6bff3b97e62778b425ddd50dc71401e7f5a6ba73e6ece79c30c855821e322abc60f10ffa65f06753c10bba42b05076eaef17ce3142f101fbbcb8887d5d8a1f99d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104e529929c564e7225da3f0ebb6ebd92a8cd98deeba7cb48d4508f4f45a1173df505abd9b939a1aa50261934c2bd98369788200146aef0bb0bb48cd3c228d6866462c492e3263668a1f9ccd681603bc8d1cf40d42562f6e5c7c61da050dd7d2d93bd5804010ed1ede4bc8cc65f5e43ce87a44ac8f45d3945;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d9a2e8f3bc211821b84b4b804f994938131473691741beb81a527c63f5d458f8c1cc208cddaa5a4200d4ec8ea6a3c342b2223f56cb2fe6cfd024cce8ecb97ee9d1ea14748b1fe8a94e10bcfce21fdc0dabbb9c4b971b066caa404bffdc14e99f152414298e0bafc0c5e86692b4573d41f0efe2163d6370f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103b28e7f68e0527389d2289ae8b72b25b2506e177de343dddc31d275647fbae23ed78d216db29b0d4ef89612da07eb86d3f6f4e73a6d032087648c8b0306c58cf33e2d6d22ca1239be592969eb4da8728e94502221f2bc3e9e19d68acbc3d976190680af223a42923200d980677d449f3f7e9359fe6d4f4d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa44c6ca2111baeddc097e96417748e4c6fa3a984735eb639271325522636ba7b6aa8ca56ae8dd1d4b1ab6bc3df6c5a465ff3c8e2fd96be4b63a1e5e9b27d8967d6a3c6d2c6ebfe759c66c45397c65cb5e6fe9bc49fcbe8d39d39dc9803df3056cff5971ab21d11b4c875fb19dd7590aed189260a1a187e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h887c68b2df30a2af873ce848e5761fdb1142257e9c21ded5467c43483ec8346bf53cb6c0988f474d7ca8f3dc6ab474c99d88b06e87e8232388e069562a373c134d246c45e817daafea7aa579a45779dee6e7d0d26ace549f8aaeeadbcf9de85cf0a319c3f9cfd70be48afa0f6871c530b31b50baa7e0bd80;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c86514c8390058c9b81f09f955293dcf94c599022b113e5c7a567601a86a33440ba3af46ae014a476d065a4c1f1a910a5883e0811b922d931a8d9fc0e06e217ca5dd5b162a2618fb6996f04c57fd1c48b41a4d8f328589081968246beb1fb6b81e821d19bd83abf28f6b1e173150ab7026f78c2ef2ea0c5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae394ba096373938cf88cb642f56d8eee1636a62273c31b46c4c87447e03aa307fbbfdb6f151de787a491d248de0bbcd66ea7a01e7eec28dfffb13d8653a5e28d0e54b7cb87caeee98b64a8710cabdbc84b278a8968b530aff335354e51630443621ef2227fbd9a1814d74c12c3a58fbff371a353d330548;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c90f6289e70118e625025a520ffcfff2996e4fbf0a95616fb730399cc7b380881bd11af636dab4df78faf9fd69e0f022a7c282af0472425dc1853b8524afa59503caf02b7c795c2db6abe7606f6d34941dd143696384eb02215017db494bf1fa3b673639f3ba19d7973245c6061a0a4faffcff38e49cd382;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c1960da8aa709182be9b2b5188342ebe0800096cf5fd9c1840bddf57844d6710928af30c85228720643fef7e1337faa0b617e76a95a2eee3fd9db4a36b03953dc49acc655898d4d35874e763fc7a267ba78ff20bb0ae750ce5dbfae212370564feb8462cb08fb58fc74fc7032af7de7425d065bcf2b00b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56500f3cd3e27ab48047d2eba914d7ed92232d13a7ecc5126ee641cc59e127b60919a4ece19f47e04f007eb4ea1c141a5dcaa3e37dc2242c8c8a3ae4055d58804f637418e8959d13704189b9c3e797a8d60571fb5af5721eff59b852862895ee1993e9a7b83d7bbec07eaa89a9d0c30e6a3c3caa113db8c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6fdb49650cfaaeb55e454bc9f155b2f0586aa0b28e1cb238bf7b9a8d944fc7e532c2580f068439a2909f943c057501cf3d5fdc9b506f94092d23f395ab6e054752719a970333112be4c86ea8a0e315d86efd8306ffd55d1b12e848d8e127d10c38fe538ff9dd0f01f342dc6db7e0d1e02f11f9b59107c69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34ac6c2e5ef4538301b260fad08793cb724c93b0f9d910a41f0f091b6feb11b92db25bdff6fcda1bcf3d6dcc045cb641d82f9e96e8e87a5d01e92e072bacd68db12eeeb708bdb2ed28a6c9ba873f32bb321ff7470f8d57550235b14932d8d6cf577887cc1ce8a51d3c9ab61aa93fc489c5681d9a1651c882;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d24bf55049a8fe3de745840a37d230172b9058c52dfc2cc849b1ffbb4d2075ade39a6ae4e1e32120b2a81544c1d6026c4657d2d52d0cfe18c3d3e8b3a16bd17e69785db931706ea1360d3cb2bc66e8456ad6bded1de1d7e508bbe4de3d3c202ab91f757925ae768755af7af776ecb6de2579543a43d3f2c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f22ca0fdb73a7a8dd0a9fa20b89eb3e184cc093c2b54326041e1cb0fc42b7262e6dbcf35d30a526045686e78e6fead3ffca91f652162163bf698b90a5e32394e4a46a221979608e066db276f07b214b8963fa0484912a3b0a15578528bfd004139f065c3cadfa2bdd166a970a3a9a3ab7602c0f1465754;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38e9fc3af017eced333c62262ad3c8289ebc2fe7f63d1f3893e52ab8beeda09bf5e452b747f386e29845aa7a22c793b2fbf389909dc840b9cbd1437810d7fd24f3ce75e6ee2daf287e009c8b912142dd528d873282ec1114887379081758da6ea88e804736182104f1fd4c2fb9dececced8225a23003e3e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0d407a8bd40f691d1f62389126612d12a45975bf0aef073131f3667d184e629d01b77244cb587269ebadc55b90798fdd99986e38d99ff11e60d752630741098bc69ebbbfe223824309a8704029bd868a5828e13292997349b097f7a209e57cbd92443b98cb1b60bcf0cf4ac517e8f86db98affe59d8e0d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a457ac5ce7219234db6cf857d01180fabd19ed42548a3031305aa884d87ea61f3e340c212abdd295836190cb9e8f10949e1382ae0bfc743ad2f1120ec0a89baec3e103defe1cf09bcc8099e29564fbe2fc641a671b1d909a58d2b5fd19e31cd48f9ddebd1c9a2c4880bb2e4f1e57c5cb5877b5e4f0d3572;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e67c58cab49c078a47ccf2ed3fa49e029ea0777ac685e48fc2e11cbd7447162cdae90bbfe41b06ee86a3c6f9d5289df17776797f34ff2c2317967dfb26294c7dc70a12744d6540018c8ddf34d505c232b13208b9a3574650062dd16779355fbaf7b32b2945ff60350a5ee69c9cd5254d7b6d042f5561be9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a51ea6217b1d266a05fc194956afd15d768d7a3a27fdf83096a7dde12c0aaae3c8a5e31aa09f9d2737076ffa5d5111c94311918eba75136efb4cea3e43d5faa548c28213e218d5f8ec838469a304cf9f166f7a7cdb82e021b0d3e34ebf14b91b240ff6fc2c53c09e491c5191d989df9e93fbadc0d51ecce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2684f095d98d66d522d44b5338d117bc73aaf2b9fa758ae4ac73442dfac25de2361d2bb72b09f235c9c66803b35210610ecec58a1e24a3567d2b41a4d7db59ba90f76b66dd79d3e702802594d2f1a87ff655f3de8070f6ca92ed6c602a9d5bf162d4d84dd78223286acab6a6eea7b6cb9e17c63927e8d88;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114da3f873ee154c396c3a7c81f549a9152010156d7fff2ea29ae4e6ee4409c24026607cf1fcd7fa0d0d288b7d47184a3b735455179c5132b7022ffa8ff4febdeccc721dd29a488ab9a057f75b723a7c4cabb07a07337caf193fb786321c44047bc6f3824664dc3d3f1b76e7b28dac61295f21ea7e4950abe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc26c43957872562bf55e2c34571b813d9672337be5a9361ab13c51060a1724453bdf314cafa9023bfb701bc68e7b1cf474d7cf3bae180b87d0450d0c14a1472c33ac05b1b975fbda4d89f34955dac02c4ba3fb4c6d9442046da51bfdd44e1d7684f83f1c1efede71499ce5e6911cb56524f6918e65bbf7a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a00f697046ad2c0aa35718f2ac42787185a9c22e5c87303e068a2f1cd08f19af707765cd005418511905380db5e2b82cb0206e6592f7c0c90469dfd419884d03f4bdafde8a19dc4570c1160c86c06634b79460210b624dddc3d5d3b6f28c2c70149b98f38146023118f28ab93c69358aee99c34a178433;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f60bd90d65d1d3a97f3e5a118cddf5712d90562890849841bda60f6042fb22a9b83c4ef19ee9885d582b6fcac38a86bdf20a16a7e0228ba83e2b59832f59739a0903c5ae2a05d217fcbbbbd0cd7a269cdd6f05a34193569826313f76b80a7498d427a0ac6e9ae5e2eeb99193c8ddc2ea092b004add1915a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17835c11e895aa8aff3c6b0d6893aa8f3fffe1d454ccc47695949948c0f96d9ef79f9ed23f84324552b14407368a90a7ec3d2dd558241be598623198af4b19f96fc9e1c0c359eb02d4c8aee2ce3b56e87094e6e666145664b73b1e615a3630f0874acbfae1c9088140d4a56c35ac8c10edf5c35e90c8163f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ae4e1eaf4dfc752b5b7e3b989ea8a9b95c6517ab5bf8eb92406e8040d35cad0335320bfda95f8585de1d3eabe08161a4a30f9febd1ce61789d6d68f94a0156b1512d7e433616bede1495e3c1e5fd8709642553f48600f215cf2abc072bb88ef8ea37d61ac2fe4065a94fbfc3b9f684d899df2c4ceca53ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38ccaa811f6783e566253b0a76bacdf0a504d5e8c5da186f36806096aa2128c170ce7e4c3b692e2fb4a59df9a554b4cf976db6a14dc6228852397ea5d1bc91ddfa2703561b36106258fcc0a4391238746a37d325066975037882be6595b5c32d6194847435e674466c5e921a0e7c12febfe11cb4531158e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c4f81315e3f95fde7a2c9175b57203beb04fb5224fad5479bd48677996f689553037b1a10780c96fa310881ede03f0072bac08856f6ffdae02beba58ab4e39afb2ae49e3035802b24a21975c774f0f3898c954f365e426945584038130cfcf7f1627cef53d32e373b165b5d994760dc2687c0e33055f685;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15943c1e231e8a9847d7f30e11eebfd36d22a83ad12ef0ab00b981de34ff8f53f16baea732e41aee9938cfb9ecdf0a7093256e8b5588fc42717cef68d071610a323723b302df158868eb98f01d07de707c091ce653e74f004aaba6331458ddf445ac16cf64ca7e99bebf5fdc6a9434539287dd834ce2f21fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e9d72b3474b2ba4cd80580bff88772032b1fe7d34d82ceecfa14d635235f7467360a180b300ebe4ceea8da24d43a1d34cb72292cdb9a4c8c3b136c17bbd402528ef4ee55254182ef072d83c53c3df2c165a45f1ad0766b58e16258ffade553f6781e07ed074bc19ab34d36e23cfd4aebedcd93efc816a2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e014bf9215627c213d41b0024e651986d973f9301450a61bb285f01e599cc30b404b44daec2902ab5473cdfa29ca6e166dae98f55acd134ab7e7ae720fea31d8991e84f3889f25354a9cea52fe5257751299db29bb9a3869748e420c37edb2dd2f2676749e8bfe9081e659df1e8610cfed59f5724312671;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180b8663dbe7044692eb5ece58fabe4a44748dfffe49e2a10efa06cfbeb4cd64eb8b240e0b10ac084645066dc556b3f397e6ab3a78e9808dc6c7bde7deea9ad96d9ebbec6b85f609f283b21f4ca0b8331e85f232672700b7b14481393691433142c50fb94561c23168695d38dce2e8a7950ac4683adf8ace8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h743840b0a6bfbd2cf34fbdc8c49931f2f06418e61512d5da975bc08a80351ab5b1938f27451cc3b9cd0e5f5ac99ef1f221d7342fb7e85211634795d0c68ae3cf3deaded39daf9ec3926433ee724085da947cfcc9d072fcd2d5e276f7b6cc9b273411a084044f9768657d3f8e62059d43f5dff9244e7deb76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ed789abf9177ecc78516da84a58cfe09d0658426d70b23265dc0a4c71e3c2145d6186b9cbf565979994667dc1b4808158a6a4f490c945e7b6023a5a1d78de12a856c8428e4592dd935836c8c2686a6fe8d543cccefd1d8eeef5903ce8dfd54dd8c01e61fbf107e58148513b701e2dc18b87d0de325f84e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1264ddb96f5dc507ae7be3a9da3465073dbe15faa23efdf893ce0cbb6320ace471c2479848372715fb4968a8dab8a5ea715473b73290fe2d4e6d843a47250db9887269de52a1363f652713a93980136b1585e7debf5fbddf28d5a24fc424906ca8b4b4569757989e5438696cfcdd76859e7e0976a11195d04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0fac4f87c446acd6b897695decd90bbb4d9d2ce8b4474a81895a29b74d44fc7379a62775a8b13edf298c4daf8717ba8d9e5824bb51fadae1e17d6efbaf5bee7ffce4bfbdef8400610a19b2c771362d32ad572ac4e64c7659813197878fd768f60913c1e13cd7ba7afce4d748a3e37a94f1fa19a66f0d089;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3371bbef44ba37a0e69367bcb20ef5db194b223b65dbf74674e36b7e2e36f4598851f9b27cddaea333d889eb9c442bed1b0b1e3b115906c1c798510cb5926272da76b17e2a99d99786e41581f96abd853d46bc940415cfeb424fed8a10ce8583c770f0841e4586faace320b5fade380da82b227eae6d3fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3616fa62f8af3e90ac96a819b51ee09e021d44062cd5489d178ff2ed11fc291eeb98575ebc2527ab1f096472a04b409b05a23b5157248949af9fa2bdb8a2149c96422cc87cff65375ef893bbc0dcfd8c594deeb2c049d94e3a8a86ceb6d81c411ca315b84d6f79e60b30c186add9ed3d9f8d4fa36558d202;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10668a3f88f5ce015c523b397e06ba133a1eb0c8ea2b05296517723ff022fd2059ef930f2e8d0959f080c34b82775ddb56ed30afedc577a484e9326d0f1317c8b767b2cc5356af02d422d8b989867566dbd0da87f872dd994ee3efc3272364df93f8270ee464f3bf3b36b165347dfa27076307cee32d36b37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e5d7787f17d0bfed158fc61c751c7315ad6878f3e36e36fc9cd92dd2a597e33b2019fa2ccc43370fc6ae707d766a303055b174ffe8cfb45a1c6f4eff89d70ef3f8bd215b34969e00046057031e90775d3d8fcfc802686008e3b35035e7cd16fe29e8ad4028a3f78cb78bef1cd26049ec3d93f0755808062;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123ca5bf1047a57347e7f7272d903ff7c53faed1000103c02ff9f1624f52f59f6383d6ddf9f4dec05299967206cedccff6ff8351c54b19d4ef36e30ced2e51422c0cf299a00568f093427def64813b0648a473d933b8e0d587721f8ab94b521dd8dcd872a3621dfb69389951103f97bbe4920657f132d4e00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b1134b2e4dccee77cb52bb00816242cb4c8dc3257ab077df2e11b25983419937996399ec08b32080c41e0581a9cd038025d155831f1f070c9656041e30799aab307a060658bd898f5443eacde750090a45a7cc5aebb0ab281bec5685e215eb5e7c02f9c71c304bf52983383dbb82b2896018a9784eb4356;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dfef97d9b9dccc62b1a9002f37a37832e57a2bb4772354b3af82283ea5b85e838fbac987f465cde01869438dedc4ac49f0e8c0ad741cd72c60fe9e4e12fd6b330941c4f11ce27fc50352216ae1189fee4b51d4d796e46265e09f12947b644cf26cd2d10865ad175c5548997a924b0ad62cfbcc4615dd9d39;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a21fb21b2310f79b815d9abcbad8f934f6df6aa965f36b4e9f8ca35ce7bd86796eb117cfd2356b6c13721f6339492587d6d0706b0f33f8acd58f79fc29a6ab72fc9a6eab6bd4567e04a108cc4c8465d5bc1f06b0a57a3dfc918f105c8826f2b752a6eaa896e8d7a7569c8ba9e92d255eb9b44b6cc7c3d268;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18005d4586fcd38eebf2e5074646486daef24abb44fa8999bac32b1950d5f5720556057572c86273074d9c1686639308aa809b3bc028ba3594a9a46c415193e5c7083b88cc54f79340bb8753812aeacb1aadfd67ff1b815239ea1352baee55667fe926b423f177012c80446060703d134b8d1f394f38cea8c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6aea9dfcc9e5823c29b37b8ca3451f371f992cb776f637962d417d8db794141ed4250a6600972767ae933b3fbc340c397027001754a66e5cc17d67ced69a5d63c7fe8d27039ac69bcc6d60032f93c383859a4e16690afa316714bdf124b69142c480ffd1ac39596aa842812a643ae4730e685ba4e0c9d21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137bea5fe92b5b67d112c45023a455dd92cb39bc50a5aa419cec41a6872cfddb88d58206fe31ba2db0468e28ebf5061a33a25883ac2f6d47bc65906e50d529855383aea34b9beab522e94b5a18caaed971c55e2af469f573283916903ff1cbd3c9af1cf0e4b7f273d56deeb390087b254bad9bb8bb3bc11e8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3b03fb6bd31eec1ff46d43a9e94c71805f092f41e19cecbb54acddd8b0eee490b4fecb7e8199e7e8d5e3d60e51fceae9f1e04903684b0c73a8a9342b04979ee570e43a0f0b85f6fd5cca57541cc9fca43a569ae6526016352134f22a139c9b98cf3aec7227f01774137e10cb0a34728a436659a11d0bd6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1906b6210e49815fc2e5787638d51f3afb5168990122dc9937df5f95229590a87b8f5a27ca4df901738644d61a486e56ed08041ed46a2d89cb70191f4888dc96f2d1b484a73aa81a3728a4536a8b8c523830091d7453edbfd9fbee2e02e7a6e665046d77e143abf2edf33ddfc57091516444e01434e5ae051;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27bb07f61cceffbad604b7cc9a54d6f5eb8f20f5303fee0439a6e826bd9bbcb8d2932b7fe3814a664133c2f9adb405afeb6233bad3c9b7c173f7b36b33208914d786ff062c28ab862cc2fe896b96aec572f618e77dae2ed64bfee6d6e07de2cbd9542d09d2b7b0612188f6f97c5c95395b044b3235be1f37;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4d9664d18d1e0c8421a5498f177833f84d5c8cb75e0d147fd23bbe881f651417b28700b3305bdf23ec38dedab395f502e776386ec8b39eb6e20bea04d2873f436f9c12bbe4e19e5878aff0c5af09d6fef02383c03dc15b303292377c04c9917ccf0aa0f3c4d64ad9b4d2feec378ccff15047966e0a9df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb645bcb9919a9e259e3dcc00dcb61bf514fb06123aa2fc07528623e006734edae761a93957982183c920200515394035c7d706465943ff022e8b365464695ddb338cad251125d61918e898cc0946f36a199e84d0c01db172969a94db119d270a1df6a8e5116112c6af5e9bb08cb0c6e41c744e8d07877b7c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63c4e0c8fa168e5f742f3d32a55ee6e7ead167829b68f7053556b2ddbaf220159079aa19c5155957715345095d8ceec1ab2b0bef087805e86b66dcc8ec6a9a9e4f44a166c6ddcf226629edbdddb8d69f521fb4d14d60712a0258b3a6c3ef7ddbac21d76f8727f920256c3e342d41b7ae1fc41a1132e13761;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcce9720e95a0df4b718edd0b593f7d13a67f98fe15aaadd62c9cbbd6819e825258628f851dc4de912e4ea29ff991b6a72554ec8d330aab1a248ba122032348108aca5679e2fc3f767deab7992947081dfca9903c984f95d2d2f7f04d6992b2581d358c423c2a58879e9e940a6707fe4bbe70ff7f3155fff3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb9fccd8755a3ad8172597cb7733bc349c96b76fb7594180b5b23f64beb41e30c3592b158c590f5d473e63d9ce202a26ecba5759296f5d109b095c2fa2e9db2d8e3962623ff1cb219900c00d80fcc7631f97185de03c106de2ccba6f43a992fc5856a1635c6f8ac7c46e4f99339c8d375ec98e37f3eee872;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5f81e82dd71c1dcaec95316f5f7449a9e3061938c18293c11e99a90fff7529f42e4cda4404e79819b1331d7352ab17e1e04858b4646ba84cc7e1db5982f28605f6981e0e6e3aadcede4de1e3483ab64aa5ccabdfcece30313dd5cc55606758021d7159ebca28bda8f2fae270286cbf945bef8aade824145;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1212ccf1ee22831ca1f31678eff9a23d087652031ad0f610423ba79975cdc82b090a2cff5f0709fa7a9826bcde5a2a6c8b17c78f4467898353439c6614529af79a873591c978a6b08fc395aa95c5e109f0006953370556347522cc424cac4e4d11ab233dc2353e9bb184b110450b3d456d4f3311a77da0464;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha26a38b379120442b1a5c74a8676b8234eba0c3e987a8927dd2f0111340cd3db770588924970c013177f1d55fc222f5412ea9046088132957030e3a291ce96a1fc8095c7d6257b62c3e3717a5813efe1f270875ccaa49c96a171bbb20e0033edbfa98592e821f634c8592e7c9efb4db27b0db53a48bc469b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdfcd2813ca4fea30fef92852b190b6e172420ff816c7fb21b0234089f0ea8752889cfbfb74f6d576572b72a7df6a2277aa09ff5f8631464d7ead7be547165f95f79ddedc4d8ae977abe62adfa5f7b8eecb6edb1acd006c27dbc8071664c299e15399c1b53383e907b9ba6ccb27da55fb2869e07f896341a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab62cd19f21cda7236706f713c8f80dd3431ce9cbc306b32d3da655619141eda063759948bc92172dbc7a5bbddcb59f746a1ad89a07bd09d79884d4de8d355827752d9391cd58c0b5e8b8473bdc9a64c22fd067be83145f2d8fda65ae14c98f0ef3d43552bf44d4a35f974ee1a425cd621a139829afd1f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3573e04132b86558de7dfc8c0cd4274787fc4e8adabb3a24821f140297e143eea07ca52672b5a16118cf8e31a55d56a7428e73dc475962d3d943ff6b288fda4d94e92b336e98ac2b2710f556398d869319b94b60850ddb16026d6a273607a95040017d9ebfba9d3ad3b7d6888e1ad94aa3d57d720d1d0d00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169e863433b734e3f32f9af3685d071c6ade7ea7a210485d028d3af94ad0393b2d2c93ecb6795fa4e6b6a0a0f27a67f80d8a08f80bea49aeca1506d451cd00589b1ec52455d7d85b42e000b9275c412565f1accce8b811b677f382e5a99b438403cc758c2411f4927a4d92d06c664bd7726532abab40e1cb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bbdb1c0aa317ef1a7226e11280a9cd90c94e9dd7d1758ea7b4404eeac093828de24ceb49607606ffaa27f1ed990e982e91aa14655164a90406ea4f4fa5059746a45a11eb9049c5af1db9054e97711f76cc48463415dff3a213c27d3e2b3666c5c709b4760441c7278968651dfdcf3d39ae0cd4c8fcc7ab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had23cd03804359927e43ed00a14a9b093ad231725e3e1679a716a292fbeb2fd6972360fbd8cbed8051e68b496679712c7d8afcfe713df21d71c224bf4d30143ffa1b772efeb7f242f4bbc465abb11def17d1b71b130bb38f1a933f3aa8758210312251102485a1ea764e7d2dbe0a4ad10f4ef04f477452df;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d0b9a0bd5356307c46f17a15be89d3a31922c36c03759b136b91a7029b4289040a44fb3f501b180ae1f51432d80e249377063d0020fc95ec20dcfb7803ec738731687b09ceee0af0f15f43a84839fd5e75829723fafd80fb8e945f69875b98697f1d3c0e34de3faf48d3b0e8b7d7e128220286010c45248;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3971987e18bca5a9e48a53189d7ef97a1761b3d34184ae6e0a1117f43b9d8e42d8d27f6da12bc8808c01878297f0fda43da48586423f5c860b50ba8e97b24321cea9e7e39cfaa1c071ac539434ea3e9c7f3342754711d85b0149f408ca965bc61e6c500ac2953909f92cedf25708dbc31879652236b7e486;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e8aa7b4c40a20df7b34e4229cc17f5837bd2c91546707c998f5751caf9e85e50856d23af4da741f242e15ba99d06de7530b8cd79843954254defcfeb5200d72bc1a4aefa89270f01e5ce4563b8b390c16a05e06b91205cd35df2876f82c9ae28ecd8eb746456841f0c18fd931a5003dc0294042736df332;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2621df418f10800e06723127b4dbd88bbac07351e33e69890369b887e32bd58550085fa9cd261c21bef0b2515dfca79f64fb7997b6ffe911ba74b87fbc93d76f0b019b401d86b7bb8fce703e20e81f641ffde60238bcd7c1192668862d5c5ec63f25327e9abb79ddbb3d93702fd09bd4be90cefa202dd678;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc97378f7e4737f60d0d80267b0f8973a6a277ab5015a4c55496a2dd2bb49ae1df0a826a016efcade93867a08f132cced063e1853f3edabbf87896d8aa58a96b58c9f1d1c03014e89a7c739a248d725f60f2651fce4e7c1fe74f8830c27d6e38e36fc355cc4a7a0ac99c1cf0a1cb90687ef9c456d9ae31699;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f95d039e29ce56d650de90d9ad03040081879d8f7cf3601fc3a7650c3879975fc327e9e98afbaeb6181bb81fee1651bd42cb0289f1a31d1f2306071abe30fafab08ca6da442dfbaa47b224a37d6a978395d2d21bf3f1486ce8bb5f0ddc7250f90e0f3533abd1010208ad5ea39753fdb8d45e5d9acbd4c1a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f5d109009c7f5754f28e22b9f7c3dd5d8d8c7e6882f713821689f559199567fe772e82b6e4845ed1237bc9d7075c6fa984095ae3e58e2a3fd9216f9320459f925f1f2010961acffeff94a049c65f48564e8dfaa66916663ef3b9a90edbcc5ae46183322a1daa7d910055d3d30567d98dc89de73d7f14263;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd79f7197f8014d2f28390b889b459dacefbe437bdda957368275718046728d3cf28dc65906c3eda61e748b04b02cbbdbd1e78d21901746707324adacdb7f45eb07ea030411ed48890322d8c6d0c179a075c965aa6cd71bb7f156a08074a7dfa2614efb4f98420614c23ebba842dedbf8b050d9a9d49d957;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h174d76eb1353f46c42c4bbafc0a91a58bb762756fa4488dd5efa351c35d545a84b10a7181e500cf0459517281dae5c3d944ab25287a713833dceb65a70a181f6618d6c147e8872e7639370f682f55c2bb14d828e4bcb956023687bf87a3b8058ae5855ffc07ea40d5db4bd3dca8593d67bb1a773fbe588dc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h619dbe8bff06935e52ed85a6e2a2281ea3c0c16be9b41e7ced5107d2b3d292e794d936ee9b811efd842651f1dbb40622921995c7dd9676ac4c708c82196cd7ebab714890e388678a1772aee61db439386e0572f4196c4fa968ff9977f2c1189db7c3c28b2e3af5dded3b39c831e37fed42a786cab5f43eff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aca619422d803e767c4c495962283b8443c116b4df960af9e7ffad9648b52d5c88345887207994e51b91e58367e7fb7dc79f57fe112cdb794b39362c2f5eddea74e8fa6702bcda518eb667b395da91008d9bd731a8e7f0404c90f4eab17598c645b1dca4333b3d23f70e0cf8b38ee9531608d9542ae0c9ef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1feafde03f30dd1a19464c2376d4754ceecbccd9b06a000fb0e3116c39bfc6c06ef79fd3170277aff719ac985761235ab96e8f44b104786937f5246fe221421b44fb69c00ad235a617ded95567b8cf6ff89992c8a793b17494536856b6ffc1b2ade52cf40b45115228c66421c488c806b6f1340cdbc9297ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79d2d93b049ba3ac6c9c359dbe943a4092ff898320df58b5563b114a90cab5c0cd79f77e7a512a9166c6a832cde8579b197f57393b3b4e85ebed19cb1b2e95bfcc97b337fea24adcb23ff2aeeb4101a728dda393afcd7e8c433a7e7d136d0dee44397b54dcc157b245bc1384dd40cfc0ea8dbe7ff9f685c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb81eda01f24a077d5f54152b5c4bc80c5bcd06f00ac09aa38d5f70a3f19f32123fa97b78130ef2b7e13d211b6e9dd256ebc93e5cb8b4d128126de0e33ad25529c6c5db34accd82c62977850b554f04a38b78955edc0653854ba0c8e6b68e1c5ae8a96c0c86873995753570a97887791241af036adb438cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139b040f2ca7db6cb90b07024e36b3ff93fc23ec6c23e33828051e362ffb0eb9b9ef04adaa17ded0a5391143e659737eda5aa848e2443051ea3462c2154b79aa1bf29bf4cc838f4ee09d461824932d71c8a037802cd4590edaab991a4a8e5e55245aed66a547d0fd7966d1b3aa1b52be455cce80878ad4030;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b318e4307465ca2f641f90342141aff8351bc700b6635321cad4b1cb32e407042a33eefa66a6a4f4069d2d5fa5fe1f1e9d3abcf91b7d54c47ef09ea4d79d3394d3874149da6f0fb1a0820f66f5b6916963a2a8723a992e8ae67c1bac9a095d1415dba53c229e926ca46189a0b0a2205c6a092dfafa1d318;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h174710dd282ff9d935ffae6bbd14e349d228492b27129df93a691925f23683d9186a49de677ef6dc70c522290ead99e214fafcf27ff482e202e98780f813a0921499aa10deff85e8c1cd38fc0d1864bfa7a4489cf24eb693dc26d5d659ac9b2e918762f8ad67ccdd791ce0fb0819397dc864b479f56aff667;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0efe82bac81d75725f09126ee466e262c71bd5e4056d9ded9988b78b1e6eba7c6fea5f95629fcca722b55611731df4373ac73f76128b6e2a1794baf0ef08642ed6cf54b75f808454abed0f53bc49878a8ae52ec44bd45797f16bf7b8b7c48d14713ced58920179ff55fd1ff19205fea13778b51f3c9918f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h412fd1bb22bdd2a699774f617e1a2cc0f6708a8af553428be0e46dc9a24accfa5e056a1794be6e33192f9620899f3c7e326ff68783401783a9714be7c1949ace85978e4526c1a39a3cf8e22886d9ab4cd51eb3c9f4f712103fda88f0aea0d98ba786b4b7567ac2ba337199bbcfbf98fb5312f0134e83548c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h687603f1104799f58b7fc3048c677fc5633d98c645888959351e11eab4c66530e0c42a293a18da0aead9b421cbce191d6c1cfde7902548e90f028c2e98a63471d1c04a2a379f4ee7363586344e5769c6619f388fbeaba98028c376aaf6366ddcd19aef39a6cfe84b4e3cc43dfe72ab777ee44d47dfdeef67;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f2a43039de2b80c941c1a3f1b81236e98df3016ae6c737eb497f58082219f6009d89a4c14d27d0aa568f1299a2e1bbb6aeb7340a492b02dd6ef1496ed9821db2cf1d23dfd49496f9e56d0d7a0cbea9ece1efa19dd070d88946854c267b3fde696ee32c90c71dc938aec36725e4d6641d9f2051ebc7be453;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1677c46e6b12fba989ef045f3a586b4c0278311bed71519524827a63a0b98170369edf33821914b18da4e5023d8ce407509564913984ce0893dc1a2cf692947255b344917bbacc933dc10e225a7bc5ba3cde748d583ea6cda3a2a3360ff54ef94bc557e84c889c40f2694bec7bd711e3861080843371b9310;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb44ed08ff4fba54b7e85f270873536449c847b0d987a39326ae1dc9c4f5565f70a30e475f28b94a69dcd955c09a17dadbe0a5440b0f3469aa42d07cddcf27078b118291c95df1d8ecb908865e77be612dd3a6404ae96a8cb2a06886b77b06b519abe41048c58a385ef6babb6ed23f7ee6c2d0f9d42556c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94736a083cfb611b564d7c03d3a3db911a5f3fdda2d4e413a5e6537668bfa6ef716d2326e498be20a52d64079b2a03d68450130fc5590969e08319556cc4a310de1b7428e58ada704e82e40bf9d2c28eed8aa8bc4c458c796c0d918acc180f3f32a319cf1f4d52d2cd815d58c860a40c0effe49ef6fd3e14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2086daac2164163ab4e29cf745db5f491f756adf1e45428bc17549f39a02fa3192c46e282ba3458bd333c4913ec0350e18ccd2a8977e06e9c430022db3af368f04bee0b678eaef33b5a33d4388ea7d35bebc27beb666c9ea59676333642144ff29cc655e4549047cd85bde6cc682d848b6992f4aabe513f8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175610704b0aa8f42ec3b44474ccd4c69bbaa499d3108126863e1ce4aea718edc141d18325a3fdb12d1af1700566e8cf47ffb674897ee2c74c1242fdde038054732bf8434cd4c4b3035c0dc333a757e5922cec2798c94aa9568bce4d1dfe4c2a681747c785294dbcf3805a95b1e9582acf6985c75c80b2dba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf83b09d43feee2b01be7c03b02ea0d9bcb4ece799bccb15f53b31ce7d5ee9a3c0091b4a9e573ee91cedbce6e69cbd9a137cd6ff70f79bf42b89c5ae95a375870805f6b3ba70638c8ec7647ead9168173f3bacace15664771b11229043fcd326131adf4fa1435e22fd1b227fad6927e27f6a5af3d2b79132;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e6b68d22fa459c4f1a5aef01cb0585bab2e8a222755efd7b3e811a6b1bc71b0769167abacf5a3f75332b16f5bc7b615e9ab4c48491aadc0087683ad2597f5044ba89904185c3490c9e778351b90ce1657e0ca59a13d34a0927fcd27552317f4303407f1302906a30a9dad2b8cd50ec1a562c700fbc907dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aca52e1b91ed21d2ee1ee4e07b0639f9448bf5641dc94e488d4c4b142c4b9158d6c9473e59a230a70c9a4e7e93fc0f3deb6e2f9c7a49f220b26fea4c0c04b182db3f2c68c6b34f87eff4fdadeb739f93766f13e76911adb7b27cc474edb49dacf7c0aa172d81a97ffbc3c2846b092ef7dffdca0e9069f46b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f83a2edfc9aae6a81cfe0fa014a11f1e54f9c1761294d721901bae2acb376c0687b10ae7f861d6eb1e49dc183ef1d12cfc80b6f01a505ff749be0d8d44e7fe49b591a39b525463c34f21b2070cc286b24ae2bd7aff679f1c966a6e617b59d7adda1a416cf800a4477eb6718e468adc0019a39ab477484b95;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da8246b9abdefc9d430dca7148a05864fa1169a52f0d143cf0fbd39a79091d3eeb670ac113b3f9483dd8b5660803ddf584e408327d9e7ffe694ddbb2545423098408991952e4383b87cacb56bdbb7d263ed94d5cdae77e6024ac05fe69365e4275a30dcb754fd79c980e24c440b5f599c8c50a96e5aba5e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1020084d6c34bca570023151a958d885437cbb23aae80b27f7f26e367f755f30aa080d9db1175e8717208a5bf9a08ab521b82af2ba809189d585c68a5c7da1fc23aa6dd926793af8acd496c9131c01ec93ac4d50174994bbb0c7301719186dc375ac1693382a37007ae84d079aca7e89fb6218c46e4310c6e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b8e8f442dc4bc5e62b88d1b015d511bf8cda67fc8ccd054ac9987c4c2a7946e3ff357e187c16705903ca948cc6a8d4bdd2338b207726a9f1469cffc454652fb8616117ac8df14827683ce7d2633d3fadf35499b0da7f2d54e95303adc8fb4f385e249dc3ae019b18f714581689cead7ffcef9ee45d88e98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2907c81e7a1783739f8944e26e4979e6ee697a1ebf6b1f14d4b0bfd6adefbc9abd0d4c89a9316a002f813ce7176df1f700c7adb8e69553f03356e4ca1b722888ae396110babff986545b70244cea947648d746078beabecf339f4d0f7177983441ecf05acd35950057378d96566dcfd2691b5e5eed85ba6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9e48540f0110d38c227f0ee204e90b9e45787685ba0960f50c7fe5f4e05068154859b8e59fd6e510a31c8e15154adc89c2363996ef170b4095ecde089f1eb09d54d3578df2245c5ced64487b0d90466beecabcd5df8ecf840acd01fadd6197a4d6b55e206f33ba23a7a38e86f67e4d59bb6042e3d762f96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b35bd08df56fc99f2fa9eb7e864b094b13c4cc440b76d5d66d5cb9325809751d28c517232f585aa4fddaaad2ad509dc3ce96a8ec12d96e785a96ba7e2d905d052a20fdaca2e19b36adf500092c26890355f21e28b153f4603a4a007f10136c600b87a2800fb2d6afcd34f354749b34a4acf169c4a5c8e85;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181ba992803ff6e376d8cc8f22c0f2829d87b3cd1cf31757b609ad26145e923337aeebe80bc1e61449a736581c1cd0fca50dd298a734c1d212a2769cdda388e46a3f9cc67e26cb6b820921dbe031b9092566882c993f1601cb2fcd4f89bed668724d8d45c55a5a53e065d272742e572b7d02508bdc03e92c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf44ba2cbf93efec93b44701d8de42ae720215f71b440b240dce74886708de32541e7ed0ce6dd687de749227f57c74447ca7ad3be573ad0e95235f86092e870a831de84924bc3d73f1b401a160c5de2fc0008d24bba163474ad6c3007e64fa540c6f7f21e62601cb93b264afc319cc172f95c7784f04481e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15546a80fabdcc62202500efe1b91ff3a7fd8d89312a58f14b547cf43f257cf7c3f20e2ec3ca67f0943f5cc8da51850f9950fa76b99f16bbed56c7a24203d9a8c33813c98baba3c5f918f9c09188371706a2352e684ff5682458385bd308741f87a3a335d592d8e2e3024bd86e4ca0d71d63dbf46223f6990;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5b931c0136b20cfddce3a1f45fc40a0d7e781edcb37862fff57936caba9412c495fb39cd846339ec6a7191e9bb2b02b29cbeea5bbe701414fb20df22634457cad95918775042648ef4b436223b71fe5837db2f65cc9d4f506b868cf7c7269bdb8848838f458e047180f53f3d7cf1a126a64cf4088ce3c65;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ed2c172de61d752105389bdfb5748d34f6684b190948105ab9233314a629e453bc4f46edaac01e8e9a2194d756023391ae6ffd6f4ea6666bb23c31b82a2af9dbc9bfc4067f1215ac80bb1148638d1291504b8e8a7ca24ca0d1786010616eec37b2c37fefe8e0d22ee4d1885857f36353df2c9e8f8046c10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1569cf117e1e9f3dda1d3665c52e9456eb6724f370269069e42de5ec45a68e0ffd111b3a08cb0f1575a04d51b752e7f8bb374681ebed8a1ef78cad2487fa745535964a122170e950d645dd0503eade57e6a8fff8cf6ddc3915e9ce7409a3517b8517a524544c8a2bc358e5647ee1fa9f2929e748fc4c54b3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he195c2a7e4507e3b9a04c0d7685394a881b4103e01401d07558c0a544e018f474a4969a7cdea739db67bcbdb0d37744525d4d96eea3dde915d60377342999d9cf863c309b7987906cf99ca1944a26abf8a9d2fed082004721199ec0bb95ac8bbfbaa000b992f313244adef1c1862821c4f9dbb81c39dcdb5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4eb8b2ed9fb394cd2132d16f87e8e43d8af9d6c85527f1d0f8b4efa3ad0158c63be8d56895819560a0b4eeb563a9fcff249cbaa0e94559da9857c540d63452706ae56b84c3617ff222aecc9e8dedb0c432fcd1178ca657d5f3a032a4e79b1fb102c3d428c0ab90a1548cb852b79200fe21c71de678ee2f9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4d015fade859240fbd00b7ea10bf9244e6b9fa6ee3d2d2103ea418e5df9461aa2e58c65eae6d4f3a213957b85c16c42d94d50958438858691d12b0fac05000c12275271318c71d6cff1695fde021954f1339fa9741c9c56b62d7d0907ed65fd983ca06ed050c7544a8754687dbb424124c4355cb1617191;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c2cec7ed06b8bfc167309ac7dce7fdb08500dcd1a46002c7c2ec303716bbbf7ef414cb62cca1a9af66b489d9f3dd0538adf9b054fd3277e40271d41961c2aa743ff6e29eb45d746405f00a89dea89795655ea5039172098b001a70ed0ee3ffc708afb153024dd2f66b45fb301d7d21a15d657a8e16f1902;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187f8e2b8c6bf85af302089d61a6255cc80e91abda07af4f458a6c547d72b919eb42957c2aa1ce9f688c3aaef13299201f6357ac6ef561bd711ac4f1bf971c700d3f21e649016e26c88a28ffc0137f51661a60109b0c8524e06af52b3d08147fa0bd5c81e3b785a3e3118c484d3b03af651fb2a41bb8a9b51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fda2f102e46900ddd4f84c65fbda080db3de2a881831bcf7210ecd512df660062acf1fabba48c6db8c0f39930cbeb0d2fbf30db383495637fe22af0e14acce4b7273c4d693b79d970b79c4302efe3f68e42b7055a21c35746bffa6d48736a6be55f1a2459d1fa8a9c6d024a3ad2f0f6287881e1a31e8e238;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1497dd6e9f44dd215a2792c387162169026eaa123f26cb4299a8216597570caee40aea7d0c97d298e15870d0fbd30f4eb206efe5b67c6d40ea3e01de06a12d69cdf36741fe01d8a189f84c455b96aa33a3c291382a79b56b25b808b5bfe7ed8a4bac3836ea6dd88794cf870c10898b8271a83bc7c0263366c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1451e17edde58c07449fe47da3fcf7c28f26176a923d9a3d9a4ab4f4002168b3fb35b6cbab788602e6e2cc7ea7ec63a4ea19824d4920b65216229b8f85af2fd3c20c81a0b1357ae3b2afac88d6ca21945dd9bd7cd6bc21467aa1d43820cd9f041f46882ae8488c75d814110df6162749045e52313879e04cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a6cdaf61b47bb7230700ae6ca7c7e2cefae9d84b58096b97d62461c299f4a3290c225fa00bda1ff1963fe9fd7f89e064afed85d4bfa8b5cbe5c8bccf58436e74fd54eb9a5013f8fb4774eb83c31deb09846e26158f142b23d7576c83eec0aeee2ca6f338fe27ded0dc32384135e3b06447677aa04ba2a2e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1629b953f540934bd8ad1d192217e4f13158f7599cba44fdd379ab406f060a0d461c959e4c5c7f96c7e96887eb43b9cc409cb92f13d4a36b2d1746d7233bf90438574ccfba28d2d785368bae95f8f5736183e98b6a48be138f2202da450c313698ec6a3bd197c10a0fb7bab89bb9f5c7a53bfb6b00a6d3d5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb7882c71862f2ef155f2898a4987085933e50252cc037f4dfab8fccaa0f11a242d8b61475d0e00f7f56e08c6a4932be7850739bc084b7af44ff56ea2f1c0398f04176c8b12df2423414e33a8ec0c65e49cf446236c4673e44c202df4b82a562fd74f2c29f047d6750ee622de3008c7a24793b138f71fa92;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e650a19829dac6f404e9e51fbbd35361c61f9c8d6de1d0c4d339a1a508ea0080328fee2a67853c3b66700ef235246545e5680d9cdcc9980ea0e3bd49ad85182611542139dc33b8e3ca769f004e312b0dd00940d983c6beef9c3faaeeb3e8ca156e7ca5ba1e1be28cc08b4b15f45cca1cd91601f18b3698e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h311779c7b7d9948a15f88a70c2a9413e4911751c04c467d57475c79519f97d3f3a2e171d916f201a0967273aa3958a83769add0d950132325c54269c7346d9440ba9694147acfcda199e1633b65de5377a8354daee08c4412d54940a314f331f71a5435ea247318c0275317b42776c33691ba2fe01c5017f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d79fa54bc7288c388e2de481074de3fa5c34363a1c9e8ff7408f8174d0094c788a30a1dc9f42383a84f27f21a53e7db2670e1ec267e6745a774662ed685de1e0a2776fe7cf14f1926be4584957e3dd75b1ba5129080c0a87c742b1fb90e27690e33be821082a70c56fee90af507aec591044a9119ac9c07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h822bc707659741d6f7cbf9b66fa90392db08a7094eba710728aecc38b81711eebc75f4610936c69643fe498be17d83c1bf9afeb018b5c793bdca84967573cc2a10d559d7b79507f26da15e707027ec48d252b96fb31e957e58e79aaaff7b84f022e24e7e7ce42d38a998d232e21f3cfc2a8f6090a425a608;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4cc41117bee99253c842039bb90332e0a8812f28597789952e97438c58d8c31d5ce117208b90fa75fbcb5434e944c37f1fdce525bbd4e9e51c1307fdab9dd761552626f9984fc4421da55f81a45ef9ca608e089232a965cb5ae1ea885938801fb5071fec28d826665f0881a29a4adb7ee9bbf1292bec153;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7088bb8ed16ffbea06198769e863e7a216b0c524d87843631c092ad9c1cbf83c02faf3156e0f77673bfa79753856f44308d56af1e1fabca01591de62e1c64ddb831d5586ecc9106ddb8a65f03caa5d20587135bba44fa9499f650813932217ed5cc2582ae8106d96ad6ff881a1101a013a650b210610c7a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6ea435f4dbd18c54eacf485ce7df0ddcd1d54ef4877b31d3f1eeb3a8c49a29cb9a7ac6ffcae7d36d159e46fb299c41588e804f76f0cec39134fbca6d42cccaa957fc938fae8d2f17c792bbf5144977b5541d06466af87eb0042569af1c46c2ed7096afcd00aa86629f020fe73da63cfaad03b28a7c1060f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5af5446f8de80cc18131dd197f983fbe3fd95c92af02fe786c5e6db5365939c2a7518087bc7b63d67542992733ab40fd333317f62ee90a8f1c65ad43250f92e55cbb75a4aeaecf9e1b5754a3eb1a9f94694fae7c726c57825ffc64fabd20878b39c652f80f1b1a977d8dee1af19ab9e2ccb61a293c23f48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haad1f5a11961d9e882b1dc2843055812eedee8708bf9d2846fb6feb7ec48c27f10644c8c1f56f73a3211c82b83d778f7b08ff0d8cac5c73e9e91cfdec87f4bc4bcfb0969fbdd7c1c02fbe91e0936bbbd3eaa4a70e0dbfa684485162a86c5c1f4223916077ae31a1cdb4237954f2405a77433ec617296528c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63de05be9812f132c1a88dd130518385993ad79a1563c8e35bc8eb10a6d3675c0d1c541d496e5ebb050cec74a4b38e2bdc27eb6acde6a22e102e3481c65dbee4565b94bb07b6ac84716e87786004f47413f99587e947849a9cced6ba201447050128449750d474abee050b56a7be2603c90625b649b7c260;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8be5bcac3ab1899899b926774403dc933192476d69e814d57f44a8be32c0474caf8b2c9f80c7dcd7511316894d58bf6cb4515149c100d09a0a0d5265e83d3ebd3784b72e4308ddc69c47306193914998acf44f1c3c09d5c2dd5f1fafa5d69fe189038df9495ff556e229bbf62f51dcaebe72d838b1ca643;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac857efac1f5749a89dc0022532c197e7708d141da5c888a9f3cbc1e200d1eb46104de3a09152d25b88c8140306c0dae1aec18391a3bb1a60ff5b0e8ce8be497ab4c5b2a95a32d37468d5d9fe6be95c5c5af297e6dca50216aa5b74638cf46c1d119da6d1daf1e1b9baf14d83ef0e43663f4595fbf099a6a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f63e60a851a9860f8a6fad73a07dbb4cc0ea415636c35f5bdf773772c426d424ff25ad6cb19115c7351c414cb022c29c720639272563e777fa93d814c3bd4bc0bccdbe09298dee5d7bd89e1ee933c468465df7a5526177911c6a61d57d6630e7caaab9676700fa9b4e2e483bb5a57f5448f0e256b2fbc9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13749dc2904e31624b54fba1100a7764b911d7c105800437f7c379bae43947e0f12acff471ac761875462ea4fb1cb2cc916aa67752ccb888e090108f7427a3ee01282e72f39dfbad1d29d53fa156d9265f066997d2d4bd4408631ca3de1e364b0f216f18a31290dc25b57cf200511f966114c71325740b4ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17054754c0011b6e2e1a026b96734a14037d6e287af8e5f16993f2f4e2958cf3c48ba165fbc0100fcd84f08470221549fc306aa3cb0c278614d0d9d73515128a87b0e83dda312378e3579dff1e5a97f672bd509d35d8c1f5e9be908c57e0e7ab6328892a74992ad3b65e93b6551734073bb4e9336d5ab579e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b113a70cce2a6b115a027b7eba2ebc2a8c1b8b1e27f86465ba98b979bf969dcbc2da11cae01470db4af1e465e106dbeec41032e769c01c3dbcccb59d497dd75181020074fdf252a5554b125594692cc0f62016bcce8b88c7b2ba2846477ffbdeb745e08243205e4b2c1769b64c0620f44c8a20e2f05b390;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13dffb179b6d358486ebdb4d7b1e19e34f1222b4ccf568cebd7656aa2d32a443ffc78746d0963da96c2d3ac61271dfdf1df612321d86e39007eb6ba7e9f1527858744d9be4cd2aa3f7cca0a41faafee7ce520e7c03212560826a4df5f0183f46dfa21fa5fa434921c483ef55911b0c537264ca389ba33182d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17689aa3ed9c85edd1f0d95f3fd715f9054d8c57bfa7e80a7e4d3e574bbdb21fc1e809e3e022e5df64500a458bc20fee7f8dd364defa628b0e96389ea3815e184b82b244a1d11779599eda8572f01f78db3b3bb50513456c1bfc1ec84ceeb5bc2859b8327eaa01526915adb5d0084229c423faa22505f5663;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h273bba7e24cc3fa476543406b2c08838b32caf4f73040b067902039e19197a642d297e501496163c43158e675953d95c1d607b13b86330ba2651ec60ef4316bd6230517aa33cdc59b8714cdfcbed584b5c950d04927aca500800aaf5a3f424a9e69c889d9935048a296e0f5d2acf09edeb64e306221e4542;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19311d7f1f5ed6ab8d86b8990e1aa417b0475f2039688d7302e54ba3c247dcdb1ffcfb5eddcc3c1a6f40b6559bad803f7456dbf193996e710a4b1d5e15652c3e89b6497b23f2690b6f169152c6a7b09bcfd5d16f0e4fb2c2a26774354db17e1f29a9a2be8bb4983be1991bc2e40ffd3c803c62ac9c7ef07bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afb9e596e11237ddc32fe996371a81ebfd7ea601d15e2a4d87d9776eb04a232146c66b4cfebfd831035ccdd7c0d4fc0abe359183948a97f807ae87d5165162925b87155651017d3a1447b9449e665e910a77969d8209e9fbcf7187b2f29176f504699420441db30cece6b86dd6e0a82e45ede05c9f9cd083;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f77b967a349621361678481e37ab921b4a41da19a5e5d7c4a0f3efde240bf6d5a6615b8e227f928923583c4fb29fb7a00b9c9c8dd0a552476bd85789f58a8291bb090d581379c2621848495c12a8adeba47c40e0b669fae71db61da33c207b50cd2f9f23f59fb7a0467aab8a94da8d00c31a8871624d1f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121a68ec109007a35750c97dc7241e5723c692dcb3ca0e1dd4433deb8eaeb7a94ced9118f930b2b95693c40a067ae4ebf1d5e8b10be122cdc6284fae9b91a9962a3665ad0925946db4118d8e704f063bae8f6280d66de1ac995fa33c472b4c4089edaa1776d4c4b73edf9488f882daffd2470e03b35b25907;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12535f10d0c3c301a22da67104bea341b9cb584aa9250d6b49cc4604f8be64a79c4c83fb06667b0db0686db833fcbcdf19b9e4ced0614689bfa19a2aa326034e8bab944349bfcf8c104a39540c1ff8155653f413f096424020bf6c13c14f9c59b9dc071edc855b3a8cd1b6d0ba752c30f9da7ec7b57333026;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47f652dd64df55c6b44d02391d5c0084329bca2c6c4facbffd8876aba3abb735b8295cab88678a165abcb253328716e290100362fc1dc9abf48f6f66826d4c75a8d6bc98263b6501ae9535625410907498c91e228824ce206bdafac3ffa8a94d4a16c5d51dc25ed2d7a995afc4e9b2eefefc26192e7063c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18bc8644af2ee4c30a735b301abb41a25cce98e7f5b44b8f4a7382837fde10f614225d94b7cb3217553c7fce0ae90136a93c272eb21f158dad1729846fbc1814e03438d118e4c53357ac2fef4a3a35cdbe4f5bf1c0a86cdd183394859d3079a20b3007de5612f339d52aad559c055729b3635c5f37fcfd47d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he77b83f82139877c1cf5dcc467697d88db958b0870b51fe2bb55b042add14c35af7750b21f29fe2b19315ad7c7f1aaa2f751d0588b9cb91c2ed6187f39e08cadb6ed7bb159dfdbb09393832974a44aebeb9a15a881399d636c9f3e18b91fe1a4811933e1f0abafe6b0fe554b11b30a26033f5540a3947aef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2a5eb2084e32f0afdcfe02887c9dc8acdab16278205beeadbfe17081dfd7bbef259c50067d8e3cd4d2ea9deb8bb98099f7d53ac5bb48e2194660ff0749983102c5ab7815cfee95e325c30bff8f003a451d8e15d619592f62a6a361cbfb779397f158224b4a71cfe03731244d9999b69205c516936a2c977;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14eccc50ba29fc76f52f369f97c6392dbd9ce07ee6fa5890ab896000d57eb9ea4a68690e2227556413f9d456f2b0969119477ff97a3d7e7296e524646ab1d078dd2e6d8edaeb10d285f959ded01e8f452b802353bfa17d2d891cf97c57f33e6201cd720b29458bfbe577b451597bc90f2e499a4d1224d851e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f5b81505cf148fea7cac68d6eec1befdd979688151799f9e443ebb0307026159f9ad53da4165ed60b8da87bfc36433e61017b278b71cb7dcbbdef164b582428185c19e0ebb6d5b10bed87877d982eaf67220759ae7e7f7c958f111007037daf86950bb2afed529a4eec17d04f0f027323df3c15fb5ae8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hecd1e3c41e9d5955108074ab450159f7ca195cb0593fd7244bdc16154b177003d29914bba01cdefddb5af48bb2bf53c5fd5d8d45a8c82672c88b8e9d301c62fc4ea9feac13a3aece6b07a994760814d2ffef64dccf6abb0712022e3e0e8e1d1bb7712ea6043cb5113af2b26544c83cc7249fe58ae120590d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa3f71b42ed16c9f96e4753262d49c5bb6cc97fa2d3103c67d56168eb9990c053305548d2a82064278c592838e6d18255b0853ba22e362b7bf1f2c933c7029f76c366e201da769840c3bb74ffcb2ba402e80b1b90d2c502324b8ec57eeb8f303b3e5807b2cb7528b0165b9441ef9b11653bc389d1ad879f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a07983368a16b8269e04e585eb92eec0c313f29cc10bbc0ed422dfa148e113923edc5501aaa0300d8c2767b27fc6b7dce4ad659bf4c883e6ad53fbef724b900f56440efdf72f942c10a2720f4431c5525c59bd87c3a5b5e6e0090124c266f6d65ddc064623b6625b8f3b93030c24aa90f276cd8a0dbf899d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45d3017ae60995ab018d654ba38e6cd5d642e19ffb1c862a8ca1842716324a9adb27203e4a2fba78fae875aca2cde7860f697268dc0a4ff7e94069d45f5da08340205150c480214a6f7ed3b49f8db04d1304f8cbe36ad44df974663dce9e5758bcf9fc35772e3243205ec0f4d942b1a808b0076d88523b8c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9e96c9a709427f65f673abed149c7522de00e6742d9eec7a9b911511ecd7c4a526c6f4f002dc00e41fb8bc737d403cac5936e47da8119f1708085cc515a30184ff985f38d19baf1a77b043eb020d13803b803fd98c96f0051bd03f9fda274f8ed6e08ebef4721ee0dba8f9efa247a0bba19eb8a42e1d290;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80983c0245acfe02c2d226ff3468aa2c2f4d76656f9d87940d706a7bfa85245f36027f14da82df3c792de12acedaa934d8341c8bdfb4b8983ff86e1b4bcd74d95e7aee1b505e5c93f679f6de27d48c59c8b25ab27e36dd838780688d9948939d1cfdfa42026499e0eda1d994b6650451a729245cc1cd4abe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h81bc6ac1cbddb17acd11a58cf39edf09a96f3bc68ed3b44a231b4a7d9c255eb3179f0d920c24eedd1f4c4a89ff1045605e800a99d808f30dc49965d5dfe870d128e27a28735f103ed20d3458454486d8090330fbaa0338d8663bdf424efb65c01d17c76fca85b0c803c0457a092c5481b971c7ca9efdc729;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3eb07dd6ca88daea0e8464c699b8fc9c7866f826ab82483f1c3d4f291778fb97974895282fe1a2942b0841540367875935af850a83e0d85fa9ea5f17dfcd11e478da27166f509039b84be20a03f15cae91fc251998d3d0df30d63b70e0878252b1c47769ad91d72d9b02d998496128cd39dd3d70bdce3d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5fdfe878becac1e8b7649684edfa2fad8ccd9a2f409522a1d96e0280b352db8493a9047d974298b51299718245076d0f551076b694e81bd914fffbdc51516ada250b38c93ed15605c78edca9519d751afaf927fc49e80e53750ffe49732b7c1a79efe487c682846a1f41bf746906ccd2f199840a967a41d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha47f1fb28bdbe07f186abfe64d458673269221ef23ee27bfe251767571f42f0402db257b53dcfdc22e2e78be1801c0f205f4194d7ef6ef5c2ee0b0ed36bfb0efd2386ab2925a0b1081f7b85fc51a0a651a6222fdb7247d84b3673b79ad3b66cbd53c823c03b6e632530b6aae7eb2bcd64cca3de7ed13a6ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7deaca4e8dc5a2f1a0bca207aa0104b902dac2d526ee5705c93a5d44b82219ac491bb1159c99c1996965a98c3575bb8e363c6a9ae7d37912a8ee56b68d4b44059e6f3474343c79bacece2ec3a14b376bb2ec57f43d39b801c8dcc14b60e87c878518c9a6ad47f33c3e6f83c5491888bfcfc87d82bb7d9cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18146613888b182dd965766cce0d7ab8ad8c9862423986890096ce1646434f40832cf3552034f9378f1fd2af2caa0f3417d0bf553b4e698eeafe8a8b151d5dd1be65a3067a7f410f5dc916520498526749b073ebff8ab20f4782e8747a52389c474b7754c0b4b991f9cbe6328096005342723bb29e6642b48;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1afcbb9d0aae18cc462d819499e60173caf84061e776bef9008bbde9305c1c35dffc902e907ab33b0a5d358100b59270244c8580c40f2f96dd76043c6c953e96c545f3ebd011528cfde77f4edfd386c1e04952c855c8ce4dd32fccf563808a2a9a2abe21105614248b13b5ab8ddb9a3a7594e1d0554c77b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9dd09dbe4643ef74afc8abb23bf210479fef9294778d30c5025630f03c98e6667e1cf14ea3a6d0a6f884ddcceeb719eadbf7428cc212ce73be8c9ba431a9393100ee3cf71c9aded80c30e6657c28c0f0cf24bb038acbb2e14527878319d233f5dc19262b0acf1854a13a87fb827a76cd600172b7409883cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ca89b8b09735af6ec48430e48ea30c0c359fb170cf882f55cc7aec1ac28657721e45a47f0397bbf4852ad36ff0c26235591f352651168ac937a05a404d9958533d3261e3865c068952fcef70c607e06be646c12b8d16059e09f86e9f5ac879f61cad3bc662490c96c9e3b296bf4b31f5cef643f36eec2fa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5d41f1f4b955a153ad176122b2a65091c61fca84a3944c9e7648482a70342e243deb3e1c5ff742241246494cf0eea88cf5821d976be1dffab8f1796defce497ff44876f3191b2e171939cf5e1d85c4415f75bea8eeaa7a5f49f8a6091927ddb1135ab2cfefb228d4951c980aadb81c9b9946443dd7b515;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176b96d5e1f4a0a30b6526ec0f318dcbc3c5df9405506b26a17b164234256d977306c6340df15d4c38092b2210f014220d285f3825b0ea6e309aa1dfbb52618279a0bb77326c1c946cc9b0ccf318a303e5e9cb3a2d27eb993a7248a4a1a378c7fb89f389eb892c884a00c585aa25e84b886dd9cb97f4eed8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135c9e1b0f14009526a5d17b7415d4077774de0ff588254afe06e512e77fcee3022e7de10c9332867bc7560b4e19dfa435cfe5abbd4cdd65e0831119b70ffbc9ac988312b20807f2116d718411c112d62511b7eab90136ca1f84ef7366511299bf6393b9d2673c47a2547b0c3ecc87a7c77cd248ce82b3cba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96ab365138f731d2f0f2fa481e504cc913497e90783cf94e8bda19de33b58f778107d016d7a3f4f1b57e10894a1101ac060220ce287fcddc94818e94786e61f7141dab93c19e6c531bd43adf1d54282d444207217f20ae9eb3b722cdd62c457e7c0fbcc2760c24120cfd0524435a8e5808bb2e4fccc881d7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fd33ce3d8c416f87fdf98bfd6d3a827af4336abf2e606e0af293d98a0f765b605066c3ba60ef65097b75954519eca9e2b5161f262e074ebb180c35d9eda7889bbe33e8cbdb6d38daff7c85d06633ef6060eccd951a5859e97e47df72763f3ab8751e4a2c72c164a37b8551d1bb7bbff5eb6b7e46729d9ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h316ee1ec8062898842251886d885cd0ab5f83ad17802105b3264c2e7f532868b7398bac834ddeb307bb2e3d25a142ba35f44bf933db34c4c3600cb431a8261addf74f5d48d1fbff6fc5c2f92f826a21b67d20213c8ce52bd23a90574684ea7e846e436bbadf109487b6bf4a42fc81ab4c8bc56e2a910192d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f35194f468f55a66c901f94312516679dc6c211ff1387ec75603f074287a814c449c363f842cba1215848d76bfc57cb0ad86f71e608cc7972ac5f04ba866b194ccb33aafaadc43a3f89e6bff527099e95c0ef18e3f283b2c09d07e9e72fa84aff2fbd3e5d94e88ced76e1e0be9a49d805f115ff15c348892;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5849bbf63dcd0c064b72aa72735b08532be12606b08512a5d0ab19d07906bdda22433fdc613d3b0475aeedd5ccbd203f5d530eea1da47015b2359efc276490469192f204fd76bb329a7c4487dc88060f796d92a0e6721a306a6677b4f0727ec37190e377cf049d31b466b8f9bff5cdbd3ffaa2c87a70f50e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1080eea9a757ebf1e18e831cd03f85fb7468f7816816a3fc3d0e20651ce114c1e07e2f6cc2dd1310abb5a96173b363b018f15b0ceaa635e51f68b70ce3c9e42a187b412f67eafd5f4795afa50af09afd68475da300906e3101214eabe2bfdb40894976cacaace68c6cf17070c4a0e2456ddd5acd73b9e53c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa40861d0c7a9395ee0dd5c34bb11c2e02d7d96e5b7906639119851fc5f367afde9b7ce2efb01f592187c30359af1eb28b0b4ea1c316efc4c0edad4a46fb78531c390dd8b9a20233a7de6b32ff4f10fa2b0358661de4a53a52c7d60d8c0d232d687b88e1ca35da06ea8cd66955b12d7e2e9828417ad2d667;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadbb980ba177d7afe7cfe836e69a5d8cf519a2de4f3fe3041aa08500da584596c4a170fdc78b928fb51fc1f0d78de1cc3737386dacd39036356f27eb0f0ff6eb02332c75ce4bcf8debaa23824eeb4cde1b9a8420d208154558280acd4869153f86b7f7232fc3fa6e5951dca5534505283383f2e9f49ca9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb2f2831a3f0e17e2075cd422b51b3cddb6d64003c1789694c7a9b8e6e61dbeb24d3e507f8e536e0367dcf025b07521eeb625a3a20f801fa21f56c6c44a038fb898f2f19558e5dcd385d25b7d5a81b5df817a153bde505c7732ef0f55d4533f75940637c75a36ecc4e22c4f0cdbf49fb3bbf71847329f438;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb0954759f5513f18f21c653047ce9cad7b46199aaa60c42d2dc0cb7838cc3d945bad503a67be4a0b5c4762ac29d09d5fb53c4ef8d9121c82bc1b393a37f1fff87947232bb932bc0a86d121676d9dba3416d70711279cd501aa0c12af5afa711dbc79f05a8d3cf9fc58aeb09de9996592a822d21fe978a60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf188479e24e7d36f44039d117707e485e5acace72fabe3f78f5477121dd73f1c2d01d6b8417de0d253e085e634c09d232697ae5925cf3f9e2fbf053513103d5a0be11e888c4cd9c1f1ce2672855e1f17bbf4a5cfce4149549af584db4307d1da269b075498e1dbb3f8285d9c3f8855913a78270f496df04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h535ad3f54c8fa4078bb2a5ca32945fddff386e42587a24634536f98a231cb17a08ef989cf7535170ed940eaf697b098514140f6f345a63fe288d25ba6a1e9e23dab52255c7a7c29ee28a9200d00c2ea35d95dc4037f7805fc20d366b0d94b9982f819c227d695a29619f8a47e52f347a6f362f119f9e4fa6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1871d8e9588583968189cb919570ed3525b82338b5d2716b38c713777bda1569cde9a962ce4467630915318c37a0286604a425043f15a941feb351cd502290a5b6b5a063429f09f97487cb3cf1aba39ffcd1d72f56099e75e5cdc6755e75f08364351af7362c43e83b8f4849f231d083b6371921fa4adf682;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf46d764be04d1f45f6fc146d3ed08a5232103cf069c80291aa47a252d0fc483f1f46e20cd08e1429f5bb7abe8e962519b51257de0f15b265b70f27294043a1f878879b5fba0c7a8df42f3787fa08b17a2893606c021895ed726bc9aff3f1991f68e0513f963862a9f9b997e573877075205c48f61b999dcc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f7f6e55a61e7436085299796cd9c07c1670a7e73c687a70845f664e918791b554644975e11e010ddb715dd89b36e13cbdac57bad48cac98d690da4ca92dbe5a441880f086e26843031b62f38ea0a2bcba5ecef0a02a3f002856e8d6593027527664859f434fa00da7109c1ce1b3bbad8510a263d55e7d4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a132b676b584586aad0f49b74aa9f9f8e9406f152b9385eeb65433f32c4302234eae1b7d1d00a23b1406c3bdb52f8285ec81020a46354d675a0cde3dfa6322547bf9f8baa93b5261688ca0e040a49fadd2cf1d668ffe381ec205c7811092ecfe909d88faffcefbf8033348732d75788463150d9a09d4f8a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h933155bf9ba0b8cd83666735a44122794edb2bb877b6fc4b15876a51b652c3010593180b656e95e748c8fe03650c920b4a321283339f7581b08384f756de3d08ed2106b6720b243d2e599b1ce5577d345e5bfe5dbb8197cda47c2f332d45af881953b711f1d64d884e26f8695c91ccc8bf57a3d9fa031c23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151281dccb8938a17b6a01fa719738dd7b187b3bc390e63a93e4d58923e77405cc9a3f1028caa28277c4db45fd1add1c661c868c88161cdc0014918ed4329bb1db70227494ab2d9f571e3fb2e9c5bba8f4955a820bae735523164044954692009f9d86a1a06c70d98b3f0c196920b8f9741ef243b9ff246d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3630e92cdcbf5be920826b711d655a975fef5117312759528f7aa83c625ecd187c95b99fa509fa548792f468f5289f92fef7087dab29e366b374df1364c848d970601d099b88eb948675ddbb130800f64881ab1f03aaaea2eceb4136d35ec22a401a8ddc86407dbe72c8d22ff96be47115e024c9c1f3ecb0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h66dad4cbb9f10413d30905d4f2fcac6bfc61eebf939876ddfc283acbe62b21a42192bc47a56ddaaf14851004bb5991428acfb0c5a2e8255dca58a97edaf3d7512e1865076201358b2dec9a3b0bf5c20a2fe13c8a8296d1aa3eeb4591c52ee37db02cca84d9fad5e74836093adbcc13fe0d013bb000b498bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3d3f411a783563c6ba2326e03abe8f4120a818ac3648523ebe5b415d24c15100cf5246d5eef185e2977e5fac6f54106bf902091ce5bb263286bb0f1758648d4dbbaa9abca4ce4c89a9ac4606cb09f6eedfcb2f773025666b6922b3ec4f85e09a3d1e0d2553d6d084b7f7a95119463c6e3f2e1b9b249a82f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bc997466c59f8bade90ed9d2aa3c6cf4fdf67d9f7ce1adcde7d9a4dc3bf39170d27246c860e6d131f8b4e82607737784bd581b9fcdb949b327fb00d7f5546b12fa5dad236ea9934d24dd50962fc94caa0726ef872d49c5c304d017c17118859ae1c2590d9df42f8901bb545871e41159461bbe02481b660;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb21278fc6140be3a8928d257411b296c701e057831c643857d2c7c8520e7aaba280f071d838985495f32ee35abd3267664f59f7f8893e202619c0b3ac423527eb67859ee899408d30794861dfb7ac7e3fe8b4eb641e76dbae242cba0bc251818c10dfdc17641766a9b64396bbb3715debfe6caf9b6c2d41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5e761130b2598fea7196a8a66747f729944eb4f964c8ced59d0b17f07865cbceeb047fc65621294f2d09f5ae875bf61657a90e0b32b6eb976e3d293e3c1cd28491746b440d4ded8894aaac7bdf083f56843536026cb1c3e97c1506bab9e62cbb01189aeff08381cccf700f79bd53dafc434bc52bd37a8c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h798890f8456e7a745f2219d9c2a7fb6b81901ef1736bbbd88ba9f96b219cf66a30bef3c6b23fa3c17bc1e264a4d5c7760068524bfe76bca1d7e7d8cd73ff7d22c115d332b7b1476edf67b4bcd1d83fe438172582a018c223d751256da2a9c67bcae5f3c2af784d820bc810b650d938902a32d96f9e619954;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe2640a0e5ba377f845e731e3667174b2b298a8b3b1388302d502d9b452506aaddaf7e46450ce5210d66ee00069feacabeca7d3b07b5741e3a8538c66825ac6b935e276063b71e18f0175bf66e89d93ab4f1c80dc5f21a5641670da845e9d47530d1b33a5f4a4f9483f96e2e0e0627758de128134ca2e069;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfabfe4f50dfb22ace0e2c0142871ec10887ba4724d13aff11023f2ec290aecc0372848b26252abace423839445a0b217debfba6f1642824f14801cc0ca38ed99f6f5d59430ecf1bd7327780f81a409a1df8bf93226b2727a6e621864c35eba1ba7db5d882e508663fbdc4a10e6d073ee4ff4b992d9d680cb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6d32a6b24e73b6c0f2c8a5d3e0c4d2daecce0c53a14dd75bead768db6685eef49c6f00c94edf09dfedc8285a8a54f6277e5b0fd12c8a4f1d827eee118423e22672f6acbc2d25b94991dcbf24b7748e690c5543f340a03760be2370fe675d1a942134b3d8acb8a6c9f40daf9aa30d8502e001af6ab9b3f10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d08276960f4a12735bf410c6684d00a7cd3a8e56018af2c59f4ca49707d39ef70f2efbc4dd8bf3c99c8dc992c7624bc27109e9385283688eef894ea9072dffa52d9d5aa9f6f4d766707d341305868b4308f44df1f83e13eca0bade34812a8c6ae24101a925254bbec453a04a91a2dfaefd1c94a67ab9494f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbfc1e86923ece0ccec061e8729c4a3c014788bc7ddfcc56ded73210de6f227ca81960e2b7c94c3e4b4be6ba9cc9c9e6e09b5d2c5c494ce3cbc89c95ed9c850a6407e3ca77b4ec5a150fb7d74eeebe83e8a3c1a85001ae3578076ca46bb1ea356f8533ef96a99ec2fd71e78431354bc571ae2b0e4fb774c3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3700c1153b0fdfcb4fd316891615b8498a97199f15a5bc58f306e48e523ae423372aeeb48c871d9aeed787eb0808719b4da20cecb5e2c4d71dc5105271b6cf938f6c11e6ec3c64bf4e2e3ff6614eabf0ae97cc492dd450ab078ae1b960878a18048310a0f7362f13fc2554e05867ea55f4f68850b4083c8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f8a0199af78e39efc16adbe40030114d625073c7a8b8bf135cae896eec4909e58ec8ca34f5e2597eec1cb3f502193a67483df451ba295f6c2ba0bcb99ba114f3ac2afd9b4653344b9a87df22342a736d3f6baa9c5f82360774b375b62e6377c1220cf01222d4234d0fce52469d06d80b3c7c859908d9bbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3265cb70bfa987cdd9b836aab9382dd5281f35fbedc0ecbf5a9b38c8519030653dc847da94469f5071cde3c51a66f8ee03bbceb65690a5e8a6f24b57695b8b9c06b1e52c926a185ba0fbd9dc9cc1412adc0da2ba0b564f5c845ef077c417328b818a191b0406f2fb56082798e835ab2a3e75e811bbd1871a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d11e729c832836de1422bf371fa337d33cfcdd52f31c50d51e8291961d661d58a05153e0aed8ff3c979434aee84011fa98daddd082a1b1ab2a71b98097d046f6bbd56a1ab883a4ebe42f83a32c60bc7935007333fc7b2e23ef4d110a65d384f7dea71cce132bc61fca1fe93d157956716e44d5e986072e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1950a882c532de5274f6c00882678134f1f91bc187595ef1ec74f89369151c7f0a52a08418489fbb824ed8c020a6c4f2a34da49c6ed46c70cd9332b12365724920b24a41391b1f733e550f3a7339a596cbdac66aba9d36713d0d1b5480c4d065b48f2fdc7781f968e54078a2b0d8e50aba721a7b090b97a5f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11554123af2e3a208e5e1371eaaaa8744d0f3539b08c0836f92e63724bd0430cfd342f5bf8cf7394fed64e3b7ae208ea785887977943dbadd637522552b01b1c079809213229d20b3930d2689de05d6be5316a4ad1d89971e0d06f6a25a5bc20cac2ac02d50100e8d54ed5cc17fa77bae4256d877ed0f28c5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efb5a000ae5fca4adc688698f4cae1e7c17163f372b831baee62ce3bc9fd34278b185d662d85eef5cdbda1025d54e82683e68a5f46df01ebb0520f5b3ec7dbfc3390c1ad93b18999531da8ba06191721ad3e3314b8fca547d174a03b711146034f25d95bffa6fb33f4bce3f5f872fedae0d704374a36327c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12978104e02bde329301808cbd098a4c20f5eb18af503fd23665dffa7802789801252646300951a36589889787d8b4b414bfe17a5ddb0fc97439d9c7cfdb0ed502e96c33f0616d09e00822bbc04db5982391a7845e067366b904db643a8195e4e4518b984f27dae9a8858b3d13baad97423deb03e50c7f3af;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c252ee35046356e0896e59cf8132d61083b1a1f4f419d3c6547bf4b47af0e6670d21d55ce2797e714699bc78d90baa44cfdbe36d5a764dabb22fbf0a5d83329dacc58cd5adf25865c4624a37799d13425af1b28dac283af45c6a26d89b0d452440e2335a609afc04bfeb3ef98f7e3dd159d7fbb71b06b38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0428dd4069794c9e57287c13062b1eea39b0100baf6a2f68a505382ba7a949e4c80bf48eeaea14c88447b5aaf26a27ae80ddee50dd83525b91b571f65ad915fa93ec666fa8a001f38522126a447a79dd05522edc903b69228ddd0744e43a87d7fd823a8d56abca6da8a78aba9334e221a852837e046a2e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119c87d11132e0a7ef8f7a62f56b6acb9c1fce02b8f55176acaaffbce4a3a06302a0dbb6a1887c8bbf28cdc5ee392d05c55833cd14a078a2f7f2d9babc153c06109bb9f1610965ee0cb9e6410da309b27f82c83ca7da14660dcdf71e7a351def0a56c5ac9e5f80f82ec7ec96f0bf98b59ae61a01c3d07e68d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1161eefca8b27b92f45e264b117a00bf80919f4d567c4960a018b226d3cd1f07e2bed18ea8d2bddc3f21728585c740643fe3f9e21ac29536ced3cf22055401253f6e634a6f8646a2891b407dc1b669ecaa6a4a2d4de1c89ff71b841083d3bf6aa9fd0f742316a870c21d4d6d1ddb7442da63cfa9832e7a1f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2634ed267c7d12162a18f043ec26cc33f487465475ee4724845534c2a38c3b2b29ea346f9745e4e9d8522543a6f7b9f76bc539af5686ed6b22c2d1b38fe52f61747b0ad71a7eed0067d98929ebe0102c940c7eb8f7ba969b5443b79721948190fe31c7a61dac6505cc2f6fd2602cfe9827aa5dee940b3ec5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c4ec51eac36b39c7d8ba0261f9a70c706350de80ecbdbae7730c8dc4afd5c07b0822a1eee8bd52128bde72987c8ed7af2fbc995eab13f1b98ef6c9663cfea0b864279a20000631a9562fafbea261fe65a98bb451ae05f61b39f0c29b3608273c361f191d4997d2fa4b580af01d67af3dda7933b09ef8ff2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb7c932f02220acea6a5ef76991ee517616a7b33750234686bbd3fbeeea0267f3addcff2b9c4a5bf904dd0f4c7b7941941a2eedd129ef58a69fb67cc434da65ed3dda443d1fb3b451a78eb9e2a0706b4d91da1c76011c53c18c74369053aa25e5f9ede0b40a0ab083fd2fb81ffaf0cbd2a81c1947e367439;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f056232d243466fd026c30ae7c7441b66579f21f6e344e6ad730674771a6d259e979dfcdc0e8b53a21d3143a53651023c79e634b82b450c6edf69c1c06e36a83238bd88bfb5a6d24f960cfe47a982d28429e828499337bbc298155f1ee6de6d7878595e1810cd24ce5e5e1b7c37521132fb2ea00f63d09d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1004d0b5da3b1d6b58a661ef4650664e8178acdcf6d6ad3498cc7a3d2fe96484c6f8974250965d98171b5275d9f53959da119f0e5d256b41e535900772eb5802e45e0d15ddf712fb3026de819e252d1cadc757cfb3bfc949297a2705364c467b43702ce05e04ae525ada53e3cedd7a2056d63132bc784e0c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h522bbd304bf1e5670782c2f674ff4f30267cac1dca08022e42e2e4d0073f6570092d17c93c48f7feb745fd1a6f17a51470daae20696639ca1ec74f3e2c8f4318bade7d23aa6ae8460ce0085ec5ca7379969bbfffc207f6290a24ca7150285cf93642b4a96f3d88fec7993619c018a2abe6a388977ce33e89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c039a5c446f6e7f4f0a9a499fc5bba57f6e0029a636511ca7e83eb36b0c8e5bd5989e4b7cbd8a78276dd7b06e3c908e6b2a6e5be88aa8b8fe7de5f30541ebcd3e5206d12987c9b7983875bfe8ae2a933657ab78622dbb065942183a4a57f1aab0e64556eccbcc54852cc5082e3423bf4dd1b662d990f8f1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60863166264c984e910d9d3d4f763660e1f9a05bdb261d0a7a55f649e3c417a4c7b0d45eaf532d7698d67826084b101fea575edb20d8f1ec2a0712a4a9464e4c81ed64a43ea643eb87194c7911c112fee6175e5338e2b86c9911241c5543c404c1c2ffbab188ffd1fe532e96c92a44765b0e09b9b48c070a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcc4005d8c2a84cdeef25c8a933c04639700be46e518e3ef938acc40ce963be34cdd5829fb96092d6a7ac0102378862adbb6c8ea966d9e4381f28885000d8fc7c733446d3ae854fd7ad9c7cff08b9d10b0c3482c037e7e3ec08cd78310c4a24f9dff47616124edb2d1089c63e43e3e5cf1e3b84371a21283;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a6c5d85917789eeb2da841abb28c98b13cfc1de656638e0689f76c5be8a326c45db967e2b17ddd49404cd38963b375c129502be6124b58b43df6aa08b9fb50d6cc119253a7743dd71e52d4fc57603978708037ac0070d79fc0ad43dcd1f0b55783907760d3ec35ad1f6ebe487fa5ed0b5e7509b73e9e29a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169e571c2997e7da680cbcda18a8de8d85aa780eedf09c23d8ec38641df4e4d6b2bc01dfc4018a1dbeb6e99928b6e939f8e292e9d7db02b626576e883d386d1d2abcf90abae2b233f67af714468e413f5a67913a8027588a1f51b0bd6ede5e4b064495078280048f1f4d96cff1956cc69fdd36df4658b76f6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11da6a9e5df3bc3d4ab719e04d11ba0fcd6c3d91ee2ac736a72903169a26ee3c7b53f068e00014760bba6ba5c1a1fa97b524a8b95a4c18a32e8c9033ec2c2547d703185bda6fb7ec08ed8babb05620332635f00cd80aa647c2587b840dbff605c64b9d9f3d8f423f9293ade593c057ec5ad6e2af6b5fd0927;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52e4dd0b55c675df0018172efe5e5adbbc87a7694ef875165105fe8157ddb2523f81db7ec2cd2d942d924e324b531dc759c82b0225b9b613a35ae197a739b77813f029416dcf657862cf5ba763ca58a5ef16c7dabbfe25a3a17be5f20d9dbb93d727855d10d3fa3f11acfa2f21631993a53bb8d31221cf5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11061cc40f6b25e37e235b33d4ab7cef6bd97e275e23ecfde759196665bfb5370f7c6405dc40aad0076dc1756ad3d2a7ca7a48449d0baa0d9c8fdac817afc2a33008d569c5257f3f7c720d72cb4a254e8572a314b4bdc0d39e37749086fa2567d1f79b7ca86f8d78836e2f785522ca8ae6460ed670c9639cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1ee6c464ae03219b249009fa834ed31fa011728afb2efdaf3cdc88f56245e176fae4373be1db2eb0528b229f1865f2bc6cb8f18e558f7eb7fde035032f246ae6303bfe83a384e1792ef10ea2b776263eeb331ce721f1101e4afa2cd7261841126d63eb25191e54d0724766d0e46ecb15c1c1b254e03add6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h454fd7edd1d0f38605e11690fcd83f8f5f7c336fa5f6604b82a029181e8a4feddf2f071a36b44542e837a49563bea0a7af68d474474307aaab2b3d86c3908e5a3fb1ba8f0cb17ee1410826b405ebc2472e57e054def22847ade8b47c6d977ddc6636a5687d9fd1d6b9f92619a89b87554057d8663a72efe5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4a05e7a8c702ccca10d948f0567c9b188f518ac87a2031bf33b3a0cc3192e9db2fd99a5b1c7e5e2a6e820103977a9f6442f4e3ae3d0f0bef798060f8ee0d5fa16119b649ffe71aca952dec564890849fdbadc25122e7ea9d2dcfb0d8bc40c23b2f9c1e391c3ad98365e0b8fa336ac01013732d2a1d4bf34;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58fdb887d784fdf3b499f50745fc4c7a2e28ceb73566c8919670e059ec7dbc68da1f29a961b100321cd4780dd6805935da95919d497eee7530b6240f7e58ea7c52c9fa87d59d32854b9c470a170e4023adf5f99af9b4803a534b63cf4d4126170e4633c5d2564c7470899fcd1cf0db684b31282df5fcb520;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c62813e955b16242706407e8eec0031859f0046358506e53635cb0d693ad0c09abade2b28b5fa2f76e2b97991449e1822f6f1b5c168310593c9c0883fcba5f797c7de0913d741bc7d74f53f848243b48f0f37f3c9ec1e5c39fb1e419cb1ee3b4d5b360c9ebccff126ba66d701ce4d589cb25f7230883855;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c977408ca32dec62c731d5c1936ee52bcc8f520b4bb16d0e66f769c3d40674fc3fbf3a279e4d7d674d633d13d797ee34c3d71a15da045d6ef10148ba377b52f588d1d4f664089432033afe5947a0d46800f7485d2fdfa18d1cde2760645157d7456e59e380b686a9d9bff5992c04fb1c0e53a7f74f4ec7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadce174bb3c39a1e02c8308673bee74069e6804dc1132f06c02ad24cb7dee336fae94a08acf70549ffd92aea8a18d582fb0e2e20779cd67765d8eaed306817fbf672d76a38e4939bec68121bc98bfaa537b4397eaff303a6f41f05c37fa043234f3eda951e88e044dbee7ce4745ed65502b42e50ac12bb7b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49d0f7c145ac9a83ce26dce5a7dfbd6ce687c2a24dd1053923fd28b28497eef8896e79f913b94b46ab05b52fd6590788acc1526844e5cd7b1c5123e3fe1ef3dae4ffa33eca55d41e923a3121d20d6d5ba10b1aafbdfa89064316f10a645772ad1d8ca5fa7671d7f13d528c9efbab8204fb27ed1c7ad9499d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f1e1ea7b8b1ee0afae363835887c149bbf3401569ca26b924473f43f3cdcf937a514d5f31fcca8753ec660d9a0e33cfbd37c3c434c11264d4408562692598ccde6dc3502813f0860dfa0a2a4c631db3ffdc3499d7c17cebac7aff4c56007684718ee2eef623a57d8cd50e21cb68b999ee786b730621b6b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c92ec811632fefd920db0267f13d276fb4df95c69549bfdad2c92c2659195d4841519eec4b067ebf4e6e3fc1fe68293a477ca0fb166fbd7af05597a30b94a9a86d487bc60bd4a7e00cf03a894d6d6e66ab68af1151418e87f77accd4677402b8ee91488bbef884fda8cdaa9b5bb5fa48cbd3a83bb0e94da;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15834175344abd0bc57cda00681c252ad7c8dea9492da10031a741deaf0a2f0a492abf11b28779278fac3122771c9dd1fab5ccbe9f1a7e22a3fc1cd08cb32c2c8ab85e12c502fb9fb428829cae0a9a24d7ce8aa863f0dbb849b1574b55f0123293dc24d11c861d9e9151ccc1b07a8ee49f1cb3f3e2af42c7b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ecb05a00fee9bb37054d18529af0cb35748febaad6380740fdec3f8c22b8b01004b52bdb9c5a9565aab94efcce5b61b84ecfbe497ff4f5b1956a82cfd7d6330e323068bd2c0e725f61387709ab4960695e552686df2987c42ef0f1b3fc7d33b6ac8574acbe13fec5c2e2cb1b9b9048d4cfc10644681f2fe3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c56eeefc86bcabe89868fff644a6eb75367d4c75be33848b737f61eea979fb25e6b071829500a9b7693e099ed6a97e96a5625522da6b850dd12806380a1de8ec118c2e5beecd791b915aa1a1fe85089ad714790950289decf94d80bfc62922b4d68ac780af9637b2f12da201a86be3b8c461e4de681243fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc12adf132155e611105b36286394ff278fe7747ea255bd683b3324ed3bc17a14fd8755f916d5455e37b04b10ef54a036999b9cb148f49b68ade98599aef865b4e897648ac06f6607ce4dc0f2863d974c235727270785f1e5f41f0d58aa7de91ad74191a5a9612cc436bf15d85ba2d1c04e3729455dee4e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1808d59c56bc076242965c94b97db4a44a0d379f50ecd579e563533671baefc3812d853bcbf6719e71469ce7d789142435002825b0fd840c6b665f441389f92bd5417e25ef0fbbdad68d49de996ed160420a252d1abea72e62756e716816cd9893a9a0917cb28bebfb1595706b4874da1535a07eff07268cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b82007863cca5b5a3e639098c3ef5c291757233e847d2e1c672eb5b34bb999305bf6457651e8b6fd931c8b18d59feb503bbbef9b866aa551f51df2fc30154ccfffc3f6fa6825382583bc46248a846dbacaa0051142efbe078bcc7855ff03fc1432f329ed775a6917bd4b15bc9579d243abeb13e81690504;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e24215001db75479b3cc2725f6beee3d3794c9d7977c8a5a3a0c97f63b3300e6797d5db10271b3c263ecb99652d9c2b40ef30a8d2795372ba5911849ef12ea896c53e92e659a669a610ee014f044dbbb498a9f15a5da13135f99907373463521b7dfafc9c038a7c4788a3a4b0e5c9c8a7fb6a058b9f9b811;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h563ee2d0b475fe4461937dfb6077df32dc8c41b290447bb8690dbcd755cf725cfde10fd30b45a4a7206ab13f566a05e1bf4687fbacf6f2b86bb8c131e5634c777ace3269f5686e9b948d572794c967faf1b8bcd14a85448820945e854a6dc63bf0e9b0e4b781a1b5533ce721b0383f497118662ec65911a2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9c51bec97411e77606d559ed49fcc61ff125cd7e1095f5efd9976402e4989f53c2e409bffa938cf0d7fe3da48fac4576b0287ffc7a734bfad7efd32dd8a6d975851ed9ba4e1198276e4c69e05d0fed2f28dcfa5b9c553aa4d3679ef09ef7651df3fc59b84bc403b8bc81e26adde4b05293afe739e795a54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b9281b145479ba6ae6102aa29e8a3d1b59b7458c4d0e5ddb694c9fcac3b53851006609c91dffd18e6d664c75802391889c7dbab7c159a4a02fcd9554701b677a8bba810ca00f2f164f6fd9babdeb199408518428727e183c7b33ff559debecf726fd91ed47bb9330bcbb8f42cb98686eb785cb60bc99be8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18be8ffcb68a9138ed84d9fd6266325ae0ba3cf26bfff19c68875cdcdda70f13a81d1d9c00e0cc05e59fd5548c3579b916c5fa9a2dac6573bafcbeaade92f9fab92eae5d78304323a41d4e3747b624228aee6cfea259033a7972e70b6cec73fdbd47bfa63189798b85d501ce5e334e5f12c162ba4395b1b90;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13bd5de563138cd6869f336410c3fe159a52697763055009779e926f51c2230ece622f792a49bf235ccaa97725b30142205f6bcd0d93ef794f97f1f22f1dcf3157379bf62f3abdc5ce094b169312079bc711e2b17eed0ec4df99965bde67cbfd9e93fb3c4acf8feecf4019f0a572c2229dcdd066557e891a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9c27f394212625373bcac5d0116dee93f18a3c4fbce76933d0e50afda19485f79b597a7a5365ef18fcdd222d2fd5ba49d2f3ee39a013151dcecc8afa80fe8e51f0f27f88ff2d0ba0987a8f4633796737946b278cf46e17835c965d5150015d8f382b37a7649a82cd87e00a7b7ecff78fdcc2f730d1c69b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5ff1c6565be9faa0f8041eb4d1b807cfeb0f7dcd57334459159d048b9698a3c59d3f2da9f0fbe9e6f05715bd2e000f15de35cbfaae565bdb8f16b40d933a31dc8ae610ab2fc74a363009623bde9a0890394cd345bf7f71dd9c2e7e82ad5f5fd2f155dc2e6ed86390064ce1479191dff43174778855e1004;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1241b3472795105b15abdb66439def21e9a2be8131e1b382da3e037d79f53f73c601667fd36e7a0825817b434ebe4c13cde5f32f540f485e2029af4eb356d8f94c5ed16f52894e949ddbb09c31d3aaa6d621c6542e9fbbaeaa35dee593eb6fbb26d699b75105b8fc0b5078863d4625a0f921a329c90c10743;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f15c4c46bdabd684dbce45e1aa1eb48f41cbd04178d6975fa31620ef16d820d48883b8454102661f32bcddde2b82b325a07e1416e834c7b17913abee35d2a28986e2ed90884a5358533966908645a0fd73681b2c115f048363d48557659b11e67ae82164ec5380d2127e2b53a7e08aa5751b38b6632632e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2aa0b6d4e5ac21db0080f03d5e3b78986c2fae2b7fb02b068ccd4d440cceebf3aa45b7f840f707fc83570d853b42e2d3524d7329c0e453320c1b30dfc52e56cc069f7ef3eb752068d91d643bf244229d316fa8f6a59cd6fe772cdfb4b7f970774fb1823dd6445880f9bde6899a67900eb19a476385ce4c5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h378bd0a430059f7827971ca1ef42da97090db629f12e50d9bf9d64a7b56dbc89513136f790f7118852731f1ad1d0055eabb204128605caa247c8872d75cb6ff63210cc59fd05ece972a9be791340b5614a570d6d341404fc3cfa66c66e733dddba9f726d816838fc00581d4607533fd56d0d993654f68570;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1571149210410e04906e653044c138ab105a4d42ca5e8bf498bb67f6001285ceb4754306baac3929474301b51abedb99fd4b3e8d3de8040b0701a8b048c18963436a865747df8a896b5063e1673117b68caf910b85188a24084d6cb44619a0449b02bbf5bad5a659498e358c85cc4ad2613487ff754d8eab3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1518fc647550321030204598aa39491348f859f8f2f7d4b37d0b2689fba5d3f63f174cca78b20b8739e0f181155e515a8d46e8ea53426a1758a9607ff8af9cd4c05880acf371950658bcb90edb93f56ef704acab6df474e4e4e73d68187ee1cc672f70765938c629dda4a8659e6e539642d58a665b58b19ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49cf4c5ed61ee1d83c1cff547b543e03fad77dc8bb9cefbc23e90b4088ac37d3b83dea551d4162565a763c17b8bf9770884c2a2b3c9cacd62914925815bc14807e89e44547f17c1f268d04e35498afbade09117a6894afdc2e21c3230bc11fa2cb135f7e9c8eb793a96729ceee9dd03712636b75af41d3c9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27745ce784984d251fdc96c3b1e477284346dbfbbf970baa27c5493e48c42ccfb6c82cbaa132151f39797dd87d82b28feac91dbe6582f8ee12bd21a373caa0f93c8114dc9e5029001c0686296dbf6b914e189aed4159f6909d8409c22d46774afa8a90b637e13eeb05e4efab79076559b4ffd36ce1a06783;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102459817a3aaf8e50849b9022073a824ec238d973cac4dd5727eb0b8060d67656e48f7990fc65cb93ff7c8a8cb3bb11fa3d3ea31f1277ac46126d8287dadee5c387f6e865f8d263187aa853a38a406520654b7819a99ec11a1bd0ac09c8e0bbdfc75fedfa61462d888329eebb2893858c29ed2a0c8867b5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1885963cf8ca987f28d19396cea68e2bd8b9aaa274bb2b391d03f33336be125ca3a90e9b9675957f1bd44948ce1caf11c76a279b8aa71d1e2171412b8aaa23cc5cd8cd5793cc5c1b92387e13d97b24a42f06cc96dc7baf5456e5e6c2a4879f3df979801c488adb33f6f3ab50574d980b4bb925b0eeb05023;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b4e97c81cf80f03a70bd012a36a1d78ac3e99c03299c1cbd4c171bff51d59e13b53c6524255f0c0cd69a915147917200d4f633420fbe280c8b39a42e90b8d846eed57e7758689f8425b5b39f615ba6009cc2f21e25d091b60e27a016ce0e651c5f3119ee3d9abf5cf7e3e3069044852b3dcf3fba6a024bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51e5b3ff49e5d1b4f18b1a9bbeb9e01543c15afd5cdffd4234025423897e6892e9d9ce81e359bdfef3d8127d912b95ad668cfc6dc38aab6686c836a6a42c8e068cbea0a53f88b01c3195af8a3a623f841ff01f0e86f12b853601c84f624d428b398c59eba9487b826289c3092fe53cc2ba8b67d8bf993fd8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed3902a8ff9ce760f557db35226194243c3e9c02326ec993280817d3c79779b4785048817c3e6fd4f6466b647dc81ce15d0202acc06df13273d34093c2f785d7304c6603cc4cae1488f97a6f53b5c2e025cc2ecbceec816c613dc53d712af4a9e39001ea493f07dbb543f1538578c63e8c1a870e57830ed7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151c56a702fe8532c0eead6e58d0605e61297320ba05277cb5074b059a53bac0497e0fb344c8ab3414c68de8df058fcc89b2c8979a96662dcf5961f9988a033452be46f56d784fe117c4142c383c66bd67576ac67109a2d95e74bb66e119e2844590328208b70c4d1272a4eb99e55ccc81d8c0afad321ecd3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63bc65fef20caaaeffa40a618f4adde26fe44ee4d909a3ddf61cbde2ab76b5c659c994634e47b2d302b3e738d68f02a839b99f0d7ca261232e90836a249f0829de983f418169067fe9d3883b09d2cceb6e84511e2ab562d3582be60e88cebb5bfe609ed9a3d33a31f42823b0ff804983958959cc7d991a7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f409b90922edab18388c8f6a3124ab3d5c3e32f40c34e18e84e05e47a745b6d58c41bb411fc5e9fb0db7d732cceeb15ae645961edcad549106eeb597f5dfc4ff9b7524a36f3070bbd4c5f30f354e4aa78995dbaaf41ae411e9196d207e31b8403258738efad0c5ec0205a2bc346320dd80445a84ceafbfd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1718995383fa5668e30536c8a682d4352802ff464e113f930bc6d89fe4a95e3be6db63e1bc77120a264c7c71e272852bc50ddd81aaada0f82668c0e03425c77bede4af98972ae82ca552d34d859b177434f7e62f1245eeaac9ad84f20389ef905f929333e07bc7c545377dcd010c88a0cf8e1967bea961398;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c4a2b020859c87afecda849c732f64662a7e99457998b80d19a0d02bc3af8842ace71d95d9f5c066bdb6ef44e10e725ad9e320d38768b1d053c3b086070317aa486c191225d3c6fab4a9ffe7c45a017e7e2c230267377bb37a558886c9491deb172921ffaafad1e241b5624638ce54d99968179b21dccf0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5b975fe7dd6d072291f6899b7dd24a311e3f6f7a34fc2ec6ed0db5f18a13eb4dd9a32447d556f97c24b069e81b7e89e2acbf8722de418f4ac040151e74c063f74b45d4e703326f7d6a7cd81d5cdcbb3cc7353d4ae8584de1f8631fecbcec874d8ab94da03076d8de2e35b217338aa176e6700b120d65289;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b2f02fda4f99e02ea0aea5206b73b28b34da6479a55d9128722517cc01d6bd72aa46e960f1cc972df8052c8379c1f7447d59d4c555cbe297482ab7b554cd491e0ef420e99bb66e9a28a0cc30f91f2701f169ba7db27ad16371f0b9f5610b0ca8463a93b46cd62eda140cde527f1725c630974fc5f983584;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e84e3045d16491f77fc11ba9d7b5f4bc1e3809efba5e35035e9da0ca51db370b9516115a53dd7ddf37b4dae72985ef85b11d9ea9668c67541ee19b84142c1e893a38d96b5d950f7bb467f610404c434337d274a2994361088048a4b71e2f8d36f7fea719eeb218669341da7065a521cfa14da04787372946;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94c3174766d7dada1d229240ab16c2d3bc243e6094ca794dace22c92f2c73e248432069923e53805093bf9e170bf53b69456e3e7f854e047e85abe0014f84a817b73135988fa5ff18bd2f7a7dee9ad0a9adca395683e83e8e32cd6d05b3180486a4648c4e9fee97658242715cd664dcd634c32fc7c0b61e9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea520dfb915c02d5af166082d09a459db4c55e68f368041beb42cb49af9f5cc4396199cd9639eab5359a040b16f1b093b746698d6acd77140dfee9e8a3d04bc27cc0d31e3a1ca0ba0b8aa700b066bcc9205ffab0d4344ea170897c63ac6de8a42c0dc2bb26530609f43445d6b6e959d858ee73e766eb80bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49a2b64408249973f4ec4c694e3418413586a5ec7a83f91c8ab44f726eb746334647a8aa3cb40d345ec6d088c17fb04748f6928bb699f3f58a8c6ceacb1aafa07fd8f083687496c103f63d3516b0571ff2eb1ef88af2eca8232ee02150d72888a8080a5959753625b98a95047ebfeef1b75b697e0dd3e787;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68dbe38cb814eae215a14721bb2e32f4bff1e2592e1b9dfdc243c5dc2da0a7e151f372db191c647cef1a8a92e035fd43536bd4bec62d01a2a24e5d9f7c1b0a9bf5e63df14250bef838dc193b3edbbaf0f8c7ff0137e9c16410900200be74dc7a1774c925879ae23a8ec6f39a3fab634de629729b34169baa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h155f3c245551f479dfce26712b6ee1bfcabedbb960414ff57d4fe533b9c6a0dbf6cf4cf0bbb05c751ce38b28dbcfe836f8df30050a816cf8506761cd1507c971d9bafe6d16671df26c8420c1c97e23507482bec303381c2e38107a62f3dda7cfda3f45dca94c732cb6b755e9013153097a47cb6d55f01f6b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h931315306c36d054d957c5fc3bc3e0c2a12e070270c5f28652be65b8fb9f1f49db1c907ebabeb706122924b6a9e0a1838549f61017d560c1da3cb6d2149f55abfb2c9c76642adb0b29a93c158785103dc45a145f40bc7f04327263b4eb8287d23adf552bcd4203d8b7c47d3f097d6aae684a1043a53a0d8d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e90f943ac2f1ca52bb4e9a3a5a423bae63864d1d0e13e46f8df0a8f097b3d97ab1146db067d0ac3f4d555e147a4d24f135c0d1dbd88b6b41541082d9d5566ec2634c3a08101a174992bc6ca7aab0c79c36b758207882795b248f2574c996351b1a6f153b9ed52a245713460bdc09c7ce39a5b27124176b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12bf81d00738bc7239e62c3809288dfc45b5021aa335a3da47176a2c12cfe41cd84c18f623eb59eb560f9826af7a33623f1f2ce1d7968b5a3c784b51a0c85f938402ff6868865f02588469a5e81a651a5835c5320845f8a2c1e5ea0434a334a7071e54fdf9a2202cf052efa365c78073a32bad9f06963f6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7e7f1141a44d973a2dcedd249fd2dc4abdf27376148396364c496a488fa2cd3ae539b55f2c144b0700525faf589eceaa1c4d86bbb8fd7e150c37166a77101796a717359ef0d22f92a15cf03753ae377fb1f1a5a2ab68fc72ae60383aec016bc9364b6e2f88b04668458f7fb89fdb616a6c37e4be4a28876;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hade5415a077ea3b5ea438236c2fbda2740fb5af209125fdb55bf0aebd149a6361dca79272f49f5acab66ec487d4037dbc300e959c78f1e24c3bee35d30faffa91352bf0b286f9dd05afef0a64d2dbaf01ddfed25eb986cdd99a9d34aea4f2439061f7cac7ae2040928b979d9b5a84f03f2e4c7c55a9ea255;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196ada8ec89d5dcbd7946d3620cbdb85649195e77b712e14e6edca27c9368c1210a9f9728153dbcd5ce185205e2be9db360ccf2c416055f3bbc0bd4873433d24ffaab14e0af329076bec408048d0fa01a56373ce5e3df710dce041425c9938e3ef111cdc2c1f32ba0515ef81ad8efb57cd8a9df45144b6706;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h717aafaf35042b0ba2d37db3664263d1a9d9a10a1939508f6ae6ced6e4f3e5da02ebf89395ad6c672d3b41234eefa501a8d09d79b8f1b2862b47f04cf0c7067cabc18a04138d49fb071dbbd4084d0cfee381337c4447678f16b8fc74c1fec2307237f814ca71d462bbd6378ece9b3df209f691b1b90bbe91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc24f078ad503862152effb49640e7bc93f29afddfd38c7295beea7472038b10f37441cd3deadc0ac3d092a598f8ee1353423593beb12df158bdb254142fdcd294ac74c2cc2956c533c5b27e1ecc781a78eb4c9ecba9424ef57ef69e03a656c0de199dd0ac7a7e35629f7c3fd81b0b1c1949d76aee7187356;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a544e39a3926095aa8cfef58322170e14d19fea507555cca91912c4985eaebf8492cc540aad6f984a725da4b3b7ad459a7b648b435fd3416cb101fed5a0dba4727bf1361518418025e17986a332f1f8c4d6b2c25197ff52b3209ddc71502a58a27871abb05aa1695f1d8acf6888faad1468581733307bc2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e079d9b95bbe79600f910523e08dd3ac3aae77103b980b12ee1f02fad230dec827a1e16dd44da604a5f112c7c6bf6c77e756436ea08dac6af334e436eed73d1dc36e3e78d52c2f741b5a657e7e0247884f9b26269065d4d2ecca18b15e58909079082de8209aaf95795f52b5ff76309742d0e98dd1de696;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb9ff858e75bd7919b66bc6fadd638936aca828b31c281f9e2178b3c05ebe4eeba29df8df7fd3341537441b9ff90ab1b22ede06864232c7db63f1e12a4df071a8603a510fb8ad17292f82a6469dd8ab7223ed24ae09f3782fcb91565510a8ca4341834bd65eae50180f4a7d98726844569542da97d293206;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29fad8e933cf4f2044e9d15a64cbf26ae74a7760731d411aed2b25d152a1efc3bc1d513eef40f184da17ccc2f4e99e7d1f89b6f3f89dc080da818e43a04eaf5f4cd4ed3bd835b99ce67a7c705d62f5db551d12c3f5bcb1de9372e0d4ed1f9552d263c86298b41f626c71ed2d9aa5dbf729d8c70c86e1149c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9f0dffe8fbbb2758eadda830e06e5ad86b3e04c097ac6e9a71b363799f7d0aeb85a3e985281e67b36178f81b9d92aae7e493a9aa308031db2f96959ba6f6935443e5e8fb617d60ed47262af7deea6a5bebaac386f5612c8d57b058680eeab470c18149057b76dc657bd28da71f758c2514bb3ca986b6eb6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cb8111e60854c7887e7e893070dc1898e98ed3e5641b0a36c33166c35e38c422566153a1175f6f76f21665fabf6b53c32efa06ecada8b8dd5d05e5a2957db35214b6a41a433ad033689a812aff4536667e32a3705dd2bf75a1010d5aa5c3833882180cf6505405385359f4d29598c5c79bcd32fc0297f08;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6bf299837760a89dd5e0e412e3927c6c9ea44ba141bcfd9fc3cd72602f5a7810ec8f604852ebc3d3e7f6d116204699cbd22090849871253f1f1b2e7dbdef7f64b7a974167197c7077df43cd3ee9972bdb241cdb3459aa742402be2c38cc33fa7310fd563cc0b57d2676893be40e8eb3704b6874e22f9b76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc08f433f19dfea4c435809aaa9cdf9d8732bd3cd51b8e033c43bb1bcb668565cd408508aebd4989b12ece7272197429ab4e7788db539b1c1bbceaa546e4bf127d0d10e8750c7cca682abe8c597d9a17ab74c886f33e73b57780a86a3343d25b82e828410b181c4cd8b3edf2639a1fa59b027dbea4da024bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9d462143ab3030224e651d51b80909e6f6acaca2ab69b2d368dac0c7b8a6de88862fa2f849fb2a4c2e19aa03dcb0577ba33829223179f11712b97b28632220e4ede9868076601742a157540e2397586dbfd5e19a485f3e287e755ac1ca32a57817541a8c8802409297478786b9be5bf905e2ad6dbc68cb0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb97775e6436b39c580cad7e66eb9e92c5ef6542ad1c83839791c58041541fac0fb806c80fb5bb4eedd71b1053cb5ea57f68166c96c17e5fcbf2ce26c946c978778dd88a328a3ee8bdd4ef71de445a3ae06849119eae442f35a1c28612bf55277deb2e29732afff5d5021c57ed0ad8945111694c35199bca4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc237525131298a2beedb1939a9a5e8ea3d46fa80b27447a07647e96bc0948ff7fd9bf985eb78495de0b8380e36ac9c9441c58f0d1135242ce5713c6de47b6735eb8b4ad3608a9f3ab8513b675715d9d217ce5f0da7d120487b2acc0d8435344f09e901cc920441cb55cac23ee1bc985b78c61eb956a414e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6551b06f4288afe1db18dfe04fb89f0ba8fe7dd17b2a52e209e32f61e9749d564214349759be3d64f4fe2858984217c277be45bc9a809e0a270c38ff7cc7cf98011693c7be29ece0572b18669e872727d16b4084e4f2d26bc542be012d64f0e91f147dfd66a3a2b16c9100f73e08e4ab2c88a97b5fd3ce5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b380f1441eac5b1050bb138f0079bced86db163056b62b5d346a52dce6b63787a20b0b25b351300f0f46ad885b7708560ed9f2fc03ec76afc9621560fd5500e77ecf6bc6513f6a8d646ff52693929a93cd2331f8121ca6243cc0b55f73d48e52f8108fc91a385299b480f214522d1b4daa50546255c87da8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70b43485d155900749a159574a9e149d6788b9f4f7e69baf0c26f1d6bb424caffe543d07cb99610736a08bde240bebae8102fc038acbdb56263b3a92799c5da33c6977591e0acd8107c9aa9db4faa8f4bae5e758d1e7cb2156a39ce1cb2471f567d08da37c4c35c1b5322022a5d8915644b259a4d33bdadf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f3948993bf87f4923d621133caf106ffd528f00fcf71e917f2ee705a632c70f5a903c5a562e34e1b0e9c87ecb2cbd1f18ad747b75259fa88823b6c6c0d43de40b983ac71f43cdedc3854fe99c64f97119e048b208cf0be4addd43c18326abdc9f18fa3c435d83cd01b9d248e7dc377eab39a1f8a2708c12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c0b848e07cac70680c708b0e30de1043be40c7ac1c53ddd566892c849c126fb44d45559636aeec97d55dd6140ea6f3cd81f0803b54726d3a998532ec04a9e5b8c93f22a2477fc92de5cfacc00084b848ca81d2f7a2bd70b040095dc0cb6c18dbc5b40db1dc1810d41a684a14cd202712b946e195329561a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168c08a28855228c399c3ce073f7bb4af1ceb0adebb67a485d68c907c6a30c47f64260bf771b205deada87f6eee7eac92016f90f7a4203384e3a40c989eeb69578d4c1233126735ce9e335eedf368090d265d2908d26337e8bd11a349113bbc8c76f518965e4b14b5e513d1b82d54bce7915f3eba20fd894e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9015076cfb0517295c708681ef21ab6494a9b2dc1458b7a1856c75c9839a0fe88505f05376eefa4f38f082ba4edc7edf04f32d91730d3a6b5ff4c301685c7501ddb9c6cf6137361fb0510b2c88c4ba3ed4b056accb1f7a80617d5d80bce9093857db47b8a358cb8b3b5caa91496e409191593a758485e939;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he0e736071f8b96ffe80adaa1d03f761bea01f59d416c1764e22a295d7650d9c358d89cb7b9ab8d842fbacfa5d8130aa57f432b5079ad9f021b5c021d96589c7515c9871b84682319f25e9ebec98ec5865251056bbbde65e7a4331dfa1f8ef01d1f9c85d310ee3245a239fb764d11495b271f54d144e6c505;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1438f11643796bd517f67312f96a16c063be77b3656c5669226a9fe364d4eee00c54a9e28906fdd9652c3988c21803efec0876d23c4b3b4d7a669cd47c57436d48a66f7f76c6c2183a479972e4c7352b60e22befcd6f904c727a6a0b41d2f72aefdd32ee672d6da8bdca31854787080ee7249055b78861415;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a20d152c643722d83e1d1f10afeeeb7a9e28c30649545d069e235a282e662e0e7a5d17d01b1eb38b82880219579c2e808e2797035adbe43d35262b092267074166f3fdf3733d05dbdab2e9c03920e2e7528c405c5f248aa3e3d6f0b1bdb962fe01086020d74bdcacad024e8c22eef250757ca322126316e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b543d8fa70d538ad492cc3d7076150ad908418ce407f44de2eb8cefcee933a55343ad0a4667c053924f8a6368b4d0133e55a1dda4be9d0d11e38a479a531ccceadd9126823065a4854615fcf0d65493f9bfbd2eeb023f87068afd22d1652de0dc178c77d4632a089b902808d29e071d59568e075b083d24;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h825fd81a38d9121306938c881bb0843822b04a81130de2fc4141a5676ea10a32a3f7bc0b4e5db36b8a09b3b05aa8d4e270680b71961ec59b453dedb6484510dfbde59a67dda4e95dd96b27626235f5ff1cc4c713954a7f8e82e2f59540c74cf24823df8d4c555fac6e3720eb382c5b491f18336c0a89dae5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a325907d25d39fa65ecbcd8d64ff4a01181d78fca252c6af9efc46a451b4662a968dd94ba06e736a688ca3c75e3d4ba10f6755334ee471ee09e918f72a51e279d74c7bbafe2a683eba6831aff97a7965f4012042587d75ccc54fda140e6b75a776f44d06f48260a9838a19f4b8d98189969d41b1a00cc672;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he599979e022910446a33e327164a6b284722c6da9a5bc38a6278ce26584eec3c33a6ad77c04e8b1669ef4fb5afd44865ef3993795a98c4314dde8a5cbd82733f2168ae76a71adafe61a3437ad5422d58778bd868c3e8f7f4a13877d1cce0adde4a5a9edbe0bb703cbdd9d7e57da498352e44f6e0866eafe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd774bf1abc628c51e1032017f41930ffab129cacf32fac6197a6daad9f43337b5fad90453400ec8b70605eda0e83c8e6340a2bf8f554b8550f42bc6077f88fccf631b168b3b620b9d2eabb0a21064580ffc9c5c01b35b9d5097ac5f9bb94b68d0a8aeb97115ca2c39742d5ed958127f8f1db8c2b110c035;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c72a8ef77d613759cf511b32de902bf079cc03c3a38dd05490c5e56fb854da7fd05722f93a7cdf67d3b2b85ad71866ae4fb7f011635b61dc2018da7048534734f9634253432ca08b1c017b6a26789faa1dd15bd7e165d178863bc209aa8acfa8b59bbbceef81a218cc94c5674d067c00525ed36b5fd1ef27;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c70c487295af402a8669d76bb833d7313b0fdc4501ff0a0e411553354903fc55298dfdfd219f3d725f12342cc8e12945e918f833111d44f539b16843281ed972aeb6f38a8117c4dc6147dcf57b5e558201d2ee31f3a0d5d975a7b4345fec78c80c321ac378aa51163a5073e83e444e04b78debc7a08ecef;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfe2ea9df53f2fb33d0c8ae61c381af1fd2606b1a119c87c6e05aec59c8f93799391ed83bf45baeb55e29a01a3ff6b6a2bdf163f5dc6f0418639643592b7e3c55d482784518fbc93623e18e6d9c488d3a0211ec63a5553f6eab181c5a50e3cbbf9ad7557e0eb714e324f3a68edfa79f88af5d2197265fb69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfecd8af53eaa9f803312bd9c8914c17b44ead7a4162f0b1fd4e007a91136a22bbecd688c2a745aecea4398bda12f258515134ab31c6779b17df4812c32557679af72fdc8f622775ab1c5c57acd9ec4b1fa4a16d78c68e302603d3e6186d96c95a739f11f419ef37cf734fca824772306f74ac2e3d66f689f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe5ce628224d3b300f72d1ae2e303418015d6d2a562859ffddf1a2cf497624a6558a4e178867022bedf64e6c078a06f78604e612bd6772ead574fd6787df5a8917fa0fb63901e5a610069f4f3fa4b54b2c65534adbace869b86222d75b8295d5fb46a62a351f65857365bc5015c35b1262944ee98841c3f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd91b0dc086b744db3202a434fa14212ec0d1a20b0b0c47c80fa1b41dd4f21729151860f6805e12ec0b90938d9eb16fbcb11e16a66ce6314ea49cd781dd35e90c6490ac91bc3497c899ff3b8b46d3d885df64ca75b4f74eddd8e6bb2b94ca2965018c45ec63199b3a8fb1d93fd428adc5e00b88c314a51d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5cdccd34efc47197d955d8a5c40966d0fc9169180a88cbec17a69d8c6ae9685b8e4f5615f9f051eac1f76965ba71b3d52dffe63c211e48e67972e8c441934c9fa829e018a63fb88711831db30857d2207b65d89bf6d9e8e31e38432072198e3883ad60b3b1e49779fd3cf579f37e3ce7405ffc439d057b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee1348c3af80495be2adf37e964fd34c5d326aae7cf72a6ff7557a15d29e66d8e444fa49aea2caf2b124da58a9d7abf4a106ab6ec3ff3459ac0ac9665267bcc8389f2214ebe8c4edd94de923a1af50e0f095d7c91d64b2bd15873a2257a2b2e214f88caa33dda304c06f92937f87da6b63c32954fe3fd848;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138a4367f4e37cbd6ba6614abe9de567be3f24ec944f1946ba3526614e42766fc94fae0bac9df184e1ce5c93d61a212ae2b724d80cbf57f04a2ee41e317138928636609b469b84fb4fc8070ce6770466045fe98cebcbd0162d759ccd6ded2198d67dc76199577189811352977c5551732c78e0c0d63e2d4cc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45ba4a5072995c0f68ef6438072b608526a1e92b0a544332d0613e159cfcbb18c8995dee06f491a6af9985926b042e03c5350bc5e1861e2516a1917de89970dd545e48eca16f8f3a982a45e3e066c43892971246d9190ac64154534e7a993ec73bd850e82ea6df04342d9f6e7927bfbba7fc8f74e98da312;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb70df7900ab31608cbfb15e868a27ab3fc17a8c20f6eb9bb405a0aeab0b98e3ed79e595c320e6ab030a551fa245a1c1585518edff603b7f8af03bb8117fca6b66e75d9a23e2d73fc11fb9ff2706fae7dae64a3efc2191ec02c65b1c6c7d87516419695ff59e267dd0cd40b665e3eb76f6178cab500b573cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bda4eb013bde367e218237fa6505bf4de25cf57b1c0db2898227f80aa86e2e4705b169dd068b338af5704ba73907a51063edfd924a36e191b0465c081695aae7fcf6a1205c3cd04422700d60b4427d6c1f77d003e5bba33c5b5f7c6421a7dac19a81070ffaf00364e0613783c0ae938366819b1725a5da2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc5a52da93e27734def13a7d2ac8488b2071d2eeeedf56a1b043fa5794b5a10cba9f424c298697750762cbb3de4ab7f5def3dc5c6e43e4333161982b96fd15163741dea14e17434ed8ef559570eae56dcf16aaa823a77eb6542d95a6d2c38608345108df4e3d359d05f8af5b6fce9ff291586803dac9015e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6f8e91540f5b883241141272f3ead6c03614fb68ee3201add690043cfa783d370be8db0c7a03c3480aded0e945e5f8c6d99f865c5ea68db45c80f861f9b8a082dcf0c217bf7a57a064cf54494a1c2a3926f525f90852ffc9919f48f583d840a2b78d64e2ef30b7b27f4019d97b7b8d4e2205dc044b15c00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10488232fbcdd033beb2ff8bd5219723dda0ae1dda4ab4eb197f7721844fc1e99fbdceae9c7c873c272d48b6f537e49fa474f27431f74d16aecc66e917b1f6df640a87b55628c3d5dcd0fc5db96a16e7ab4fd5bb6e7390d9087e8b21f61c1a46eceeece2693f140c6b668a70d885d11c0ad19b936e28442d4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166ced9f25457f7867ac03c5d172e861e922469c0181cf319fc970b3b3fb4e23d259a66841dbf896d1aa0420ffc8d266d21ca36814bc70eba98dbc2fb8d060045aaa4bbcfada29e5c057210c7900df3a155c83e3741e4a581c097ef6f6becd461061310c02daad04874071687dcc7c21c0355b2566200693e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3662c383eb4b34a221b753804abc83fec510c8b39c6b7e2790ba9f54061c8997d64075becaacf0d2b83b81aee72c659cf25234af014ecb9dad05eba0ee621837fd736ab7ea062d2132523ab141cb61ee6011d7c6e911c848121084d063ec2ad8b65268d787298c855444306928122c056e7c20628410599f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23c8fe319f2d1b21dcb9cf4d8760ab990ed5dcf7f91a534d4d6a302500d631b349b8b3701c441d84f269e18d923947611c03e0e80aac2a776b7449cfee6388e7004e61bf48f603f2c98b74d868a0b8650861c3b66101efb85e450ce32135c792d7b48d5284b2b1ae055e9931d55e210eda2ad9fe26725f46;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196ed12ae9f27efdfaf7e06f397863da39eb2707d62983dff8682d23677ceafa165ab613b0a4106cbe334fa4a73e0ee1c1f7d61a889f3c3475fc07e9102c2bdeb224c05e2b959a6c9a58506013c53d81a0b33fd46feea7c2faced4c277b5a59a15ec51be153553cccfaa556111dbb5b74b4f0802cee0a9780;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de9354336b89cc6ede96f0c19232d986ef02f3351a58a4ac6447baa79dea2ca2b0892251233b76fc12838b8f59fa7a724b1f6a7e4fcf6c4ebdb54cf56a52a396cd26e9a602d9f29b8800d884beae7b47b65d403c8383931dae1c1a7917a21f7f97a61edba2ac10093caed2c7eeed54ccb2728bd74efd1976;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d798009d6b4f2ab165276348d7910defcb6bf8525b195897cfcbed02c3f0191ebfaa6277c43c3c73dcd758f449f08507a26ac881696756441bf6e0901001df5272196a583084aaef5c1fcea31f1bea6c9a4bc78fe91d50aeb3440f17202a0ee8030cdb7d036c5939ac8b2091283ebe18b49908569ca3f33;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1370fbd1dd2d0e4156289dcb4a17c78d0553ba4e173c1ba71c8677d27774d93d9f08713a03772759cc18a11b64ff1228dab9ba09f592cef288d4dc92d3ef3bc388cf45bf8af2cd051886ed643c282aa8b32a29c9c8b180f464a3a2165d480eb6a53e00dded66ec011c584ee2918d868b7c114e60a50abb62f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5392491f729215b0defbc254dce415e336500ce4ab101b2334153f1a5208815e5280ec74676aa42b578aa656fffab5135b7a229a1293605de89528d853f262b7ddf072f34c20e7be1db7980f1684419d559f29f4721e857df7b93762f102230cb3d29ac27465248e2e87e162e15bb45d99b8984ab8de580;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50ce2b1cc6501beabce6b9496dbc48913f13d801ad30c7af0b18f2ea1c2647ed1bcbfc4a8eaee0ced128c557fffbd4abc7399e487df9ad9b065613c2ed9e3d15924d2ce46f9fc9381fcc0800cbb11bdf6cf2c66da65daa1c7345632a7ea41439ce09cb759e61930a09721151ff58c50bd724f8d0b6c204d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h403385665f5cbec0bcc00448b9fb9750179c9db82274f6d97e350cf416d6e49a7844101096382b93d451eabe5be2266fbf569cb5ed09536410b92193a8857d9a66c735e92836218e71efe76afb1a6a4def23226ea9c3f7f4ae00387b5414cdfa910bb70f9407a1ce1eb541c77205f5785ff4c63fa6c669f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aba55d49f576209a619e596dc05e9a35364a4ced67227f812dd24ada30cceee3421da8eed39dde84075738d53855124294fd1a5e838e0975a9c37f6e84a008e17fc55768dcb3ed9b30c8e5c397ddc9a07601ec9dd744512a41d351713bce628c726d83d114360bdb940d65cf2219c7dddd1e05c2a2180076;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e62921fb8b674c5ec6c26ca9b46c4015901b3e09232e33357250d92e3fbb9fbd854a97222f3e8c135ee719d452db813d721db11d54a229bf3dad16177f2f54834b23ce47185f74329bfa6df689ff6a9dcb1b9e5f1004993bbc9d4d911b0d8a673e777e98b0479b4db474fb260b89c6cb79bb55165da2d357;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19683ad4677e4438268dbed6ea1272474040893fd82356adbeb40f8fba0a333a52e5c87d82fd24874b0311e443ecfd60e0bbc05984f6f8c8e1bee36cd168695dfe97a651e5a3acbb93c030dcfa06874b21d0f6492c5408dfa72c013ece804caa66d5730be3618200ecc15ab581065bb2c491f838e3d61e9b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b27d263801c6e9e543653187481fca3b7b69c5fcbad3880a43842b800b78cb4300a7479035b3c9d001ea35e926d3a37ac6530c6faac153f5c0d906309aae31141e0e5d172832602d4698f1faa191cc1e2e61ba7f8bdc25891479c8125360785a945914bcfeabb51231be0a610468bff3af7637a76b84ce0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4626ac1c4c5807a26c7ccc35c8e2c88a6271138c6e4b9ccffeebbc588fabe935f6a090312663fa078a45a09b87d72b67af5bb86e41a5ebe9bb7234abcccaaa38a73157224cc670a51dead82827e7b8023a021547defcac60ff772b357850b052db8edc99e622e8c962737996f1a5ca11406c0c9b29237bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ab2008e4a83054fdca444c80b57c00330474a6c6ce17f69d2162ff963b591bbba29b2941eec232f25d377905b40cfa3da69b7479b4db0183a2c9f536eba6605ed09c1132b4991a4914665801011aa630b5c3eed2f7c41503c53f868c5352151624fa4621a18f9d1be40b087a11562c77c2b967435ff97a0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5826ecb95cb02179eb7cf5de0d6be626bbb5d637e54d5315dbcb5158434f612de87da1ae90e47724c1500ead2ff921a5c2ddcff6d82d128eb877ac04febc7c5c33def317f8842ea62eda5bbbc7cfe08d199e015a1cdba9d2a56feb98a2bb435da02f8847093c4f284539ef701b3167c589ac2711e566c1eb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf14d11f9484558a2a68629cf3100ba59d41762f3b78f4b5b896778081792f4c0595af7c9c2d6df5b72af861ab22f7e1f6ad10b3303fd7db3ca11ba540df494efc5dc27a305717fac5ff8038707364351379b48780cf383c3d7945ad17c4c57a2026676b3f4a7e7bb6568ffedd3e47bddbd4d10e402ee28b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebfd4528d26ebf0c4ab4b08e863a44eb58c58ed2224218c540325d625bd919125404e6d93e57255e0f19e85ad936308fab1e485da87f41d5415787c960d37e1b21a5aa129a826e050bedbfc627cc436420a7cab71f261cb5a280c13c8ce76314cbe69abf97e493943493c933bba6ebdf480ba0b249758af4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60031b70bb7d8f52ae2a6610ebc47d1a779fe3c4841bd5728beddf58524f7033fc046d337d0777bbf2873ed1d6cc7184558309cf19b851701d4030245654c7aa68e54776a73f2f7617e43a8ba7dca9808d55531958891a125df2f48f3497afce95141714e03555014ce046834986bb6983ebadf3847f3668;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c732bc041b9825e794323392f50993f80d2b9e0d1d970a9dd00fb500500f1ab9782fe78c4a8dc7478ebd964e4b925ee044f79f57862290ddf1531b7c943d36e2956848048049f83065516d5f326e3447145c6c624a4b5c108c3f0893e042e659961dbbc012e8a78089d5abd6475fb6f7bb941c946ceec5b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68a78f815bc963f2b2b625a4c4b31bbc26f03cc1bda0e93adfddab7600f3351d77206b1fc6b7fa9f550cdbe7e115724f7290f7d950e2a5da6c0a77a5d513965155294c62c74185478a672f59e81b10ef0ef96c9c3be0c9714fe196629713f740372829530aee196f6eb006fd446dcc593c996d417891343f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108ff6440a373eb5fa5ae3ea58219b7d5a6dd66e2b38ab9b9ddff0d8beb9ef4b4ca14c2041c4dbcf36d675ab6c9225a082274df6bac054e92bab641ca48b373db44d392564c10193a83fb6989101b6d3b7ecf43434495ae868b470ec1cc1b16ea9e35f5f17fc96886793651009cb369f6f58ee8f6765ea425;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8a31ade4b2b2721d7f6d5b5a9bbbb8e10d93a49869ac0425e635888e0b4b2133ad2b27de6fad59b011401ea79328f507a01d20100af5c4ec47b2f117a2ef13075a8be4cc53d733ca66941608082ab9361a74425ffa0513769bf6845bb28d8e5894f184de72ddf8925771844b5e2946f89129ed4e9c82d9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1180230e885f4e5fa861c960ee46152d615004387a02ddb8d954e4596c2675198f1c92a495443ce6077ee8fc94ddba82231d5008855ce0a51dd93754a50a606d95fbc111a9f276e56a47d2bde1de2f7583ef0e2231b6618222fbcc74eafcf911416f6e25bc3433ef304648250a677952d0fbf40c6f412c351;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1987d289473d2d7cc3e9eb259b0b287b940465e6a62481e725660cecf5205df6c6735c9610e4c413e40d0ecb9d83bf4705f02be2fd141cd45ff9e989776d48b1d192b8bd136257f82343a67109dda211edeb44e5bd9be9d25c64d84d40a93ec044a83e2603ad2d9453a725032ebb90772159c7b4c975c63d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6b5604aa3ca8dec6d12b5e3fe6139035891fb0340c997057b4e6aedf5e212af2d3549108af0635f5c078424a71f38d1b9dd15588d9e6ccf9c0cca9e0a421409242cf98501b43346e7fd99dbd2fc88dbada903b9d93639bfef80f039fd1f5572499f96c3d7eda1997b94c8b1587ee2062ed2a039de835f64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1feed333229f36599b8611f8f3593b838a7d34061e43ff35a0575820df0a4e5786f81ff89fe160f2163bae55ddf5087e19414737345f6932e22931719851d49f303fda33d0a76afab513cd291cf5ddc4ccd1ea7635cb820013b6beccd42e28007503eaf4644432d5ac714d88f298adf87ebb7cf3032111212;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5564f14d5b667bdc5c8f75d5c0348aab873d2e0c49bac154498e8266468dfa5e6dbb77bd147dc2f6511e87d50be93b89a1e3e652cedeee57b00888a114e962a5c448465cf904481d3c6a50394b1248366f81e5f33e53c8761fd43723f798b8bb2954f894a5e0803dda5a4595430e450501ee8b513c31193c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad0a161b423ad6492b65d6ccf23ac53768836ded671c2ac7db494ea17573b34f4bdebd089641cb2ad22072541b049ac0c2cfbfb518b1663788ac2993ae59fccd7307b76e265281e27b07ea1dfa31ae38fb6a33492d7cfdf5c04cd9e4510d1ae9c34c5a8b099e3f9199aad6f168a898cb6d75e504488ad0e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha282038bf1ab8ff4267e5ac98063b95629bca810f2f80158e014bbd37472a267dc7c0a4b61d3bdca2cd26ef61fa1d10fe5219a6c74e6bd132562a7b17db52fd0219dd8518ec8a8bab0eebf6f5f878972b9b6976861c0bf74ab45479b0bb2205a9af96efc7cd0022259ea0ac305a570c32d6ff934a4152f97;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6739fa260658e112ce239557b566dc1e9d6d7fae55487c5ac736b277c78fd43b1698ed7da7a44508af1fb731e2cf8f7ee9fbd41fdc5f84c90a1243983001732cfa57b42499e85f8682f89aae09b73a648dee320b5cd3653f3e5af1cf6af6372f009de5b812b866cc1f0c78d84d2081315392a9fb35a078e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16817d2a1d9bd4fd719c1d81c9dc113ff65b4aa20ed57f077edcccbcdb03af3c440c09c8b29bd4843f7789234cd4412d8b95fbd9302a81a1de4421c1d5b100659a0e91bfc538caf0c4ae33a2c2481506afeabba2c71f1a62306807e09ac176ef4d101bc5cc652a017b74b79674ab4551b02bc667a21538a57;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19bab63fcd313c98264259a8f710a1a3d6bf1a6d9cd2c504892906b308919adb238e9ce2363b7146d1ed9786cd52889f6ac2eef17ae811c67f5a49e8708a771fb08d927b7e390546038e9e27b038a3339bb5a750f034381b816be3d911a24b916642e4543217e65ba4c95206c458813b1e6c7c64654637834;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d3f68f8436e690e2fa6f6e6e0a560fc2e71f7d7d0f8c2fb66ffa095f254c3402a21971ce7c4bf64560035cd4e93371892c3850033ae81967c84154cb36a31c0f46be55f325f8c2cdcd63ff7f5e29c8ff12091f06aa7fab6eae91936e6e93368ab2225c1eba32a969bab0a28e2469b87cc32c8399c938cc6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127870df20dca5e839a25c1375bce952f6ec73f5cd0528556237b7034fd9271ff01f47734dab57eb4236fe8b572ee32bff59f97a45c5bf9256df22c5815e8e646f2e775cf2a4a48cbe5c35d5e42d04d47a4cb3137af60e1d70f4514168210d687345030f82f9aff8823cc41bba7d0c8b8a7489b3b106375c7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1661d7773d3d1baebabe6a3ef0d00c0ecb9175d6ba11ffc488d4eb76a7314e0912dab6f811647ad74a37734157a5b37691bc6defeeadf9b1236dd65b982ff093374438b00a0af19f72492e56ebd30f939fcf2b2c814a5c7fe9159277663c3f778bafb3d20e87c95cf46f190f4577cb758b55c3f92c233110e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1acf3de44d34171380cddfb1fe99563c5cd63480885314ab05c9e8dd2112b13e8418eef73f68bdc04f12616a6fea3ccbf3c2e0e538653cc611fb3a16cf2ad4a8a7bb49f29fa89bc575d2690742d93f2bb6a0b8ea67d1107cb27fa1a1beea73065566191f27cae98ebe40441b5cd33180ac2afebfeaf12406f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b7a20e00f859e546b5b9c3663c0242a8057ad0a385b68d18b4c07d968b900bb712d86ffb0ac2e1709fbe82d2a93d32076fad3c9f90209eca1f808809b1717c28668f6a1777237e11893452b90a6e36a1157d5eecacfb386e4691ea0b297137dd03f38ac31a04ee2c7e78bd0f88e297df86ee34364856e5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5fcb9e68f9975311f9c531ad79b97152d3539dd5dd9c131e705fc618175b1eae066c1f2265373e19661b95403a6634faa492cf99abe5d414004a0157d3c1b29bae3c3c1d989f7280e8dcac5f96cb1ed60294c3705d78b11a7863caa148c897dea1a53f9d2b1fb1ef3917af6a3a80824ec1bc1c9bcbc92650;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1b9460d20decf6317e043a2dd6ea3132a17c4e588820932c6e79108633f70055078c51e86fdad541f5e8608ddcf67719f09c06856d6fb2c727394c323820f818013445f652dc010ec6b66a1363f19198cb1896acb9f7893d44cfd9fdbacba0e18123bd0d64f6da68301a1d2354af41cfa67c443f8c3f27;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17671887475aff0a444ba74ebfbc4df6c2a2934f89e42a5c83ae082fa8ab738c0b3ad32825cc7f825a085c57fc6b9330007ef3d0a6e82f4d69276f702391537ad112a80783326e6afcfded14f9b427de830d7f996db30e451ce8d4d17ee03ebd7bbf1637a080a7c3979034d57999df1aa4b4868828ee9a9e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h990de44b1412c2c834cb469e414ebb61349d130777e7d10f2afbb53a7de6b1e218c11595e3f5bb7bac383d09d2c8e13044cec884fccd52bc01bfc6e57b46c1faab9aa2a58993d88093a435bb5a24a0f63cb5e17b0f4a31abb4f36dc1ded4c3061d68a0920034ab38f802b90658bf55a400ba46062808c1f4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e4fdf3a471b32220b90bf13666a26d272408cf8254be9d5ddc1736947a2f8de826bf2c13d8e06e21ac8227a6a72f43ac3399b5d4ea6c469916779253615596cf67d8056e5e87ca83f219f6c019f464c86520411f4661adef9b6c4215fa248b20226fe40756d5fcf059de0c4e4adcf87d0c6c574dd010a66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d0c458d9ddb83578e3d5f24958c79cd0a8d5881e92f47a4486a62a15b569c532fbeaf9758466e5844c2aec86f6edfeb8e16080a07687d38c824bd909263fc7940e8e658d24d7849e07cca5cd7279b151030525d2dd2e72425df492a68279c10a2812143794c280af8be84542563ab6a51cb3d527d8e1b4c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1481e7cbece52e2400fa8eef91bd58463745f085d7db59c24094fbf5017da5a36100c2e2a95de0aba204f043d5d1130d8e6215e5397b0e4d110b9d034d74e2e06389ead73f88fd284c113878e9184b9072969680865b8de5eccd43e34ab3948f36bad115cb010de973e51480543aea7a27b103e7e57f7beac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heae9b5c73f5cd8881d1e7be9e9d3ebcb67eea767d7a431c5d4900a0f4cc36204971fad0bf1ae725c0aa5b6e59aecf1cb09c02039d31a1df6df6475eb2ec3b366e3146019ff998b70e0dc1ab6c1afe2d75610866b638d36a43aad3fc650041a409b2608311d8dd428d499dcd8d9e9c247e0974b96ab95b716;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c768717d7d4a9c98bda01a3909ed328e216b55671e79e289c1e2a943ecd383a5b995f32dd331b7cdcd9c1fbc2e2a75861a69e905208a7b48a405e73a04b509027e807cbaa4a0be0e0f0f42aaa13ff5f86be4ed803e6e6cc589271cd5833b3cdce1628c048ea08d3d8ddd5c153b9d90c96822a0ead267f83b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cf250d7bb7faadb5de1545591af1f654451485fcf8a6c74041353f3ea772c26e5348f474a412f93d69cc435fec437b2b7f54911b91a643a2f1d8339c0f9919a3c163440f459fe40a411484278731c08786f96d01763c1ffe67ddf0cb722f6c702f2209f81abcc8f4a6b67c5be2abaab22705c9f6dc13600;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h798142efe32eaad708fa8ec9d5283ea508490caffca28b8b4ef4060baabc66bdfb7a4995e42640007d0535bb1551b2b4f57c23d405faf2749f2f75fdb918cf4b2545d60d4df1c304d104a2485a3da6d9bf6d2bafd643192c1c5e280936b7eb8fda2fb1b093d5e31c74292e29e7324a69bc873620f239c1a5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46bee2182cab2de735daa618f33e489b74ff45d37888009e04dd34a16050628c61f2de9043f66af5c61d491f712274eede27727c632eabb60ca68a5119e2f2ada07e575226f84f26637c9eafd5deca568c07cc5e4cb6ee419d5b4bf26384292556dfa1c016816d592b9a8f6914e3d088a42573344e15d6d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5523ab7ea453a46a4516516314fec90f4bac76478a285ec36ee4b135be0dceb1747cf7c35e3651d94e2355eab0471b88b54f79f4ed166eeecc6a455030b5d4d3a4fb02fd6f3508270335c3a4fc36ab12d22d308dd5001790a417f598d2678c9baef23697630872b6c30fc1cc6f1173054ddbcf6e3160f3e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74a830077cdad80e98870ad446ac0375ccc0d08c6c63b42970731a6db7990b2b9f900abc5e422688512cc387fbc8c48b08fdd9116a244a5354f8d5a1a283a6a8482dc3468db19ae8a9d0515dec5b5353d1d52a715c475d8251cdbf1be0481ac2e56d0a85d13eb1948f0382c887a32e3e195f25b1c89fb996;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd61e07c494c5d5ca3452aefaec07330d09be31c8b832d2d793bc048dd38346047405ba5bce594cc5380c86cbea9245c4ece8063ec53501330c0aee739ee9ac98c4b0fe0f894984d464b9f366849636400792655ea6132e9426950afc718caeba2d1644129d6e03e8d04f8f70ece0358befcda7b9194f49d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac42c423b6e74253773fe9643b787cb48a34968035a25c543814b958d18f5005182bae75fb8a0318b98de9a2e244e3c85734b7d8cb7e4b2cc6409c6f71edbcbf2ef2219f6d4036a5aab9f53af2f2fc7f0c4a0d32c4904ebe057a61f4a953ab801607395fdce41e8d059763d1219e586131b49e3e2e7eed12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdeb573ba834c080781598876803c235ee928df4229d514bb82c930f80c341e8ee24cb43be2f2df38063f0c7d96304fd5db4ea6f0883c046454287ba2099e12d60b481b5eb62083ff71c7b729879a50f07e7eaedcafd3ba3af887b4a1554d2ce6a17ed8163e94bb174fd7b4b551fdb0825a18060624da4eec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7fe84a08f8a2bfc0285fcb562c5c074bcf5766c2a59bf6b141da6040d3683b4fe8fb176a9395521651e3de7f742bb1e01f53836ebc8d6ea0718271e079fb4a38e3772ec030ea46a263fd832c66749b6a63597d400f1de474f29cfddd56cc100872d52e7b2aa7053f013411f1d079d4a622f485a64fe3d05f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189143b94f7226ced8d6c8326db47d55d648e8ef03138a05a8f92ec4780cbba6e06c9521e564ded1004fdf32f89be620c39a8767a3320e6ed381dae54604d3a3a91213ea46a06c3e6ddf746bf9546330508d177ea1617fc47195ab07e57aea670593e3360e92193dff8e98fc5ad2171c05b0546bcddd71d2c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heeda02c9f21d426cadde062e1a0c25480638d538dc5cdd1c9a1597e59c0ba8d88deaf102b033727b043576779464ae6dcb7893fe5a931e29438160d8dcca3c58e29ac2c91bc96173e24bb485cf6068bcd42230af8ca7f39beb12a570200e6ceb1fa2a3384028fb92adfc2542508780e3da7dbdef4746377e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1689fe12f681b91f2cfec6c2652f83fa9c019a7ae744e80ccc52860d8f9c7184e05caf7b9f018365f08b7e9998a9e4c6eb2345594f2aa4329e85be2e6e04a49adc9eb717a11fb9b3311f28832b05818e7858c13b692678e03d4847a545f0c634aa55a5041beb58f2d94f258a64093f838c12f40080fb5d46c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22451e8ce231429afd46508c031605d071a1052398f23ea061c7f1da22d43dd81730b06e0c39919f13122216bb86d0bd01de98ef0dc1fff040aa5e7bb64330989b0ea207c14fd593f75016f7e1e20326521e2a88c4a577429d40f2ff7d980cb58f42fec817fe54f880eec35d612a77b95d1a370da2162313;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52d81ee92f18c3f9e8676289f723fa961bd69a97ab811fdcb7d3b08850697c22f81826dc0522453d798c5059e0fa869e11469b6f0f2fa16b485907f24592dc341507b48ff768242427faee8530b08bfc68d39d1e62859ae49d83c92749133f46eb14d4f2a84ff547600d733d6280124a667c11561d51432f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cc40479bf22ef0e9b783a597402992455456612eaa0a2e844d8304be62d156633694c312e689e6890c576dd5100b5e52b63a4cfa938b65fb6d51f1848ee38714bccca815334f3c14b0939ccd4e8fa6e8bd2bf9e8cabab64979439421bbaa5d69d36f035165e42915d937388f8070a7b26655b5afd1df33d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31be7a8b807717989e21ca60ad70f9cfed17829848f967444b91ce3c363e1d5ed2b980013e61bfbf11ec49684f4888536a98266414f55fd1d32c5d4d1e19aa2ec0d81963e947b0f4e6ed8d9487a1ce609637ddea1d85e7067b2330ff9e08102d81d43eea9a2b39f64ac53b2ed074836c3897e60a53ccf804;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h829332a689b99860e904bde2a0670f4c0d08959248a7d88d203fae702b54a63a34bfd18a74ef1fa15d253f429f45c13d2788f3a272a08c03f73840b2764c43f0d77a71e101285a4f081c3b11a57d99bcc66747c236900730508bd18150359aa9a254da6dfeaf9b9db7466fe614ee3086029cc637c8f4dc1a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c48fb750342ac1d2a0d0db022b72bbb04e4dc68a78e8b82f92feb2b93ca610902a4e20dcdfbd6c6068c7da826693409b0c2bd2bde29093f81525b2aadcb3e7877df681102fed4c69a52ab0660acfec6512fee9a77bcd2db52abac5272c63eddfd0ddb300ae1c52b415fe7ae04a89cf4f3c08f23d712bff56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7e394486c0076d8ee6b4454b1338747c5fac0060eeaf9135e67795e781443023609467bd7a1d2d1bc2756d7d2e990f489766b111e2d5de57aab98a6439aceb6ea2878e4de3dfec27077b617c3c429a44fb5800790de7f69a644ab4b53bca1c4b7ee1598742634f7245ffb6b9a6f06e7c59087973178c777;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c959bf2f1a54ac487cda575a58ca7544c3cbd15e3573307269982434d2daae2a383a1abf35d05dd59430b6e64fcfe2338960ab1b4d83c36e79235d32c47957f5a686383b2a15c9a394926a637c10e326d78e74b9af0d625130c981e1907afc9b4def928b5f08186fe1876d955c7faf4f405a031e73619f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h351434cea66991d67c85132edeeec5880f21c23a81ca54406dfbbbbcc6fe18eacb41030a29e7accd2d7717fafd8f6928e5808678d8c6c803ce071d08dbcdd0db48f77ca870c8e46d98d387fbaed70ebdf1d7ab11a541887385ab8aa8167a7d2a696b12a7da1839ee9b7a23a4f1b96db0c7f98bbb3b70da43;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1613cc9902b0d955cc6b99812d81adbefecd02e5d7adc26b9226d4127aae078c9ebe98e9950fa68237c6863a2e5e5544c3d9d6536f70507804d00d1d4f95462d36e90fdabfcc79c2e10cd2be0c88825d695ab8bf0657aab30b1584fba4d47b1e1582c9dda2126b171ea40d28e084dd6decb39660286189d23;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h716411d02a9f24c5278be125f8bb417609ff3548b7b8a47549608dbce144341e0e1886c2849d89784501cc12a9ef3eb9f3fcc9b13608f5730cf8360da368a7efeeffe20f45f1b4c4af833125d30b9b5f9d13c9d5f150ed429a497270dacb49ea59e9704f8b0a2804a4aa8c50756bea24def533107ba49734;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62ec0ffdad5f83765a598678b02d6dcbb1d7ed033b619ef855b96a2e437d6f8fecfb5929bf3b507c0f5812d867f8555217dc66d4480ef7592f28c6ee6b04a4b648fd82f029a7bb06cfbc71ef31a93030a4d9b0b68dddf14c0c4dcffec5ce882454a0a6950e8e9fe5d45599c8a99e4e6c726a0a0a9ff8a546;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbda9b92aa005f5a2f31940e1e379add1105a6b5a993bc487d59fdaae91b211a27d021c1767da91e90ab986775884826869fc4b38335b0337cc4267a37e5a141ee7e9ae2ac868d35128dc0e745a9a4da15fe46bf4151be325f96c168e9546d2d2a6dd42e39e0d5e0225b31e96b141cc9cda866ccb27c7f8b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf223e7ad8f044d0dbc16e509990421102cdd883e4692961951f75a29c4fdf23e364610d35af9ccee0097ac095fa8a2bdff960277a756b1b0365e5f77c770cc0028879ebf794ccf1d3f162dc00db9e93b5092f8c3e5ca6b4899ed51c1c037ac38ac68e80d0f0a50b5ebef2141bec487c86694b1cefdf652a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2318d0fc4143fbbf21f6b40f1b1ee716dd283d1e7f5803b22d0f7321ff1216fc36e187d4e24241614582f4369788b97275110094592d3f941b51efedbb89b44b8288c7c86d03210fbcfb1b8bca278361dd5c1d071fe87ef500ca8249ea8acd6caa409d63b85d0fc4e395065c5a21676f57e55597c2d55c06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h389aec35bc7488fab6aa063b9908ec517474b21577f56d4709ecdaa6388bf871d2b53503e459a1c92fef6c7fa91b588f698b86faa93ccb70316e650ddd61182fcac475dde68dd482d22f0524d26491ef93bedfd03447bfd14b7ffe16d91ab63abe26d6c1d1b4c66ca13d49ffcc19e2d2820600ce3ca343ec;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2598b3b6d5e541697825911b162ea986be8579ad248435685aba52d756e545afab47219f0c980da318d527eace784b7d544d7f3686deca4af4bef3e5e68f2e5d7564ec35c97edf1da02c37644d9107431a0c8f37e4dc664d7217e6c1bedaff4681d21a272e920099a9a590d437e9aed2c53ac72cbd2c5779;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec8924183352826c4548ae3331ea043c63d834920ba206b4b25d3c14ec1fb925b9238bc62e89e1eb7a8122655efc3e9c6e0b1e5507bc848e4e3697021c67454f4230edf6cc69b673a77827feee68d159c3baa7151e6b7bd3260a9a86c71b146af8d7875067b0e8bb8fb797b05c1e3b52a240e3ec8eeb7d52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c97177fa066640e8e8fb04e9852d3c9b140394a016c389474aa752a582e0eb5a076d0471817dbfd15d8d5614904123289ea4339eaefea18bd8f07b288a57b5d3a3c72019244a8f0445b2bee81df1602dcba73f6b0c5827f60dee6cd5100587ce2b6532c410c6907ec6c6a0edcdfec5e8f75354f805d71a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3e6cfd11698716d48156eeba963e0aac3b958018487bc4db1d615f19679058ce3759fbc07e88a22b7cffc7ed04066f8535405c44d94834e00910e92e40e4902b81149d1767ee1109292b431f1fbc3c76e6221429b27556c8c87bca3bdec6095f6fd2f1d40baeaf95b101f4592f00e481f03e40ee41d4ac0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7b8512c9749ba86444b6a2b1248964bb85f98e8b823c54801bd9150987bad64e6f36dfb7f28ed5f21003a6d16d394b80bbf8156559aca69f1960bb9c6553c8bf6d5a3f81cde8c11fdb062e5dacc21ea5687bd17d798434b86cb89a1f7041adf1da725c7db6423cb0b0d10711ed32163aeb57b8b3e4fa2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e49bb64c46bc4b8c34c516e9640402a1879789e19bd7f5011c9930e2769c11bdc8d23c7d955bab280cce12d604c6a6775d32e690e9bd10954e722cdee637584398fd856df6bdc7fcc9a64bcec46d7f8f36300d48ece3fa2a1b9e54b6019bfffe89172cc057078b336a7a3c14dc7d252f3648100b6936d1b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146908bea3596c41d176970bc72b5c5bb6a807d3f603062085afc1d8955087c91cca30a5a7f704582ee50be58605c184d624ad6ae22a82700acd342ec189c9666f169c88c92a48f476c5deaab4762cc76fe1b3b17d567bd81193483c3b57722de24c09ea7e64b5b917add3044abaa1b072a3c8dc3232d55a1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dce2a3a8701e89abf499824e9c1ad3a68a9d52b8a0b357365d9223696a05d1733829989dc049ffd838c707a4e3d91b2bd6b6315c7751abbe02e93f9ff88689a292e6f362b378b52f2fd2621c59fc0d03d3504d906177eb2d271403ff692ba37e988ebcb8de90534804aaf7b8cdf1a5a62e936315695eb76;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8cdd45c91e1790f7fa3d7b4af70ed68cf0d2a293f0318dcb230cce5872624d1c5b96ed63fd93571e73e38024b7cd0f118c28760d0e5d574a6da090b6f1b5e9eb4b0d6136245b056b707613c1a79042aa72de19894ca058af61964a025e93b41bcd33d901dd1537c2ccd62354b46f6f9de7f86c5fe9725d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h859e60e760aedd27e51ed2e6d2a472e170944e37565e4073dc3cb0c918dd56e8e6d3d5de363d393a2ee64d74dda7cc2860b486b706634f764bfb58a2205595d92e5efab87f48a2af8c5856be4574a2c2e428d2ff36fdd884169e9910db31d08a4fb52cca5f12df1b028d1abaaca46c08b53ff0c8a6f93b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cd81993f47755ae8a92170315dda8f6c9ffdc273a7027f1d031fdb47efe5ef5b2c656a27759855ce0f7e479cf9477ea5e376a7ad4aebbe62a2c3650f56a3914dcb62a3094375516dd67cce6973555543f2f2e4d5c6af7e5ee72a6d20b3bbd257ce5d556c9b01ec466fa179c4cf408ceb1fa2506a303bc2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100744a60414c71547fd06ca5ce8d0d6440c5735870401d44fbf1d7797d856d4fc38b32f34a56f1fe4d5c32a3b005bec490fd4c93f2d42976bc2ee82367ba3e098bd40eda073dbe638f1a9cbde26a43fd22181570af122d4846bb6cc814567f1d57e02c48ecfed0cee1b5e02a7c0505c02fa35887473f8260;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196bb6f5c5701a8b8a507f0f608cdaaa1a719a61244daa93501f6b06ca5574568dfb29ec13015a2e37eb8cebbc2a135760c89f4c70457f1e598d96619fbffde52763fc031deffd700e68232e0bcbd9ee83176900954188568cb85a982a40bda9a2f6bd313502667751851b56ee9cdb21f9784092f2ab3a298;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151ef499e8e591111c33e777d39ce9cba9c3a085ed51bdd192fe8eb28f7172274c5dc3f0076b744677c0d33b774193f871afda5ca7caea7a087f285b6a5183435c0db93b85b1429ed0dc02b16b3e0a5fe2e62606dabde851f6bb9fda0f2b3c6273daebbe35f861013cc2e18e79c0d9edf46a17b423e3a6b10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4d63848d04c8ec309b5c1c21c224ece8b3d43b22999e4cea5cd36e973acc8e3c60f6c0ac2c75ecd3b00730fc5fdbb1ca301bcef5bdcc266da3f5bacc41d28056ca6c1b3821e380b3e554e5d8a0697b61220bab766e29ece418cff1e2e89adfd8f3d867dcbd1995964ffd071926157e3c1163109078c4283;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1553ef8bc63ff4f2f4cd322234c513d89216e01a459d8752a0e8b9f4983f4836bf2cef0ec7e3689e7d88f30c9da55f53baec8da247b6b4a406f36ea98455024d5c3c8ebda1766d13e78d042de0becab837a548792acdb31ad411714b89c5843e95211578daadd3b8fb7b3e45c28a1cd8a836f1057cf8d46fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1044dc791a9e92e2c305c5d5a905f732426a638d95e0a774388c58efc12a7e057ffea928048143318cdfdcedbf4969413676b5d86e64baabf863e59043cfbed3d3ab28aa620bed171f8d8c8ae474f398f54f01cd3c6af7a54fe52b52d1def017e952a81124e2510928d0d52129ebb995a17c4b2d13a8a9f96;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17105845adc75fb235392eabe4be3f03cccc2391f86ea4c9e09fc8282ff28d171d23751e945f4287c318e14db16689f9dfe3bc5260467462b060d61898feee3d6b6f5d17f519cfeac55895268ed189bc0cf859550d8f17f467b2b4b5e7b1a5d1fc2c00e629296aad4f8a7a06ce95ecadda602a5d950cb0ca5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb85a84b81b69a7efcba5c1da9c1a074ebbab95bac317ff1d12bfeaffa8f429d90eca1fd645da47bb2eae239cf4f5ed48d060f50d8ad5a5dcda4493801a625c2c431fb65d1e06c2488e497e5f3ffd0aef9ff3199ab041e3bc0850b9dd5a0ad190713c7d1d54726a84fbfdc8b8e8b00bbb48c8bc5a6baac89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc783e1587a5fa70298b3dcd8eab0498e187bf5542145e0fd98c0a0b9f0c2292403ff5dfe6907360646ea1abec436f3f8a6bb759c91999a5414f361c05b3e200dd41e71fdee0e1b80e54356e299e57c45845561eaa08d43f7abcdaa5dd8950990f904c8c50797b61bfbf60241f5c29e3a319be303e61986b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b7e920a876c2d3dc4590a51c3df332c31bf7ab44dc03cefe64c193431a55df871a5ca63d75b39aad68f1adeb07ff28980f907d334a6feb73cd7b33a4735920f9034bf4b4fd88bc6e8e04cdc966e9f2b403c25023d6755360ada227d8d2f9e02063edc3ba15565562c2e312d6491586e4217437d43f8b846;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1152b1bbf16c619aa872f6d8ee0b745f3881fb2fb550f415f92ec90e096443adfb98072c6e449933bdcec0200d0f485d95e7c395b8a452059e79224cad52878d1550b25fadaf00da5fa79b9b99a3b49d95bab90fc49640f81c20ebffcda308ffc27d30dae01b6961d84b37fd911554c202be9b50566c2de94;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1918e37b5fa39d611284adf8f891ee66771ecd6db46ae8f2992e403a427fe5336d01b7105ce98f13256a912a18e6c6392ec9d55e23c8b1f122ae21d9a71eac6ad34de2bdf0b647ac7526cd98305745853e69814c54c188acec74745e9c7da81c1fcaefdf1b6abafb648c9b948b8b749df778548ffe8602b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75af86fda90e465c99cd09ae49cf49fe72ee44d515f8134ad9a6f1752e553a3188f4897ee42cf82602862b55aed39a590f1ee6978c5cab202348977a9934f8157f7a8ccfc96ece339c546e61340f0ffbf7d12dcf8029ae5f87494657f671b6fd39ffc7403897e7555f59388c9ae38748956693c19b55cc7f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf6fe0a042b19a6c492a35fe257fdd1c0346ce51f9cf018719be78129d33482a8f9c979392f9c2218fb13d6948d423d528a7e3a1d77e5c1d7473746d8c184323b2dbca0582bf77eef116f7ad0e0dd6246487c7c005c785cecb7df380701e7e2d70f0f22aee5231888ca1a19e5b39b70cb6d0fc3f9ad58278;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31d3c39e87e882d4da91ee1c684cbb678826cbeb64fbfd026ae23edd661847394f5864a8ef6e8247fb2f51e13cdf61d5921981835563d0708fee69e255a05994425a1951d7ff9fb0b6335af57f94c8b8d941bdbc0970cba3a14b8ba85bb3e62c9e561ccb5fa8f9b2532f03d179bfc06e81ad89ff4e170c91;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140c6948043bf560d337eb18406b2c245838464be58fa1d9759752b91c073463b0a72720c9fcbf6a7bd20cce6066dd355e2796f28ed21927323f68a54f329bfc69451df6c163abdf01e209704fc7fa8a9576f2aac49ae32324aa536f34849e2a470610ae3591421f05f0eed9181c577d56b37272f0ac3185d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3606a737a9ffdc9fb8e8f7f9e9b7b66b81144c330fdd439334ee9cf658cca19b4f4ad831c0955fa3653dadd870fe2756cf8d2fd7db30ae4226d0e4f1ebf69b97cb724af1d83fa0d085d4ad491189e7523a12a6007b77cbef9f77a58bd389c87f9cfaaca7730fa18c167d2ce55ea2123d0ad1f1bd9d58dd8c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2faf86fdcb031caf2d872d65f758173af45a8b738f0f8e9cecac6da46bf46f08c091ae528459648742c56dabeeb279aa7b1fe2290249105c6ff6f0c6c965c509f22498d12f40282cc401c068611557a9b8b4a6d41b144de15f98e1ae8c8d982a44b1f7e039c0f07b3ad02bdd41e995da9d61b212e508480;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46a28393b087bb14a2b86b9cff96f46269742246b63a4e477a2993ec0cb9349f5732172b9f4582a625bcb1dc286fb787867cd18e21f65f6b6c9104f2d9d2d6fa342aae39919d900c77ba8d558e39d3b6d608f7aec1fd8625791e18afde4a40603a2eed0db9ea50500f0ce3796205a2d467492e8ffc649eca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8ecaf51e10ae106bb11b4aa9a842f56c391bf2bf762ee6c38fb96c2655efbb3f6072ca382f5af51da1c7b160c7b957ecdb678f9f2e8fb69f67df518e6cbd36757a02e7451214312a5583d6558b281ec43aff7198152cfbf71a6b8c5654aabe81b6040e72127526ea4e652cf7dc4ffd0036ad2e01847a964;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d93edd64ba5bf92957a47f46282d3ced8ef78867c7ca041af0af40429ffefbef0dae86f86ef1fbf5655a6354aaf2f3387497a72cf5d766cc8bbf66f7d18125b1c1997206a35514c2b03b42097a6bb329850cd1b33f4f05db4e8aacbf96ced02e9818b5ce01f56199c8a417a381c3f8961517314019013ef8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13afbb1fc15e1a594f95abc2a252ae572bdf41f9c257de687e805c3ccaf1962e00018afc4fde230ac7cf4bfabd371261ad2c95b60728f107c2199dc6879fe08a05144385662720bc0bf76d9e237801f854b6cba7e018c45f74da8cb44cb7851a303aca4360bd09caec6d07afec114f38b94c28c896437cd5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae1ccd9962889dd892861205eca6e264f17bb81e45ba1730934575a8533229166ac2cc8706500db448e612fe35307c56f08ca555cf69d3b3fe6bd8c9746a88d1b4dbca132c0bb2646b37f2e0f19d88265ca09289521f8461fd7e497c4369428987706fa169d90c7d55175a55f40e79ee2a7a0b37bdbbcd10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae93f497bcd8b6552ad3544bc105f37107c54e316de4bf9ba67542f51bd1f9e3a8b047c83b26660f1843ee949d0555d4b32164e7ad3dd437da60a9f962ce6791974cb1b6c49ca766b1c92937eb79be407185e933c64a2390294a61e372b3b0933587b16dfa938a5c01c550a2949c12dfe8e972394cd2ddbc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3baa09ae0ce9a26f13b7c6fdb57495c7acca4309aee9cb5ffed90e39826eb068be8391872589d0801dbfe0636e120e28eea33ad5dfa01ef95da7e9d8d79d0df689a46d8aeb3a8cd06fe4f3c85fd8775df674eda02296b8f1189373022cfbc975f953b64b433ddf71a26782e91fcfc6a7be77a39910bfac4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1832dd777dd3180e28b34768c239873d26d3d5e9540de906bd6cc3b7e2a5a73253eaaae339d7fe5a58ff1ebb07c9439942c19efeb801f2aca2487c55d20887d0d648268b38916aaae4d09de11f5b41b501ce076c6b59e85d8711e70a2ad417114c5aa62ae03d5bc4aeccdb170e737552c51a09e37d8e3d3d3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ba988fd98f9a5611e489c7c5ab4bee1f03c64cbbb5b494d3849042ebface8f422306d45323e9c959206a78e0ebc17fea55e8482d805735e05b3a340ccc62b2787375e8382beff8b252665b242191f5d1e4dfbc15a87f4b1d19ad81f2508df2dcdd1e0a202b85d0964cf355451576e428042ba1a02c08e09;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1759aaa98aad397ce8b7515f891dbc471249c45c9a1ee1f9a6cf36e6652f8676ed83e47eab51b4b7f22646577112f0cda37d10072841a44868f60cf59adb4747af50f2e33f45cf6ffc912d6c688ff669b88bfc2be5394ac8236005a48d01ba3123103b389014da96dd9389d0244b853879f28b6ea9dc48592;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6922900aa111ed4addc0df68c3b13ca610f2cf667c1473b6805464437c90bd19e14f9d0e9e19208b7c77c70c1fceac40a8fa0ff6fed998a57dcc40ead654eb1019136eff010560495633fd8f17c8e67beeaa073e4e424f4880edfa62bad02d903c171bba51c562382f65cc1bf8744d0852435715fc39532;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h642d9610cf6f8d98733ec6ce59c6b2da8b68c158396fbe25ef04a039c6c636664de25c47707a527b2d4c3de557f914c7bb960ce3b864e8f1e6f4a71a2afbbde680aacc987d1da9d241b25e76d7265a8996ac7736e9c8f19302d940d1adf105a44b5fa815df62c9668c16feabf694c3f07b751bd8626ae335;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a70714966c537bef8931668f08c628ded321308785cfa1e5b76846e1e81bca7ba0d99c7582409f7b465d655f32c4ff5b114a09e2aefef6f95b935cfecc1b3f9594e6962d10d0e24041e6b8155259bfaf8a8928adfdb3cef9cff12497887d517ad3b79c1f2dd584318617fe23080cdd834784603c8fc254a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae7e1299efe7f0cc10b48164aeff6b08def72c5995f048e0da55e87d3911037f0c36a0d979ae641e1751cf68fea96d7e443e2c2da3379a99f18358182dccf35172e562e6dd0a33b519ad96d0464b1a44fbd9e8549ffb7680b6e9b83ac666f82cae62bc7bfe7d6bf23907652f2095fdb1657cbda2588e5045;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9decbeb76335673fae537e52e6f4a2cec4e9fe0f77fa2d9a1f950b147f36dd52f18e93d888b264c33000e317af9435a94fa92dc83f4cf27e4cf79d787b5ae0a316649bc7c340794ed53854185192dbab66d080aa35cb41fd8a131a4804b2ecec5d934630ee2eba8f958267e6c9f29c9d1f506e70084ab9c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1365c8bea04ab657ece50bf0678b31e737e50d82c0750d2ad8f5780d227d6d9b80e1043e933b0ce8db49273cab1baa354926af98eb97b6dd8f3744b6858a68aa75c2854b51721f4e6f48f6f87ce286cf7ff6b4e2b98129a337344317459b2115f7c7141b3d4763eef3b1890513603dc374dcb8e8725657cee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca8b22c7aaf7a49800c5743a4473b7ca769a1f125b44b83487dfb46e54a85c6930fac678c1b041a96b3efdd82ab7406d26b4817de75b6b57afacd07fb0c242cfba4a107925ef2dedefffb6304557bbcd6a3d4a7fff358f9ec1d74a12b8383bf222d38a7b0ebac52c75578e3136e902f8cbfc94ad6c62df0a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5fec0624a80b49eec88836678892a39830033a53ed2c93b54270d24aeba0c61531ca2b718f3bffa063e6f8d9df143fa8624fec5d74f439290c60e7e9b7b54515a7fda50ab217144306d34e8631ef2e7db2e3374a0640a1ac4c0ea882b2a537d65eae117e74cc0873ffd02e67b901e3f33200a64a91ba676;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12283a9ca009ed29c06f6802ebbabfee00e8473534cb72f9b405976e6167a1788ddb1a7e51b88745429ada1db2c0dc201f3777db1e1182c8afb0f0cd545fb3d0d1d199f1dc9e5eac677d454c20fedbb652b9fae7e4e2014be2f71f767595ec8c3534e39bf4d7ffc4d15fb280553c305aa74fe66ac04a54f9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7b1d1036ef5b58c4a467b28e41e5d27b68261b453daf24d1ee939a4c25e95789b3bf7cf921be20b1e3500cc9acd6b72e926cbe68b3e23cb9fad0a066b0f0523e789d2d73037072969204fa91b0960eadbaaa26382bf2b798a0e954858dbba0c370d76e59cf7906aa666859ca61b96ac02ae87dc27ca3dd5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bdd0580cde8260027c72b5882970d0c3fe881730c4ea3d61a5b95b08728acd3a1d2261a6b37f85ed82ed726df24554d4f37b4f3236ef2329eba84bfee74000a696a2b0a83bb1eb07fd036c1a12018aee71686dc49338345335aeb82b2d629fcddbc118d2ce3b04a2dabcf373007faf2879765a2cb52df858;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1774ba4bfd3ba437e216407404e716178274706b7ba77e4453e708c55e03e00549f132157cf443d4b87383b6d9e474f49699471b2749c725f52a81d0eddfe78f64d9c76f0a2c4d505246c5f86bb32d29cd12e8cb1789136159c530d663406f9a5551fa0bcab659b9c257dd8bb0e093bad889610cc664d2635;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e8ac67c26057c4674e1d2825bd3514966d7b098a3d2c56d515613a1b4f2406ba88dfe0cf314c6661d14598e575d7147d88eb77e24b10a424461377f2fdc04671e6bb86a32f320693ede34abe4362ccef9c425d83d6f478de98fccd266f0c4dfe02b74fa8d5d1edbe351f3f02b971130976e0af2bf88365b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0a170eeee73a844dba06238cc0abb7170fc12063e16e6c85c8a617ac3d25a35be7ed0d8be15047161b88b1131d1df8e123858ce69701143b6bc7f288aa70f8ef4cab451b5c9820c3bb5d501220d41256855edc9ab21ba7ad645123b56dcbb37b75182f59e0eb2dc8730e040cbe8d586701d458340752d5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5ee9485a9a67ff11d0d8992e3c9799894765bde72cc0657e0146ddcd766052a8b40734c5ed8879feff7067d069a0389a95709ea7047b4264d85fc617dd82676b9d4e6c15a462ba3137dc7b8493917b8dd8a952bf98c5fcf3f03f930b8b1608abe5162d102ce9638e3e8a43fe502472ccc82e7e260c33ba3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d40f0b6e59797d12740289a19eeb94979d2b584bcd4af0fd67042a08a4591334ba7acbd6cabc0ce69798fe0c457ffa5a560f8cf5ab999b9ad6c2c8574e2c7b1c7c4a86c8da011ca4109058d66c095d29ecbf1d885d0008baebe0e15811389495b7adfa14a82db6d72d27e3c37647ffb9ab5c8d733e95d1fc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf709594b88572d87d3392244585b938d273046097eb229314cae5b73f52b02d43e8229bd5e2dbf72b14c06e1a3c79577937753f08f6bd65a379059cd89c4b85ee8b19a241e8472a9199a63357a0b755026b80f434bfa5a6da8ab943bcec79e851ce474e113918fb338619f0f1c9a5462a71857e42586ab3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16eac01e6c99a4eee83e6901fcbb06e51abbcd22f039205df6a1c98204da60ba7a9d02cae2c108841afc2cde9c9c41f4e62d535823fd597d24898755215bbdf6ee4dbf55c3aad5119cb1ff99037fcd2f1d2166f7b85f7c0bbc616f74a02ac74ae82afd7b48b632f6ea2394a8fe4c621aa2799ebb2ddd2ad83;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbbd05807fce2546aaa3000519913860f1ad184e73f4bc6ec3746895f0c9afceca731f2605b46bb93f9dc76fef42b8a1645cbd0755c27d46440827620d1f0389df19f3cabf0c1be72809e3bd77733118e037b3fa7772bcf78a59463731e9100c1dccb05110d06d35090af157f49e0c2fd78dfa9b3af8047e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1796e50984b7fcf09169e87a5b8e730f724d592c12395c58becdfe610f953e4736a2be1ba97e6efae059a6ba479691333504c10a0213d02f783836d6b61cf42b5f065107da8fa2e12cc49d0508b825ac01b7e91610b4d1de4e6fffc98851517efd993c7150d1e97748076d06181a4d555d2f086ab7ae99e6f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1effb99dab80e6112f90bb2948c733cf74327e40eaf7389c089da986f5ff3dc47122fd6f5ddbc55246f75fd337b76cbdeda6df841151d59146f46e2d9966cc4030e7a1d713618c9fd34c08fdc3d2f7fce96458b362b613aa34e06732550375c1cb287315cb560c0cc077e5948f09880590670bdf68aba7063;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h240e85ab78a5ccdb6fd869ed867bb379d7df9a58c3022b67fd1efcb51b8db448fe6ffc775ef00ecbba785c2b80f963fa6a655527d76b53db924308e4b5d304fd0e51f688bcdba3bccee9c4f651c674b55c0ec34420210121369f594cb0161d231060f7de3d04179d030745b50e3d62fe3831030076deb9ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eca48e8de0627c4bdc167053a589effebb15cf402de3eba9fea740fbbd3fea8f69293b3d5fbf72d62f65dfa4de8986ffc02881064d39cdba9685036f6c4f8e6e5c684de1d844cad7b0a53433f1dbcab5df6263da8f1fd1501b91344e69a2ea1e14e95da0dade30eedbc1121d3ff8e02e55ac960a33c26868;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cd3415fa0acdb279ef70eaf73724016bf51604d88d67fbc7e98254810c48b5b290594331fde6d9be1d1dd7f9d98ab72db5b979d0d1f0049d355055931fffa8e9089f942198f7e0552c74ebd063512c3a3adb0837a3a542410ba0d69611f9dee7777fcf9d0ebb970bd9c981dcc466916f91207ef0ec0d751;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h164b2cd858b97d85cfb47af6927f71a70d42463fceeb30b027ea03aedb9772c7636d63c0b7244a0bef922a3d298688a89886030c182ed9a5bf9da2e2b93cb555a383a21197b8558f7f4efdc3632fb967f3fc16ad190ffd1641daa4472b9cc29c3aa87d071548fcba1c3204a26cfbb6310dcaa434d73ab182e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d46ea50c240ae6c4de2434f95078519044df62d5cc2cf83e43403a2bf9af8a9cca6d6ad3302f355052979daef70ab825c7779375fd87b93830c2a40fa09a0a87bb71032281a51fb3fdc0009145873bf0aa8618d28ba842d439d5cd9972f08f2dafe572741c13077e3102323ac73f4564cb63e65a0c25630;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec89908a1823d75179277265472b5ddf34976496b0d0452a586b4296dfd902c29d0fc76784e3cff93b968c01667cd3544218ab593d8f8ef854765f17e5141794144bed0ca8c1247dd1f654de57b9560646905c4fd00f15a720a4d803b6041088c9fc2452744ef10e6587d622f70e1d33b0881fd4e3c98200;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128bbe132c0d5e83b40c0e786c1940fd7db0ab3fb2351db1e185303159be7dda17af9c505bdda6275844dd5c967f421b7cc3afea13778c17873543b40223c0d33a6dc98303366080a21b0b5aef8f5ad8af302a829a0bd363e89c7853947e59c099304b17f528f56b7b1b5ee65e5d1487edf4694b0233c6bb3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h361f6c3b31c33669483bbc59e83d92893f4e6e88682315fde123bea609f656267f897eac6b94f70f4f7d61450976d7ff55588b206243156ede7b12b77e7b00047029630b902e517e36a835cb8384980f7f7500a8c3f2adab420a3ac8ad315a3c76493d1aa4eafa6c5e21614ab2608997944b9fc2558fbb21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h360492c201b6975d577373078a4cc6e6515eb41765ef0d10e38376e42f6819249adb5b03b1d9eab90f646efebebe4de853d5c9f3f3751be774604c82a5975509561dcf151626613be9261a565993cb4664b273dece1ae4ed1f79accc78e8d4de370c4954dbc38f210dfeca6b1111a59fc5d7da5ce4c9c2f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ad43e0284fde822c547025451b9d91ad1a6989213786b6e8bc1ece85cacdd89a1c40e85fbcee17001cd50858b54f1b10d446f9db91b309768f179b9032a19d70e27f7471a39932138b1cb1d911103f22e1ce638a3904514c7d66125b9988bc9d5ec21eadaf831f8dc01be37349471f937e7a15da78c6df2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf0da494ac0fb88265bd966335d66987b5dc57ba26ddf851b1594cb166019584d9e268f41bb6708aee9d7d30fed260728047c3a074ce4bb3e2bb6b4f0ffae4a6a75a571950916dce4163d7be1a7f4d52a92194404221e3ddd1bddf0d608a9fb8260bb85d63d02743cf5c1d0b01ab675e2da3eca8497d9220;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee96184a05bed286feb9f34657bc754c287b8496b3d6ddf660d57d1ed295fa81fbe3897b761a889523ca06f2f8ac1cbe7afdad3b4a3389cb69fb0474c7fe0b9de69b42ac20b8a7b71daa00f67501b22709aed7b300aea0de0e61b0803c39faceb27e572f93b2907df8f9867cc58c445a229b1d230afb9723;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he662a189577516e815b41f9e8087d75a54cea8c7f8da88aa93e93d2cf71720b5cef809d6d54d9991c31dec9dd13d8cc3b82b9fb8fcaf5283fdbc0e350b1143bc78ed64040f0d2ca1e575babfcbd6fcb5cecfd92e7d872442d86d0f628fa508153973e1185227f53885846bc9e375580e5921dd337d059ae9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c0708ced98322cf2ac2ddaa6bed3717a7989e39366042a5fc55e6816cff9eeb9cd87223c28a57a0345de8f627d6946e3c246cc58df3a4f75ce9ca018764048eac0e4e61f06c93f2080899eaf5bacd7f9004e4d1cec8698dc2826ce0044e8ae861793c1af7df9180bb2eb906ce0990e9a32e38248c5de5ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170b542fc7f10284b908e02d622339031f323503c17aacb900e8ebc3c42650c2bce3308333839e4a179dcde80fde9d38a45c10ed984ce96fdbe75f44dc83110d885e5de9d8fe3a3f659cc4bbdfe0e20ab7735173629c529ddf7ebc78cc9d9bc20715466bef4b35a7de23e80e3c0a517b13665d8d02e633cfa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae01a5a9b593a3b1551d43440cb110c9c38fe182bb63bbbf6a4f8ed80f788b7b685e3c351e2ab2cb6558603aaf0a50465051d8a4c554b3ba7df4fe75b6e950fbe6aec4798cc4c6008f8926087da96ac2699db4d9d5dd85778b43457d650e18a45c7d2ce045c70e50139e7611b34953488d1d2a1e5e23a877;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de1027a618bddfd90b056efe9c248f3c14dec6e18bf9e68efe8e54b409b630497d7b86e7827182367345f2375c6db7f0e5d65b318158746d267cbf682f9983e1abbfd8d5f133b89445b7efa0150d1372cb30553a91f21ae4a3a3b0481930ef2bd7d66bf1ed7ad3649d820ec265a0ca501ac1c325f248f44b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8971981925f6a73f7ddb50b554e2df05c4f460f542d61a95e6e2e6c13289e832e5b24df72a75924e1e7fd0eb813597881a9a3de6ecbc82c066a0c999a40f3087ec4259a6710055ff05e2a414bedb5cbc4c9ce3d22c36d7772f4f3262242ed358c9126c4f75916a2c105fd5ee312fe739321ce5776cffe289;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a6cf085993feaf30ae71767113baadd6d1568cc16f69e42900c561ca47b65058c401034af2be76916665a4cfbeb7639550b28a57e03319e9c576d838b3e21fd91dc5383713401d114624c9b0c577a1803c0a4506ea4643cb7777a2fab2ce2bcc1dff1bef80f50454ae5bbd4500e23c5d670ad3d39e89aacb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf298c85bca458de42f4db561320a5433e04f16aecf5c4560a643eb3dfc131c4f43783bf0872a412a6532a854753dbe1cc1e5fb34d529c5240b07f580ff67f683b141216aa7378e44b9966473cb377027fbf59e4977e8ce42c37857591b942a46c91759fa37a7a7b12f0f578512e6eb340221511ccf61c2fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19314601a444e6402b6a9ddf44d51da53a004df8fadb151f306a42b4a476aab017adf1e19b0819cc9962e491d41824dcc942992bc1bd4f666f1d0a3b09875090a7dea59db3b9b0c0868a82e3bcb9d762c58a9e999b67d0c61f75854c65160433dcff5b1d4ba3ecc7b5288918b1d903d2b7904fadcdab12544;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c3ba24149033a69ea515f2d57362ae5d2d4b4649806ea0d9b990202be1320ffeefb6e9909fd87011d438d836a4b858b8fc23554d3fa4be6e598461798bd0659091dccdc0e85a0d8f8fa977c75630cc0ffb454332800877d96d040a011a5b9ad3987f986a6d7463568db70c8fdbb098b73a21e12dfb79391;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcf5472a41da3462095ec71c8fd9314d2890d3fc87cc107d158f5369bdd2a757bb662ae05ea3afd2a4a17b44d764e6bc2df1b8b0ede40e0ce46335a2e908f191adcf1e5e000c0edb1b5f0d844a8acc2c293c99db8f8664933346445851945f4ee5c06bec2db8b1870b8ba8f71b74acf8b25e151e2d8e204b5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9258b4b6e4a6fbb97e8aa194061f76801227007343e37a2ec7ee7d7f58db1ce2637d1ee1ef0da3bfa671cb93ed3dedb87a8c708de51602ffe5e3f457310bfc0184c59bae981a621d0f0bf39957ee58eb68d3fc467fef35a5925a99760e6eb8da69c1dcd63015676a29420f25d619796992f570e8c530fd7d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1500b01ce3228454d257e95989c5c87cfbc8aa0f4024eaf18b78292946eed02efbc4106fd0270b13cdd41ce3e9a9194a8e3e7b42a1c4ba5ea1667a495e5e9e0e16785eed962f2b9c187d42b6d9ef2d0045a4b59f6e62f74169bb4510d39ef7f0e1ab6e5fc7287d541bbfbc9e67ec3f344f2a5d1dbeeec8682;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h872609c8146ceee22854925c05c26e6326d69c8fc777d12426e2126fe2d810abdf07ab12d5d0b4daf0c1781727ab54740244a08a0179cbc20f0849f8817fe77224f62ba1e1f9ccc5bf4372ad67a7d28af93eb374153b284f2814e0cfe77f8f3660f5c50d92883004ab30dd92a683ccbee82a8040decea666;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d0234847619da7bfc2324bcf0ba85830a477ee1e398261dd0692228d690f52e8f610038a733a0bd80369bad73e30094f464b5cf3b69afc51fef4c4ae9108b3ba4f16f8e1ee85465c4d89438a0b65cc96ac429e1ba21ce6fdfe0e04f516b22ea9589d3bef138278b8bc89d5447207a255803205e51b08b30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153506a43ea94418d438b2836583351cd8cb34602bef6fdb30ddb963c42b522154bb156ad0c34bcdd2bf791f731adae3c0afe2214b987dd61ccfbecdd38e521d5611d3d261a77d6b5dc0ea79755d790105b6fe490b52b653bbde7833bb72c9d873c95fb126a9279aa2f32b17eabdf85f5bfe57e02bf2ac60;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52e5a5cfdc2bf08a0208434b3f56f9166a466487dc88ac18d954c9f03ec4e7865a363bd054e99ff604d36db81d8774c9385954f14b996e12cbe67c4d2203e9e43ad4b557d6642ddd66daa620ff94097a857bc1b0e7e8016094c27892d0b5c200a8bcbc7167208e9dcd9e0cbd162e1b05d2889cdb26b956d9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18fb3b800ec0cbaaedc1f8d364063f9cf1d009bb4794e54dba0f7b75104d78ecc86f6423ac74acbe96c3f41ac30c34e934487816b80ca177da2e6d86b9e559b85cbb6f72a4a4fb1c8c1283f9b7d313c488247d225fa108240146ef47e55c93e695d60c7c164a25899322cee104c1bd6acde8cb0c0678e9271;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed7a8d505339cf534e94ed62cbe3d840ef50fb0b9fe5f79867095e66b98f4b3282668c1b7d9a1db35a1f67c0b17d07deced25f08e15c719e3182ae7ba37cfa5277896686d09e9f715ffb9ea67011eba93ed0b7b2a943dc88aaf28c389c2a8e5064f64ca274851da417c4e575bbc5fe78a3c4557dd1a3a14f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161a52ae141ac7d2c99c140b3e951f4fa4013e753de7d3f18646598c75bf3176b64d46d534275142012464ec586adcec933243888432a4ecfa03ed0824e56818443ececa8c5c03544adce1cfec777ff35cc21e20bd40d6ab67ce84145040b1b95fac4805a24bbff3a20e0bae04b7f0945ded090ef36e3f439;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2b598867522b9e9cf5823798cf78dea361d588b29f7a136a12cd42997ac683ff53cd559409568fbbd34e84d05c9b2f0e1e2981cb837087c8e2c63ff935b7fd4f2eb5583f785144826d3abf04850097d934aa0fd79a7a14b9664da28047a90fd4c8313e777dc7548506513d391347a344d7c4b39515a0ee3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1caf5752d38dfe7b51565df6f737d744a81a0fcfd9ebbaabd8c3bdffb4725d7913c3f8b3cf6978bcf80ac4048f9d06d29954314e6c52c8fa12d4e2bc5304a637acad6ae5f345746b771d40437452d8dca59efa0473d80959de3352530092b2e5bbcf193998081cf38a35796d3d6425aac6754b685f67e8c54;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfacd6257e536a650742c5c1c95aab7a22411b4732a1f27f91c052fe63a6f88056f6d4362aaa9c0fe9d63db56af3c4e1812439774d6718a96f4688c0e319dad8d74325798aacf70e79804e2a375f961a9ee02f4d3cea6f44e5a027c81fafde6353337c76a38b647c5e032223a039eb4484f040ee3efbbd36;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152c63b81ff4354b1cc22706d74880e0854c0bb3783a06347e957a38f1b6f67558c40355380b63e059e9d31707c6c9df53b4f73e12d5754a46dfdbce14ed8d8be96a8b7ccbf3a1c9c1233f7ca95edaa3e001d81aadd8b650fc44fba14a13946e47288ba838c1e3dce8ae5bcdc04d5cd658e2a836288b84bff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6dfeeaf50a2e7f2e1ebfc475c588b7f6ca6b5cce7fb547be22da199b0d34963fbfdb6b41873796e33769dab35657b2f56604a51543db94040fad8c7d606819319cda56e8889e2685ede42c787ae6b851cfe68b96dd67a9cf1afac9f6727dbffb54ec959281390593e10dc36579e779a3724106f0336be52;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac6be2de939de0bb29ba28cd08d76ab964c0296373bd8fac45f02e96f634b00f41b40e0b4803afc246cf1921d9b2c3d422065185fde0e18fda7210ffb5139144d7a6ef9f27ce20d2fbbf37cbe25146cb1d47d7423f6aed22717aa99c19ae650b104fc9365d6b82050e265844be18e37e30d563ce6cf332e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcb128bf4d6a56303f7e8b4e03ac47d10c493c926906be63128b502a18fbcc8a5ca3b200a6057cfe07e357a822dc1d5a67beda70fb722804c6d628120909c02701510efa939793811438a9d8ff9bda10d2fdd1cd55d9e38569bf2f235ddd735fc1368b989fb8e0b944f3fd337cddf5596df26be85c846440;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h628970d8ed4d201d586164fee228298312fddd4c885d74f924e449fd3fcb7b9be8287a9373810f8f3fdaf7b53b9956b576dc9868816502bd5c9b1e1e21f10dcc0ceb261c0f1d814a2f6e62ec6047fbafb0daa830e131d7fb5f40d42bea069fde2bb51a4b876e3760a3aace557c562aee1dbf658c643f3803;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ec7efa1e5d29ea5b324fa095f2104f01e80b91826c2ef8107e77401fee6561a6b8ac9d67a215a1450320cd640b04e2454ebec687acc5ae81bfa8dcd99ef54ca53bb09720aab77d0babb3529ec4fb258c3aa94666a7c3936008d08d8cce4cf31c9c35da080038545cf0b7e2ba559386c52f742273ee6a0e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4aa7f915b70fc491d4538c062b064bd003b7514bbfaad0a3d12d86eb4bd7ad9533911541a8a43437feded7eb666ae0b5f640587754cbcf6e7d9bbe66ffb0cd62bdf9698e2ccc3555319bdc15048b4392e10cc62a983f8e40273b6a447600f8635f4d012a0d6fe396dd984432933a3ee73c0e18bd94a1cd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f803bea0e700a2459d1aaf9d9892e302ea6f9833448859f475e10b08ca378ca0764bc8548755fa53ddb56f5c2948b48aa85455f64b2dfaf201c5387130eb53adb8115df269b64e282f660bdabd7358e8e8219b27d212659e4df98ff0cfbb19d41ef211110d3239e5f6252b984965dffb14351d7149f1f93;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e785e1842178a657980aac4e999c690460ecf819e93c2cb7ff1c15e9397385e27d20fe908276521ad2b9d8d44003825916145bf97597482acf3f81a563ab2254dbab0f0855070636fd8f5deec7a231c48cb01152102c01688cd00269498cbcdde10442a7d09067140de2587b3dfd10ec378ebaae8895ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bae1ef881c04bd2eede6a8fb6afe2985fad97ae6f9295000d58100ac228206045e720b8879af1f7ea9a7b3922adf45e57188457badf1600e47ca581fe7f1acfed9b78ee2dcb36a8463b0fa54186f8c9a21ebfd6dc0a88dffa609edea699dcfb472c966c51817b30a1bb1d4d4079f7fdcfd497560111f9644;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7aeca3651e217091f8907be590281cb2918133cec5dc85d536b6babcca9818de6d52afa80523c83c4c4bb75022a47722dd7a5c67709273da3c7e20487b7b899a50cc5c1d6b15d5fad197e76a89bcc9c20ef6bf5882f535b1823eea4fc4545ec2758120daaa8d21e368987fcb69a5f2f38c61c91cf84ee38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4cd4a9cf13923b147b86231deafc896db72b85c5005f77215307e8ea150e73b0f1bcb1aab38d2135b41680861407104c04753fb3f9dffdc43bae1e43c040b126e2294377796ae4bf4f005e81496a8b12df634d2a28d4ad7dffc24d266b23f2f6d54e17e6ccbd13574e9bdafeb257a0c090ac32abd8d256db;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14bd5eb51289c197fb32317363e5176e6b3b28320aeab2121df67d529a7925f219d794959c084dec9688af7659d15b36be78e14140479a0f2eb3e60fbd1bd225ce3a2ba5c23132b29a20a0209d04e9d04421d6c5e7a4e632eb31961260cae5a45056a2fce57eaaa7027525061f117a542ec5cfc50e9233c4a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c3b7bc7955b69d066bd3a424504c4a8357e30590d722e9ad0374137080372290239167452b8b65773e79e264ff6fab033ee3d5e2ade28aed71737791e7f48fd885a08d2000d442bd397cef1ddf275e3110def6d83d7b8fe8e938e63256b2ea9977792734e4e2366ffb246b1df4a81259dfd8230d858f5e2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d89a30f2904caecd83599578b62aa0fbd466e005be549441ff7d75a690aae6b1c253d69f6b9ed58dcd4bf76af738dd728a3686eaadd3327f65ddde974618f7172b7137e2f36eab7ed670ba3bc49b726e3fc53cbc9b5631bde6d3b98d64c3eee53e0b38a19643a22e0fa688c3be1816b339059f518eda306;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d30c8e09ed0dc1c4ebd03ee0b65e7a6dcdc65e1b461f9a1a7c7245372cd6984459d4102490f033bb2af4849b3627c28fab40f5316aa04e796d2afc672d2e84f761af3dff3a133d2bfca6e5009ff053bdf960cf019977b486237782de15e13eb1dabaedfabbac34307b0eb9422a756a2f94c2a67960d58dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16765a2fb2b23b16b7d106c5fa3f3bcfed7f580d796d71c953bed9a5613006ac5b410bae096e804d574952e4fbf501940d1d7496e34653f32934a9933ef95e72a8afa315602fa081274f436c3fd14fca1b8eec827f6e0f3d82e5ee6b3258e4a0008a4228f38040fbf18c9a082e2d60fd198a4d2e83920215e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1161649a885b21158bf0f613468a311b892b934df058d334352600d54eff3b7cabe3f504d2e30be5f7af36aa99a9c599bed0fd07e3d03124b786289a324f2465d1fa6bbeb5256e6f6d4e6ecd81d714e0536e8ff101d7bc911f97ca42c26811353576422db090b1525ad9272a175991e535115aab21a3a40e6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7057428f3a018bafafd66e09e9b3305138652519790f63766d0e3a916bbf112f945d07e942987181c62e22c98f9ccd46b4514aa47629ba5f9b554252c448d208418344fcbbf14d89a98899a25c31cdbb325bf7d0eb31293dd6361c6c53c0b6e93830a5a6f1e66e0fae8ff3454315bc0508b393e528adcb4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb44f5fce4de4485f718d72b93d2dd11522cd59921d2fb24a422136212fce3734f3b1cfd9207b83adbee394c9b8174c6afaf2f1c1e082aeaa096691e8b42e75a0b9c2bdc7ec39c3abf24b2933c81e74d31d57df6331050592ffd5f706240695918c777f7fca89537aa87892237510e7549ea6d90b869242c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf674fa99969077fded34d2c0772ba3713f19dac9a7b35327e7eac3605a0b53b64f3b41a638cc49178f31ece80437084de52c27e63e7ee38f76465becbb5f835185b827087aef9f9c838ce3f1816fb652c9924a0e6e39499fdd8e3fa9f416d8648664b2e0f436485c696e094fd8d7d19be04a72b96075f201;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12409d0e47b1bb71cd8c32259a23ade1c2b905dcc54843194ff064cc2c060605cd2b09696ca002067ee6c7367574ecf59471e51d3fb4c9f72062850170eb8c8d0c571725184a2dc6f440319537af1487f676bcf4e0bacda611782cedfd0525004dafd33899fe7df64e5416086164ea453383554f7a4cbf7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7f07d7b8bd946b82d292e5a525063469feb9c934472590a74242a3d84323f924b7739471f1b095a254246c60bb4b91d11156d701a7f059985ba08f2bf6ea1d5dd874590fd07f54c0ad69099701f7a11fd8292cb4c593f0855c580a4fec60a0e15c12a26414c0f5e5d44c080aa25967e8d5f702fb14c4098;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3550bcca969c5495f791d185dfc475f42a6d7ec07c0e10e79f0dc63a00102ad6f7da8962d0a95234fded62ad90e76dc100810d0fd6965527405a82c0a7248c01cf01fae14cfcc0cb1937023d592aae4ec59e36355d1b2ab38420914c99e8427f409f9cf375998b914a3933206a44ab9cf4bda29659cbb3dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a32176a7298c16b7d1d1a396e972460e4b3bb76703a0b010ba18cdcde6de421db5d1600e868547b96cd824650992919021fe8428b89e56a6c4691846ad0097bf133b2b59e854ce07f82b1301d00c87cf1fab0ecc7e111ffab28929f092a8a5d6d5308ac6256dff993e2ddb24ae13e1bb1255a327d8160f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b498a402c45b94564eb431321b09f402e5c81376806ce0d5c5d925f490c5ae4d3e09f0c27327a506bbb192046776d4a33270d55bc4272d286ec8f7dc2db9f41a815fe4d07e859527e80c9697bdb7fd08208f1ec51bde377d060a6fdaa2677290bce5675855cba198f409109f9d5b4516d061e0186175fcaf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e02b39eef3013050d4f9f6c6b02d2ed264c50de58d17c9dac5dec1f790852fc53f9b759540a35d8bdc5c666b879c1bf474c2b2ee246d75c6c5cd632e3789a999418010dae78cb468e74bf8a839c21f93759dfa94d95d9aa9b1265b0eec4b64a701e52461fb9ab7590f7571f25fa2ff64fe29877ddbb5cac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e03fb4af0dab1c62eda33e690059a166e29918f3fcd5a8804c0ec82dda8a76e87775ef16ca3213f74b02cf1786f53dcfeb8a2363b187043cc2d03f33927d72e122adcd20d720a93ccec103a1dd18ed23d87084215712990f5b2586092e153217ae548ff0d5b4d9926bee59a468e759491c9822a2fb8e9f6d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171d7d3c49a3f3e380fdd66b036be13fbab4866d32ebd62e0ffde78d7a482a2e27bfb61a1d35c0d7dbe7df4b5d895648f6e361f3261941e289c2686c2c0bb797e21a2edc15de2f05e72b49e26618c70104b9cd751da9cb256fba98abb3e2572f156f8a67a943f543c400a0a449863495bbf6725f05eda097c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5f897cd3303cc5706b7518b7dc36fcaf62a65048747a38f2bdfa1e39bf6cd71c09713c09cd6200eb3ba3dc2c2bed089cc3c16ebfcf638d2d85c411038a2b6fe9729ccc910ce03fc226cd8c69c43bd813e632a517304c890821a98e78e9d01c8884a527001befd33cb74b4c2dd9b6ca1812e227073407c27;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he001d7c3e8038bafecf0792d71e27f3133c42e4e9b7535ae17f09e2ca44cb2109a7abb601cb6d56ce0d898413a33da3d16f924c0a451be5cf898d934ef0bb25080f0b85a6f76cca91065d7976c864406157c5c7ee1c25dd217b162e19b5902b0edbdb461b1e63e329ce5be82d51111eb192bfdcc484acacd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1712f0951e1b1c4e1b0530d4888a6030a1ca99c4e3622d3df77c438c775623f67c21895452e0719d63f74e900b7f215fdef6cc1e290f2dff89f36267c07e153e9acfdb32b1d5d6445c90d80c9aaeeca76e3634e8abd677cf6aa9f0cf5ccef29962ca5ed97f7064f997f1e746efd85c8d24cab3c983762ed15;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddde51a9d98da2f049d21f2e96e781259039170e69f4e6fc492e67bcb54aa7f3700e8e5c2b94a2d6023aa2b5468c62d77d86bbe2d5151b6c81fd2618af3c5dfe4ac9080b9de870cd1c2dc2af5d001113fe8d91d3e52ea3d8c7a1d7b166a3fd6d6cb7d33204e6a5040935edc73e23146402e5b9292e12e095;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc44eecdb24e89860f3f9ed7b92a66781fec435ecba8bb31f60485dbd4b26f8c27e28612ea7bfc060b5ce499f6c5deed22e8d720c6f07a03695d62baa53fec4b42a0c33520a390839263d03392d810988307eadc17d14057a490e4c1387fb4fca1ff0fa24478561eab614103770819d7aae1dbc615767e562;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13529b358ef635caea3f9dd9a3381880854b8cb773f95033d3a0e4c54942a94c94261ee033f6b34aad80c3e235239e1aa1edd961d0b4ad0dd07ae2d3728ffdd48b4d8c7870f027f9627f2c829431e0db3d561c8af9bc07ad3cc8c2d5b4cef34a0be0c7ac9083ea622d3d4245b85b2ae47bebbd702eeb5b32f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6214e416dfc11210028a86218632d09b2ce1a13181d2244f31df30a0110ec913a32eccb6d01769b2fcf49bc773cb9c2031b384b338d6650e58edd1c3efa56983fdad14e88b4123b2bb1217af4a4c8c636a401509fca9a7ebf4fce7357f961de9b7c14517e4d77e68a8b6473f0f598104b0ba7e54da14f333;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52a2efa637642fb99db19590fa37a4a2db79ff0c5262642ca1711182567f4b84d65550c6cc33687f5c00bb9484d540842e3b49b13f999581d9b904a0de52e2136ac1ca0064936eed57452b9fe667e0b4626977447bcab74a009f7c38cc1b09b25f677349dbf23f9397b7d3c287bddd67146abbcf49b603f7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c749ec03a759ecc3e76a9a9c3842937e31787d31cce80cf2c98f4843da5cfa842ef732aaec5df8ec3601f22fdbda9e10a8e690823c8f03b3a0dff5612b25cb2c19fe76eb2ff8bd9a643f1ba7528616e1eab3ad91890ef000c274c8ed246e25245f0bfba2cb6f10cf4934c9dc83e09c9af2d02256d88ec82;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b2df57f8408495c19cca87459b88366335411775ee845e702850bb9dd583c35c8930df982a8b8b39c7ed1a991a08cbd07c997e9df82479bbb6d89853c80b031530222a025e28a72f017e540b59ecbc24a1f3edfe3dd9dbfd4797113ad3abb1558077d28852b6ef7edfc4000648376d3b34716554c752952;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he45ede93f8215028d7bdd068327cb82ca41fa91f749846c93b64c2418f2aba9088bcab2df1362c0e389cb31b5488d30f68844628d2ff8f429faa0d6c9a44360459d611075dd572c5d26b971fec65b0b7fc8d2c364cbd8441de6bfde479f11a13677f1d640f606616f3d1aef5188d63333afded6e68d650bb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdcbc6232323d90e9ae8737e097ee675010d6329a790d35e2bfbeda900cb28e923e66148413d8368ae62bcee3fec4f20026b4d1b402437b38cf6352d712d387a35e5f26fe41eb8606e68694fe71a82bbfd2723795aa1d155ecb4ecacd0c815dd13d25ed1a3400aa6b6afbfef5ef3942521edf5367ec35e378;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165cd9d95c83bcc9a07d39b74ba46b5c1d0597831b482d10fefecfb8266b14da2ce89f4c21a85ee643f3fdaeeb972e38d13ba4f4a2527b21cbc644dd8ce4abf0b33b9c8b1c79cb5cb9b305f3252168f06d78ecb3baf663a623223aeb32b7aacf8e9970d0fde0e6113bc127911d38120bc4256197be93bf628;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3bda7cd4f4a5e20d494f5e96440d735831cd25cc8b79b6e51994248abaca29749b7b5c3773cdb3435c4745b66d9ae51f56621b1b08d2199b4eb1bc18042c7765e9300e618694c864a9a08fd88fbf610edeeadc292350983197bd2d35f05961d470514e3399a3d31683e173d53bcf36bbd1c68b3c329de49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96f649417ae0bba7d539252ea865739a2750532e624e26fc67354a83bb5ca4a5b445d7778fcfb042121d424bebcf036e001adb32e5df463035c849207cefc492853fa98efa114e108e68431f6ffdc0ce3813a0cb27d01d638e04446458728bf5ef3338f686efcbb34eafdfd9cf9e747850f4e00f8e5de2cf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166476d96e9e8e33eafea5799e87fcb818c4ad9ee7c38765b069d70f18e8a6e334f5cc219d55b5d811d71cb7ad47193f7ddd90daf23e1b8c28f2a18ea05f20254a92ebf6a2699d65a07eb128b91cb6048855fd344c25802872066681dad260f5befc5a19eb51e91611a7935e2da5b0ed6618936dfb24ced07;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14eed062bf0bfe00e641caba8a05fee378be377b3272bae24ebe58e6dc8f4ada63b14d7b310f956a68ce6b2b0f44bdfbfed6567fa1eff187e57972899a9f609ef38c3dca9ebaebfad80577ab218b9f04dc37d7da216c2e0fc2b2f4e13e7a6caee834cb56269c209fae6b1370931306774c9b1941e8dd41675;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68fb42072773a90b1469dc3ee4e67d91066c32ea3c8030e9a7c5f9ff93ce5bb4950d6fc0a4cbfc4586f8690e7f07861192342d512e3568ffaf5b021ecaef0c053e5a7d527969d3f8840b53d961a2b674e9d1eb519d5b05bd5370a547834aea9f7f07697e2cb99dd5e2cb2674822a8b6aeb8862bea23ac1ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a963b99cdb814af03c0fbbb40bb8a49a72d1eae09905c62675ba3881a6c7522379f4ec30eaddc04d4e025d78432c103697724285d4a175a43ae60a98d20f8a1bb97c154de3d169eb74f8cdc50ee3998825bbecf709050fbdb7210d2cabdca0a8be200bb6a155486761b93fa0efa48f4380321886fcce4fb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa03c4f083474d2e0e8ddf058d17e222602bdf29ab3ddc41c3058124148def21a785995fddf4c1abde5ed9259cbaf4fad15b066b68aeec63d32530cd5343bd095b70b44611dbda119181aafd222c69afbd795a4074a03aeec077ae44ca8078145fcd0c459e4117dcecf325c90cef9cbde1f91c6235730ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h838a4b2ea52062df2bee6f756055840a336aabc2383604267cfa7da1edc30d9a283d1677919b456ff1475510be45e621a8ee4bfb8bff76de9cda278e252db185640476d9f0fa10756656d8a9f031a56e065ecd491194b9e794c72c2046f0bab11a90fbab88ac0ed4953a7876559fd159d461a4c4304b0a1c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e8ba38aea558f081452c5770d4518f855757f75f9cb902a9dc56657a195f694e5e91c282dc9322a20b5f5882da0f34c0860bed42f1cd526e977f47a88d88df16158a4b9ac7218d7a4fadca7344b06f45be094831d9878042a0a6c9bc13e9d418d0d270e8b9ffe2dd9b252376dd63e150b684b889792df98;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b3448761cb1009e7b8cd4b2c4a8bd951f074eae40559a35bf94ecdf4b0cdd0c6324bd4afd6159ada567d5643958bc0498c80e1ac8cf3ee1ba5bc8389286190d8d8b126e9d7f4c300b150fd12cd4bbb24c7eacfab1c685a2f35dda4486c4c8e4455fdeb9e5cdaa8473c60c0a54a2afa681e3c935ec4e1354;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e12fea513722bdc2a9aac23357ff7dd3fdbec54568ff0ab79de605edd392ce9973902c89558cfa2c5c69b75870a8219bfb01a87571c4fa5ca19b60b49c85af6564da584ade3b15e5f72066d6fad04aa45bb5ff41fe9669f56b29f954a1be0da7ae5879d2993f4e35ceddea8e6632eb23dcce5a6838c5225;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187d382863de661417269633632f0999cbb445f2c507825b73c9e3ac1f3ff494166433e81456bf4b38cba5fecd3ae075179be0485117e01a063bc3420958263d84366e48c8678e2542a0a80c8d0f62b579b3955069ff17e38a5ffb6af55504fb1d0844eb37eea4f6e5a5b615a79c272050870f9b7e7e45ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d312cdaab0715e565c988a4b48810a28e4e46a20e4f6c2297aa4bb387f905c2966cf7b6d9450e5aa2035f133540bfd110de59a861b4c90345c766aee6a3654a061518c5ceab38ced4f65d3ee7f102676dd8a047f6c6cb88bc22a3ffcfd01bcc4750f024fc86127f8dc5b92482e4fb29a5b58c58c642db9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec654a3b4b2afc73bd5e403d8136801af835b415fd9b0a21e7d469df0f0b563a2ee2315daa814953a7f74d91cf77f30d6246de7081ac05d202fac111e99b6bc36486b8030fb934ae18b46f42d4af8c917959c5d288733d954d25ef70d180b66d1b809b925bc82ebaa92c9c9be0c1b7feee6964c106d840ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1084669f0baf10ffe73c97a25ffa2f2d6e6efa85f173c4ba71585ae08c222c59e4206d6dd293dbad60438bb15b89a42e895d55c838f7644ab2f33c4cdca9977ae49318864d1726be70e65d0746dd7a748a588e539db0d011f6d41d0ab902e944b4cdf3d7fadc28169d0d9af880d0f192dda4bfcf89ae263ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9466b4d1a76f58d6fc0529be9abf6b21a29019ec071e7c7530a9508f86f59f3fc1b8b42002c2c4531dc1c1b7aa916b2b49837fdb6865c2fc89912594d90a8367052a7b31037404dc97f5e4963b93ed13942c46fe5f8dc65a7d9a07049e60c07b87d5a2408f79a560e62687e86cf9bb35ee85ca130a529eaa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8186cbeb794c2ec0b80134132759ac6f3bc1d5584034f551bafb2474416470114828c804f6c4613b356f4fa50b6b59181fd7efc7f7376d9fb8e831a4ee96f837f84905a6292a79d616f39d090683c8ce47cddad2c0d483d4ac70024f1f535384ad4b1a9ad4728485104eb0a16d2716834d7d3a180d5e1c14;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e3fc7b4a22becb61c2b585ae8417663fa6675a759e096b82dcc56876a0332b8ba137a04114fb9762f92e581b31778e1c7c0a8f90b63ddd956f2f19260759081183184022652fd0520f9237ceb13c51bfe5a0660baeec1164ddcdf4e634d99b0803e74627eccc7c99c4eacddb4635152ac24239db99aa8e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1847780e5ead747710a05074c96883c4166b9fe70d1bc76aa006c69958d6f76c029c0c344281b09939e525e69c0b4343e6e0ae198a36fed6154ce142d8cbef0a2206d97f15045e622a968c77974c69e6f847e4ec0163f7a9d246025ea941e309723a7d91fdf5ff9bab3d22214e2e9e9263834a28fc434fa21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1ad3f7c9b1356212f4f4c76dadbad1d8a06cb548ff15e2bb90bfd7c37ea7cc53eca5bb44af23ba0ddd3bb398aa5b43782a8f18b49efe69179b9c1a524a8f9998cc85d1322cf8b2663cdcf20688b78cb8042bfba8d9e197b6e16b44e30c6a2aff1bce0ff26f8d30923f8cd134f34512023ee8d174d526376;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5a3c30ba12cc7f65de98c6a4f576cfb31c2031b7bfbca24d81281c83c4e5b87e5d095e9b3bc5da2a7ec446b4fdc21710d3fa72ceb927625e75cba0d1047bb7cc99a886f82157b11453c4ed7cd8648bc60049db9614b7a5e038248e6b527d51fca89a06856894857e3be6c7387146330c41d08459b1a387;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h559c76387aa3e2eeb30ca10a5d498feb870b80be2de84591eb3b31a9c5db404ee6909226beee6250a4a6a21d0f096aef4d243706d52bdd3e6703878044591073018d65e3a3929884f31113522fe5b76ce8a943bf3868c230ab4f233ba519dd7dae4d26113545bac680674457170ec659b0d9725395c79611;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b37a51a86ebe2e0fdfad1b1f54774480db63f827ac0cf3b4b469ab9dcb6ebdf738837082fdfbf5ff3c5a5355e9cf1f74ee0ff2e523c90f68b6c9a4ffaf112f4c90bc0a89f443facbedaf3f46ccf06910bdc864162206d3e22ceb45b60f702fd465132efc7c410918e4fc7176757ff13a3300856781b426c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f250f72f7502ce3d479b1365968a98935c49b9c4518a7df516801f3b012f1ddd4679646006bda9268c4e9e31c079a5179bd9c05707856c1fafe4960039d362ddf8edda503ad62103b06fc41e3678e71b91eb8b61bf0e2e8a4ad2239aa074ac1440cfdfd183a39c242340601cfd1bff10c613c8baac16d2d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hccda43e8ab87db081761ae564fd4ba13b7b8c7afa27aa301360b567f5bb9e939082539e9ee5663a703c758a5ac046fc6072dad47ff96ae73f83c8640de328a90ce3325a0875831a33d35a7daa73ea5b37296f6af3e019b35b396228a15248813ccf8df6095b12d60d35ec86bcf274c65a9bfdafa995e71b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135fadf6f09e9b4b758cfdd0bbf2ccb1e515959aff409a8845f9c3e81df1eb3457812ca6e2bd2efcf2d9b3379e2b4f21dccde5fdf4f7b2c8dc3f69a014b3af2b4cd6abfa05a0ca8dc1ccdf350e3ead1b0239c5165a281a31b43892561f6f7c6ad52287a56ed79aa08ad02cf836a521c7c2170418019a6742d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186c177b354c556d3497860bc419987d23ca2c6bbcebccae6c22d636d00ca6235bbff5d5177d6105c6e827de309cd67094f3fe84f7541c149551ad69f35b2745a286230f7ca6addd5daed7c1bbf99f7cbc953560ecc5b03fa371cf7113ba54f5e09ad264377f0817ccdcc41335f6e190d8e0fe994272147f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1869f015928dd5037cc2fc70140b3862dd2b178348f5e2ce6d345b37a0c5717471710d0e3b1a78c32e1f52e8fb677dd0442b64cf2f144ce5240e2e2457276ee270cba57b017b5e776f1b8331804a327ab8a858b133767efaeaeabd7ebf433117f1a53ef82b8d053e781a31a8e375df7be40051381b0b95beb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e80d358104ff8c11548707b53172c5ca5b6f5de6ff9d14802e972a0317226e6af4bab4b5bdb025956c98974b2c929645feef71556774aedb7d125ebb220c0c4db8099a5b08f8d9a672bcebba320662fa25dc071fa8b7ef17fb61b1c50723606d7a578ec44881e5b267f3dcc57c9ac16972d7cc4e633219b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h289a46dee209293aba1c68ec90a779f038f52c7de2b40cab8e1ce71dd1b2636934981d4cb5de987ba875cb40faa967eb23ceb5b8756ecfd7aca38297eb9a9636e09eaa8cdb089541d199f8575e4a29068589e8b1d1b479f88fa3ba6c06cfffb5217dc775ce8f76fa53246fb59834d2633c9fb5fd434d0995;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf5fe539565768b2c83051e6290a04327104cfe9f864f9e2ae3f01249bde19bf8e3ff12f98f7f6100d30968d31d3e46a70961996a54202aa4f32baea3a2781111e5ee67b12a9d200d8435b05723342f4d5aef2109b6ab9cde55bffe937d190b1808c19f633cb84dea8ee0d02e141d3dcc3b2274d903aa88e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb43a831063252abde0437cbc37ce8e4745b1f2382079232df94b905a884295b8b627503c484b72ac40f833a78e7f617039edb49eec64d3f61caee53ce8833552625058c59955f9b558a5ea8bc40cad4a51413850276ea770090b0b3db4db4d53d6864132e8c309882bdfa4a086e1934e6942d286c341fc30;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd3292b1b2986cfe32a348aa7c0101340f82786c48023622308dd610edb7ad88f3a0b2af4a3b38164e23718d0c01e3bdc5a117b6953b4b290a276293c3a7960fe06700f81289dfd8898fc5a160141856b8dfcbbc460bc9da6e4083c13eec7ed310d6e24d5fb81fb36ec8af3ffa09bcf340fb12013076355;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e087efc36287f564d7f0eb04b888131477951a615073f080539c6ca58d22206210a83db2bf81d3ac0496fb7776e7c6d73f274284bd11050cb0cdf7a80dc1b6f6034f9093c55c31fe0e12f62f1043a6bb10fe9802f2f7cdc6855364be47e56442f192b67d5465e288f276007576b84119df9956675f7aaab;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163f3693d8718c49c6225cd2ecb51ffc71490ece8960eba95c10cd4ef315426022ca1e0a0af476b47c996345a05678394326620441c4cc33aad758cdf48c05af9aaeb3764ccf31983f782003c58a216c4b5d95fd48c82981ce7bdef0f04ada9deaed2e93469a91a64f775420cb3e52c634cfb1959da6caced;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf48b193665ec6d2c42163d11859d24e8aecb982a8193ed1fc4db55a029822eca209ed201fe71f387099410670e10733034c9a67606758961cca80d272fcc641e401958ee7e16d5de37dad4d6da89036e3e71d5a26664cd1920113d41da6137d3939311e0250c5e4ce72ed61204db466e451934f70128d727;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33257eff20041bb81eaf4c9e99c3b1e7fa46482d8e6539e92ac68364e62e7822a9f9919eb2acda36ff3945405a7bd7ed62ed213b9f7071a5a323aa200f38bba2041f2cb12681f9bfa4e67452416289c2470d153c8706e0cf35db910576ce697ad2a576fa0adb406451067a1ca168a267802d3d483925bec4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce8e266e68df3036c90d1fd780718f341f9c4ad509e49c2bec38bd6b8d4f1d7c0d92443d730f43337be8f288c27d4c40980d0232824c781dd134c675320d321a426834324b7022314c3721b27bfb466dcde1c104e21945ddb60f51aef7359843e39af463a185901bc2d6596e9ec414911a71547d3cd549bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7266e8ee082ff44aae59c6f76c2fd88a270fa05877a5f76d4822b1626bee95e86cb0ff921b77456ffd41673d14c945557ad92c11292230d7150b5cc14aa1094c35234f7ff296028da075290a357e180d37d4ff464ec7aa6d9541a9a3ce7bd82075a76e298f6bc5010f4942f02551bb2fc5cd0a76e9e5673;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1528d0a2bb7fe74525ca8f864ca9eabdb69e6e43ea5b16fd99a7a7fd727691408ecb45faa92cd98fd9f6cd0c6495d5389655a80bec25bcc980e95cc21bad2e6fa06c774377ee7a3448a973c53fd031c3f44c434bbc6b5d2ae1b8b5b02d64e446ec759ee81daee78d22ec4dc1fe996014a7d51b2cbc0e8f5bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h76f2d678d1c9470455545297d88b03aecb75649bb7196b4c4835d6733ac9ad478ce8d14a9679b6f90754e2bdfa13dcadb0396ab87db6c802c08881825839029b856f3bd27f4014bd9172f8e1f2f9ff7f6240e709785e87b7ef437561fb57cee72808cd76491788cff2c8fe440b8fca8b4adb7581f0549664;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9d0d623fb7c078551e3f7cc89f23dec43aac19d6d2fddbfe8407ff0f08291304f2452ca30ee534243e52b76c08a71c58ed6cb7f6f29aa92af4e7b2718e9c6fb4fb684c8295c5322087e9e6c8ef444478c7034bb6ab4b90d5b206e892ed75c2c8cd6f034da59fd204512869a6677b87e779d7e9fbd566a72;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a671b7a7cafaf184cc9715f98066f278e405c302203413338fc4c54b92e265fa82f6f654aa1b2bbda8797f5feb0f21abd1d827b8f0a982b8e86d10e7a5c94646fe9f9a288215ebb51a30f9a2b4ee59b06a7a5b2b1966badc61eeb720966ad61dff6c5051f430e5575c9217dd91c10587dc9050985c0678b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he71d4e4fce6d7504845d3c69a220376801cf1498d635fd5b7c4fa35ff7b019dcb26c18689dd6dae3ec566e9532a39829e50a44fbe741c5874be59eec22498a93354adec1b23c69786a211f797f4337f80db1743604cf3fa3951b9197962dba271e8e1fe94f91b5d5fb87623ba74d55abf319ac03676fbcd8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9f3d1d7fdcf858e8051b71e5fb1be022781773f97c1502a09254bbe0f91793f224fb7433af0d518466a735517cb6e240e0207282b3587e1f6cee43ddc45c46dd723cfc8ddc3fc7475ad48b3a8272603c6c09ec3e843565c256aed68932479c40fcd9591a3018746b18da784ef2a79875219963c48a2854f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddcf16376df302c62d34f6bc647f7395f7a6e5aecf3e4442b358f869bd93db0214df977dd7a552ad928ad6a70737575b621017bd0354aa82b83f6d3d5bc0124cd32e51a1338e98939296f3549c96b0564f29f17a319979ebca4827a1d8f1a291427fd2809f2649605e7546f31d3195befccd7bb1042a0536;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd84efde6ac6151072e586dbcfcce04d62e97c472a818e4cbff7fc5bb6d8faf67bd2f9c19dd6c7c7f3beec9ece30be1a4e8c60d87fc030ab14cec0c9b8b91fa55bf8617b4d21af02893cadbb9d2fdb5eb4ca92823400de512135feb09b8e519e926da191a57151edef183cd6f693fc6ca140d12307a093c4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2014f4d04c183fc2868a9e06f05817935b2ef6e64969e2f73a5f4fd91b3ae333677998e534fdae02ff581318ece6e02c902422ce255cbc2a0a70cda70789e4d2fa1426fc9f2e5bafc3cd01f10aaea00f57c3c0cb77d6201d25a56b6c6f16a4d90f80e09b9ab2123e7bd456215e81d6c8cd0429a5969c9347;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h299c9d703d2bdee67c2f7fc6076d1a081d6fc466aeb3bdb76cfa7557d4aff8d481a6419b1857ad60d372e9f4a2e8e73fd8a1002057282229651e4463a52b102d8fcc83ca2f726b1546d6fc0c41e1aa0e0e8cef8fa61b7a7e76c55ce6cd8e3b3674715adfc1c0a3006bd8725f117803abc7c91bbcdb47aa7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c54f36fd7e720cd1b1705d981ee3c9ad3a8080b1a5c2b8c8bae9bfa8fa350a9667b27d436dafafe31982389e10cba3dcba750b7fc6853890cf04ae547df3cae3bc1cb0cb72a3b73ef9382a1fd42366c36f93b6912de67d6e5bff10556d67755e02c93147a8299107f6efa840c6c108ad0c37b0a6965a1725;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5668310bfad6b687d84ea3aefe5eda85522d9f3aee4a26e78b024881a28d664a137d8fcae64ae386347cf8f92eacb842a40d0aa79e8737159f84ed8113c6f5ee7268220f4b1057577519b20a9cc64830d71b101eab94ac9bb5613cd341283a78f6c26ae59e755607dfceed047270a26269ec99b11ddfe4e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10831c67afa49927fa539b65e253b04fb311998a4117524ff5b815fd64ba0900c721ee9deb9a22190ba6136eb3c7e4237e4afa9b25176f45a9ca1ac0ac4331353ce26cdc90a4abfdba5bd46b817f2f65ef01b7afecf142363aa974bf68e3fe4a5a2cc427f2d7ae70be82f37197c40954c73b0876d0af3ba0d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8652a1eb336c6b07fdf011ad488d41e2667443c911be44f8777a04a77c32689df18451033c15cd62bb2b0f13e3ec5b96f7041e02919abdfa00ffb5794a7f0e2281f1fafa5a0fb8c438e2510a68c024e3903ce27f3f2c2e225f35a446fb454bad590bf1167bd65d895df9e151d6e8c9e1b21981568e35bfaf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f51fb7cbac8115c9eba8309232ab1a684334652e578f6c737e2e51858a3d57fa46c95b42af177fdeacedf273c5d88d3a9410fa5d45a67b35e4a4ffed62c846a20c7a49acfe94171e0f64926cbd7b91c24937c9577f049a631c0c4ca306956c5d48f1c45b8772245adda1098267ffc9dc152daff2ad4a07d0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109472f0bd24d684127155c4fa6ab40f16ff3117c9f97036bd2169be45c6c10e964d92b1efb9eb0766d9f4f02ca9eddad9ffeeba815ce75ce762706aa1d8328de492e1e5a7162a74e75f27170e160850d0cbe2a39ce6b29f62951987e0d821ac9ae6c3e5ca0290779b5c86d822ff07910c4e1f5551f8f6c62;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec418e7ef2a2900aa6ba2afe0e6802017ebc23777df30cdb269b95f616d2926218d4278f7ce2096e16272b5c5fc5f8e76c3eb3a9b90b59a7e829a9bc4ee22b995f7650ddfdae9aa36260e4083db9c95bdcac3006d0dd964745534af4b574b409780864edd7f950475266522123bc3cb33fb24a663f22d8b6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116fae1911dfa7c6268ebd8d4924c273784babfedaaad20e9b605072e05bb2b81fe58e8e0ea61de6ed7f6ec47d0b367ed50f001f260c6405ed46f33ab8dde53ee0d47852f7280259119f9226c483525b5fbdb44ede5730bddbf311a136c4c0e40ae4cbca43d48cbadc8ac459c66258454173a51c2f8cb119f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17bbfa125197700920da208e061e80cffd2abcbe8d625b55c34c559a87d8a87cdc35ad59c8e66b4074823103cc5d4f032d6ce7411eed48e7b14d5709add6a07db182c1d9e2176a20c5ff156923f33153159cbf65a33fa8c77a5badff1895a66cf7b9a8496356cef50fc3101e6ff34063f2ee852a55e60033;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17948ab602ed0d9fdaa88957a9ea65a042c0247981a75406a4e60c9200b9b98a58cd0057bbccfaa01301c5653f101dd4c018b28bfb6cf0744ff872a7cd27202907fa97fa1f242f719170ab1ed8c6ab6903ce7e65c30eae4e8b320982f1905384e4321866a236551adfa6edea3988d96b5ec27e85dee20b017;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36b9416dfa9fb18c4cd889c64fe2af3b1ca31ff2a380b9245bc4f88755e1a3b42a8a009883fd6b5eeb69ab0d86aca5a59816ffe3b91ceb823b653d42442e69da9d35e6718d574a7b73b55a60db47ea8a66dc20522a882ba905a4531bbf53c5aa83e2190331cd62ec82764b9a0281760b7f7374a9b9d6da9a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36a21b5631d2e3e0b5160e9b242a839e7bb07c622b3cb1034dd03701231ec5793655c8c10626cd402c180e05d1d313ea6256f938f78ed11a55c25a41be40fd49c8596eb734a6b7ee15222045f7d83c95ca1129e48309166859e1ebcc4995df4132e0383656714eb9144d06e16cf45bbb6fadc6a646629d06;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e10adbb71f5d0593a90c693930e427d1455ea896f88426944aad8224ad640f8b8cab9982f62d67b76471a0b5b48045520a5d5399ace44006b969a6b0f1d231c389639da2da808627bf0490384b89d9d7c2ff3d1e1af4dde14332b0ed2ebea04eaaf9e4a5db3ef4df89a716bb23c2743b8abca4702df56fe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h559cc4e4bbde87d5a9d8c69f4a9ade3e81f8416d110859901cf75a31b8332cd510d0e88b0c24c8688f458d3ffcc2b20d4082b8decfdc43a915fba2672f96920246089d2e536fa7f1137be761dca8469f67aeede694b15711181616128a8b71a57a66055ff0e77276e84b48cfdea5e65a0d0fc2d7a8b274ed;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146a2f7569a53614ff7716a5f36d4c85f47309a9e3dbdc3cce0dc37f377aa1e87baea8255fa0ab0b0273c7af3522e179932f272ead722c2283b2845ae2f3b5f33a5944cfd17d9af9bf742e00de642896175a9f1022883f5d569a5fabb392925f997e4221a59fee4620ffd1614da3604bfb314feff325ecb41;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe810c4a1d7d341d208219d9960060f34bf7cad17b7285509fcb03558332bd557c1f9055b70d8e29e4639e59a57ba0df772165a582327635e1513765c1eade405889b384e0f9087af9c0f8e084af5af538502ac74c09dee2d038b8e0d619a0cb550179ac3e70dcde84901e6075b2b4be839a4d7977650b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de1dfff63fc406d039d7eb98cc12da861f3b5818ac34d64784849025d3973d482eadaa8be26e0405d7ecefbc81a8fbc9d1359eba9576b148d174c6747b6a2cd560585a4a499568b69ae2653beb0cbd800b3a19c287aff7e6ffa339a4b9553503d15c9dffd1bad8c3b8fd6150d07e18d2218cd8d002903c38;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec17f1dfcf2ed66b975c70b562b212ecd6438e04640e7cf11574628c5cd941b940461717928a2c588ccb277772872343b2d3bf9118849b63c88e9c846cca65df9d4fe523b1fd2a36c09a3f0662cc663e73a3a7f264fbb8ba23a23d6b6365dfbc45ee01ce4432b735e111456623131589c22bb2e58281d2c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h239bc25cef0ad6899aa661e138aa19c5622ec9a0b2f9acf9694e4af328162c76e258e66e2bf9b75ce0dad753fae40bbe12477c85b62da20fce320723d0494eb8ba43358c1144263df153cbc1ea73173c25bfa1119c3ceda47981c2d3499af581bcdac70be62b896befacfb292b0da5fe9a91edcdd180a39;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c16672843fdc00ebc2e8c36095ff0d89b57275546082782c5abac3ee6e6c95c8e6e3c2000386a681a60dd0589ad4d100212a923f86e4a2f2302628d328064e9b2c989ebbe027637b1ec803e4463749c91b713a7569c1d9be5cc0873b0c97920906dc3d9e4972d215f6df16eb73bcb0bba48d35864ea0559;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcf4957ddf8a1c444925e9b546e79a9a6face9b4b264a159ced515a49fb368f8c038ef98c57e187aa716d183491031b555b018b26d4735469f3e1b5a71da507df22a50dfa118619d52648ed616fe9af092ba20b06f81315cf38743f06191e240e90a46c1bd2ed9e195e1da76535cd2ddd6378c74d5b092aa8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0ea114106a4fa198fa4239b7df88e45bed87b01d1b4184929e968e929a7609c5c3edf56d37477960e64fc388cb26487f88fd014ff9d86a61c863345b20f3b701dca3832273b6ad763836b48471df2ec11ee86fab7ac15d18c444643a441286c0e1c9649388fa9dcc37ee21caf6940a027edbcc90c961c21;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1698e8808eef76a1c6687611fa6810bc9b2bc39ebc30a4c6fda8ac925189a342d26cdc18f18a8a3e8c40e68718f1fd199fe11c75c15fc9a5e16b880ed2f0936026fbc75bba2d3fb3b124999bd60016e74135bafc2d40603efb1447f33e924af772af9a1bf76cf2fbdffc19cb097ada0805d15630500ed293f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fb5086bac22bc05ae66e4514ec51aa4bf6f1c8db68d740d6f08dc866102300b36e26f0af20dca5b7868b78d6c6bb2d81da643205d5c9149160f5011d041f067fd517fe0b16fbc7f163124f0fa5c8084d45026b571aecceef962aa6cab6bc283ec74977e03a4378e8449b42b27b059cca4795a57778c58dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h446fba816a5b2c626096cd653d57fc863e4ba8667acfcf85c0deae5733f79656c3ba96f7b410cae6d67aba266c3c9a19de4da36c44e71c8ec09245d0e500150b6b29af15a6f367a8638a8112ff9c66b1a06a99bcd89e6c8404a4026a43f289604159c67ca1e0a7bf2f0a5482d2de56983ae565ea86241c56;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc54ec2ab6502eca1ee2bcff89fb8847647800d9577800dafebab283bd954d38b584fa1664b7214cc5df749f49c5a9d15286eefea824ef9f0daebd7f5d9bb301ba84382cc242fadf0f4577232b5b78fe602a0ca0bc9c6145c7546f244061a4d966cb386eb4a0afc08c3155a0f1081c56989e3c1226a7059;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9396a0834662f3f8ba8ea5916c017e4cd206a41d4a81735961582a69c6a3b90ef7cde95259f8d31b85f38e2b4d6b7008ba6eedde9020770ca4244912cfffc704a7d6bbbf1e322da86f20821bf4c8918cf2f167ff55d953f0db427717eb7dc1ddabbe28cfb02fe78a5564dbb31dce1895310699766896cafc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c90bba629ba41adb5bdc08ea94e87ce00b99b915a95dd503f4d4ee3497ce4f18b0644fd9366adba1ebbe5c5591fbcc12e22043417ab7245f7f84d566a6ceed0bbb100ed3c90c84e8ce4315593603c2b3825f50d254adad3d74d5c744e3e3574d2689b68ba2f7eb350727a804be6233ae7c925c8f6faacaa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba91805043d00a4c074b03587f7abf85a8b30069ecd278257bd2696aef215d2f0507a6835c4b3011ecb0c0f557da3a79e200f76b9745953b47be896d38cf6fcc78e1cf3d0aad89e54f9041f8d0711c1b4cb69684556022e836e0c7e06325e1f8247fe162908270a5133c668e30478aee9356562a4559f2d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d612a1889ee9de88bb52a8c43cdaf1a449e53f8fcad17b2626630d8c9f3e3d7fc045a6de7cb340c10d340a828aca7edb327458f696c6e6941d4beb627d589994f36516e84afa94a6230362dc9b40366bb964ded73c134afcd4bad020e981f10ee754ee04fa6f7a1d42b22823b8192a4be0f4cfdd318c6feb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58ef1b949e6fc8ab0b66dda020634b71ac7ffb7a99b6bdf8999cead3204d1643584fa933ac34e9a85d65270820666531d5d3eaf557bbc52abc6428db565a99bdb8b33ff5d9a0daa20df493de5471821d69cecb798e96c2b589276baef4ff95f98a07eeab5e6a8075a79a700419d135ead353c9c9684c4624;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h307c9249e940cb74ff8bd201eda2a78d8cfabf1a3e3d12dafb2ae7e35cd6752f5996e8a66c66cb867a7e1702faf10a15f5fbba395768c442ca4fe02fffe71ddf766fd53dbfec8eb2e3acd36f7d9f2a0bb945e18cd893e997127a00421ebbe1aef2dae591f1edb88efcff2fa10b25f988ae56a65df3f3b4a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6d614f9dc2f72000e5192a81f7bf659ad10e3913ecd94a836f83daadb89a1f1087b192a378cda757d307c046e6f4563b4f717c8470457f552ddd73d947aac269b75b0d20c8e93b7ddbaa98c650fe898dd6b29bda4463c5d1dc4aaf3b4538942b8b2ae67df8fd4422549255cb74852a06bc3633ba13f8c2d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3cfa3eca973f7c5ebf5c4689bce73d00b014a66f5c234357c4619274199689c50db5c75ace7edff216fd788141910617b06353587789566a92497445fd7e42e78111a7c758fbfa05a5a08b0b483cefbcda80afd6e354e5591d6588f66dfe31001e5471d7a7ff4b2aba990334cdd894307022e7acf7a5a9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb953d2048f18fb3b3972daa5599b1bcd6533ba7ee7db8f72d92a4a9181821355b4b7b3de45d040c91cc9a74e846cda42198f0ec6b7ee962656e6503f3e768cd6e25a9b551d6c10947b6565804a12714bb1555a8eb1d63f20586739d42c776369018876eba00bb8b6d1fb9e79f3da09ee186414422a2a50dc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185ecc1c976ca7723c2d1645f27a041267f25c47df942fcb68dadea6966f7aa413194f91ebb7064b838210c9cf642bf34d5530a7ca4a721a7b07b44ff201f86a3e709af59bbd46dc00d75512c931bb5c0f465fe32d4a96111cb7c96f4a013546ff963e1cc0ffe7f2b21dd1bed757286f53e2dc7922d46f745;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157f9d7f25ada5c98727bc838084927632a3f8928a79b95f2043ec8a32b288965cd1152d420af949ca7173d3d60f92174cc60302e2a77962984f3df499243314bf7586d10a859183b73fb4ac59b278aef0a0a8ec00d9c6bf664fc84da35aebdc5b94bef44332e153fcaebf14a6e225a8a2c6c5980dc0ac866;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bea72927f2163bfc5e5abb41d1b2d6b331db2278e0663b731b2badc498b93fa292a67c23cd06b07f6612666da5777622d4fab4db33f345c6a86065846cb14250e4fc74132f0f951babce8f68367c65c6d865469737e136335937f1b8c6f9ea175220d2d6bdd668d36ef5610ceccb907dda3fbc8976d8296;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2c4630042fc69cc6d733477173e36c3d86257e061b737e6fe1651ccf5884e25933c076b86c37c7b7d1a63fb7f468ee26f9a86f55119e7fb0607883b042ffae2c0388c61481cddfdbaa710c778da9a526e7aadba9b83921c3815401eb54f9a651400edd50fe064fe74e58128e1de4a52064c963080d1a581;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd5e4342753b80665c8551df6a7bd865711248825b877512a7ad8a6c4088deea72fd1c833eea49e0c1f85cc97a991af6f4f998adaff7129169e99a0245f32486851f823d7af1552aece81e7949449c19cbdcfbd86eebe73ff8327f9fa6d0a97649d9514e1aec2cf920a75a880b2790863fedc0c6302c5918;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8eb9f6c780cedb22ba563a5cd6a4238ffda0a7a9c6cdc442e11d727bb21411ae7875b99c78c5bfaa4683873f8e57f996fef2d5efe958f2412e6be522728b4631c875b2095aa969f22cef6b1183350485111f1536783ae5e382c92b0d93d5552690708e91bcb5b0ac7f923ba049697f37a574c07d57aaa2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175653eab99fa221b3caa91d1220b3104f8b7e22569d05a0ab46e2bf824a9870bd5d2bf7f5ffbca749a80c67dd91444efb999e528088294f686bbc34ad483273f054e52b723acb14fd5665bb22333563998d1b14012c822535c6809b7efe24ac0188e525f6caf1d7d24e6eb61bf8fa56c99915fcaab0e4d1f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e4f40abbe0ee3f0d602a38eafec40a8764427877e18e387d73dbb2dffcb372eb804f639910f1afd1bb995a55c229f70dd84d3be2c39f62fc400e209252d52207a6ca9f227ba137a9bfe7fc830e044fd6e2b1cc2d541fbaf26f7c80c8ee8cd880338c663c8c65fa9662c93308314744bf7d7c6a20e8b8b09;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9674780797fb669c75133e90ab65c0b1c3cb829f7b8a3d19168430a3ae88543ddc5eb01543a6d38ff3a4f16322d08a9ccf771be5779586f26df1735d559822a86f145c91d0f753dc80b7bda27d6d1ef53406d9497c19f7750d242ecc9e2fabd435cb682ad9ed30dac7af6dd836ddf18e033f991c7a0f91c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14aefc42ffa72df96d0fe07d23de0deb226511b27b49c6c8293f6b085662dbb6db108bdd1fe2d258222386c027d1e17b0a281a2cc50b00ef824c6503daea7c76bc400c7835223508debb084e6661fbe30c33f3c2d9a5c6a2a93eda2ed7693eae6a712e4d6013bfafcdb6b7cf0fe939b6f3b12df197432b0a8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19af297653b67be50f52ca9094eb7a0aebce987f1b120b6be84893a28c6a1cb8b5b75c28803d680c9fcd7d7bc13339c69fe8f40914033ddb55c62523332be37784998cd67edaf9f553405010fd18e65b66272d4d2156e607f7ec15dfbd489b719665ee6293565bccb075fefb98b8345cb519b52544249a75;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1812e1c41e4837d2b512f9c6bfa39233e50dcd011209f497e7d9317c21a8ea4f1e3e7a2aaf224b17706aeb9d7a881cec08cffd5d414fc958a6c5acd79a33c8183c138f41f699039f49bd1c51ebb7e00b638e40747deeffe016841156c938219dc75d0538086cd48cd2d42cfbcf827d4348c82bbbdd0dae5c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4190121a5637f6a99fdb3225aab1dae81f579a3b19171bbd3392357e1d7f490e209ae03682fad002fa18dab66ed437e3dd79c978730aff2954269d5864e673eb379c87f933f8b0953f539072decd471064ccb047c5cd2f81bb5f13c4e1a212bb344e6e111131dc991777e76f7d58fad16d2011e0b75131d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dcd1c0483b669567f1e3c2c6294d0dbef942669f7543350bb8db4375e4ce01c9f373fa4c318d6320841b824babe09ee71f8be8af1dc49bb455a2dc71b1fb68b287d979e6532cb4980391dc0341729381c2a2e67691d98117f6b155e198ee9edcff6b63fde7d3680f1adebeeb52885b7a8007c227c55ecfa7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae506eab3df7d0d08fdd3deaf9b46020bb3c17f0a3b8312ee498a67b23c54e4f05a4261fe35677d21ae7a465a7acfd6af94a48a8ae84466f5a1d6da1ff8c792889f381e330f5a5f37b515830bcc5f8d149c2886a7b93abacc80db1941eb5b56b97fca792307610d4fb8f30530c2d09644dd4f0f13d3c72ae;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc5edc3ea0f5acf2407a7c2bf5cc166e849de93ded186b7f35ab1f838809e188281f85d6cb77a9cb43670ef8074c4a3a9d5a1486e28d1d639605f5b5181ccb42bbd5d0dfe85869f4802e7d1165b89122137b866fa515bdf76db5b0732f9727cf4a15c56d73b88fd96ced0301547daffb54fd3744fbe8b95;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c93c0522888d8eb739adbf662e0068b41c67aa274050e18d16a9ef650917ce3a1fb1567e2dedef092f9c4be93a667775db658be197e8bee97f016badf474f8f4db9dbb99ce1daffbf2f824275d2690688b16c14e000a3163e9cd602d29f7240c4b01bf775380a3122724de3d5d851ebb947f2336bba34683;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183f95e26042bf2a3766f79b56c8aa53397fb5935efcbe4eebf15c504282d5430d603252e6a10274ad2ea736ebaf99a8ce095bfe2ec5dd08cf2eebd73f534f57ab633d043d8b223ef8fe2d25c8ac9e051381c6ffc2c429a0640cc3a71de0cf71c58a1bee4eec6c6f01b9477c41f9b866c5de21f57729280cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0bfae469b641f037b60d09ca4dc19ac4ed8bfb02843864b5fadce1333ed218a8c275a8091ab9e5b9d6062bd6bec2bd1cf9f0eb4c76fe14c007b0e15120875b2e70cabf692e7405d74977e055fff0f3a611e7548ad3d65650aa34c94cf1fbb0c732480677786f05911d2764fecfb97159099bea1c8dcbb3c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a69f34014cda376b260877ecd82498c2ddac88a55d889e89845b97e49bafb70187c91d39c7d4009ab4337997043d9c21fe40479a8bed9840a6a759a0f24d3d41862b325867b943254fc8d9bc8f089670de74e190d726bb4c9a3d4bb02937636e89d93446966fb9bf97521a2063907bd55375f5851407171;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4594662f90244f7e9e2c2e5d29b6b0831e119f5ffd02f485f9e98df45e3a829628d3e845e0d4f92b759c9f2e5d9c8d7c796e34018b9eaaa8d1107002d4f4d95afdd8df707152be582aaff10288801456f59f19da94e026f7973e2977e3b4c58f595798d96a61ca37146b8d05c4dc8f518a8f68933dcceb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fbf17d729fb09679aa66c2b5412d3faa8cf24faaf2ac9cffe0da570a2848271a59c52658ce8f46351cd79ec31177519a95e83a7702112b3d665cc1aa4d92991e83dfc57da520be1919c4a6873123923ebbd2ecbdbe6f2da7330c52f9a48a081a15f838e7fd12d841908c84c053646c68d98d3a9958ae32a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8718d429e2d3c53349beeeac0609228a2369d3ac0c4b8ed44da5db65e6223500ede758e1dbb38cfa16317011325c03a9d47a368ac1004ccf8ed1c13f24b50f13c6c2ba340b34bda05bd5d9611f1a6a20a99424a3d3f5bc3fd4788b948586da1b9cdb45bfa54bc07bff5a5ba8937d459f578ebcf747c99436;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152fe2515f68eb8a9d44a7e2f76f4fbc73e91246e2af1762f14d848e5b64113ed95bd111faf0394c87c6a1171972ec211d79a073012dddada7429c47311a9edb644224dc6472243383d76446d6ab7b03b4b3d20a284278703164d4b6ea15178f78a186008c8ab16f9eb64229228855bb71546dc76e16fb64f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb9d8817dd4d2709983012b1cf3c2984150929ef62ac4be6c2e5ef85722ed7cc0963e4646561654b391dc2de44402fdc722e7c626fe69f3c5b0abea079fb90b2e2103d5628a73368f8cde8b0d372efe0ffffef4e00c1d55d54a8d3d78ed2bfdd298f774776a1cc166a782a971e803ea61cedb8f7f320e647;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13890a6722f720ca016abb8fcc4e408bd1bd92f8917d06161d2570553dcde66f03aa90a1045811673c28a4abad05ebc275bf7a8f41afed2972613a47e1d6fff409735429b58169bc4fe67888508febb60c587b9481b61dc9526010024ca11bf6826e29fc24139d58f628348c453d7472b836ab7ec5d97da2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1955ba4e93ef15c6843e92fca9fc4c86c04e457147f7c314da5fb8f044970c42b56b22ad94918d0cb447e9d384a1c2fb32c5e118a1cad39d1ae2a7dc0c92f8b6c390fc19819fceb70593c5d8a93dbf62d2c01ac085d8c0d8eaa12c7e400cd02da1f840204caa5827236c197286cd441e321b6fd7c4e71d122;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8049178ef04d63e353c7b7b1a92235bd6e4eda1558fe1fb5c3be04f692a2c902234bc252ac45faa3da42201d8bfe9473e728a42d4e3da9dc65a06a950fe837fdef3d744d1e82051634d3899b642391e70b5e9d8dfafa1dda05e9791dd461029a5aa20daf3f3853e1add51da074cde7545ab5d0a324aaffbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h419165474c295a7582c8b8ea33dae2f2b57977fa55c68833c759027f56f211a682f1685c67b4215800458371d3c8a21cbcb828082604234c9ca13f8737db38f7c8cf068012f73916891d2322d74bbe67bb129b842b968de37c1b8054f1e365b53793657b5dd6e3dcfa1f8f1c0932e097bd69d03f4148f2d8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34ab49f2de0bbbcdc780a655e5222468ac3dd928bc046f19c5fd4baac7da207923fb43fad2c80649b58a40cb99f7e34e01f6666a058a31680d667805e388f1854aeb9171aac132d1ebd31f8bd8c1172aa7928c4d4ebc0a8fdcc40494af8cc968b9a251cb599d567780025ab59e4993132a83bb78457d489c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36b30762810600420af3470b59184c5636d2d8773b73ef8a1b188b5c45ad06710aaeb1f17120a766b8a829d9024856dd9de67367788b84025a9823dbd73ae72d976769a311d92ddc53cdb221994b1278f4c6652d3d56a352be36cb43a5db4c0c3fb97dd044ccd35203b98ff63d392f2a565880817d2650b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192d01da51d1be641ff5986b05723b56697e2d7d19241726d057e4224c6d0d1b8ab7558fdb7519b73ee0f664c8ec94d7c2888118ace7defcffad8cbd9d2881563da9dec1da03ef44cba58d2920242bcf7eb5d09aa2a8a78375846567a10a2059ae253b145220dbb8c400606d28bfe72ce2e6f5b8aaf04ac0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9808ab4ef3f75c0bd311c04baeba58e2992b0bcf7a22e1e1afa276cbe451881c410335a601b0074eb104711f895cb6d1942abe6d8ac723e77b4a626d4812c9a2877251f5c92963adec6ffbe16cb350fb64c18f9c12d3a2792fb8a69ff8c5830ae8832a968d2a36b52f69f7c694a83a3e61b6994ff7d3e74d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd18fe11cce37c896ae3fe15da3f61c4684cd5c380732312ac52c845022478ab5e9cea8e9cc29bb321e3bdb3453cc0d31ce99f8cbbed918d896120123a90d0184de24ae306863cef3c76cd0e79822f8d7c371a1bf4c9c26fd9a1172bb60df1d62dc90b8670c74eaf24a88ccfbbc58600fb44673035b5abb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7bd45d07e43a5c0c1df2b078115e199073edd5c80b341efba8b631522eed947a3dceaec5a3a0b33190cfad9d58d822d5a2e1944855b00e0ff5211a6dc78aa4eb0d29bf06eee27589e714d9a879ceb35cca5328ee4d5cb1da22eac5caca01a362e308f398a8ed5e725bc1f9636dc0ddd2d5518cc1aa744a2e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16844e6c472cae3e2a86f36f587f631d24b130fc5d89af23ce030b4c47a86151be8c097e1717dd8e452a2df6fa070e2a46e88badf2f190fa3f5af669bfca47ede54f3a29abc7a2137fa09c4cd53fe294e7f17b7bd2ddf05254a41a0c27d1ff97273f4beec9a609f0bc4d74620425539afa83b2fe659e04472;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2866d0dea8c441bd1fb1dc467c46e86bc5c6b201d47f93aa86f5e063e7e97ff4c721ee45ac799943df65e96d8e9203d96522e9d768b219ac33d555da31790093d4ee5dce72f29d1485f839ac310f2a5046120dda96b5813b629f9e717831c3287560e7a5f0671e5278229dac053177a0e5700d71401c1c5e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1499df4fb0e1ddbf9c5bc6fab9234e8dd59e4e08b730f977685a3c1038bf69f3a453855398e29244ef932c2b6b7af93be131ed404176e073d3490d2ef355e17f104a26d1b5b070fc4afdd4f26b86af3eb0d6f7e3d2138f319dd2a8f40e8c7efc0dc1ba1ede9de9d1c165179ee5bebec06780c9078c919e183;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h738547732e882e9345b275e14e560e897f7f16c312d6b1ba2e749e5ebffa2f7301ff829175801dfea07ae35bd689aea840c5b4f6d4b86159df54ac87831b376bd682c0c6d106273057ed3b1825c3eb4660a75ed924ad2b039530582ba2b46d4faa263518b844e7ff996bb5843630c7f4e7def8aad8a411ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc6ed9390c4083f799480a80ad548dae365b4205cf37596d519aec409f751eb1608d19432e511e11bbfa00edbf2fb86102b891d38cfc662ac1357ebcc9c1b52b4fd1447fd6a92dc1c57aa7407ca1331c667ac47e6f1f7aee46b824baf5deb2378bc2b77de61f8b1bce609660d233caec4a80307ce2b0cf5b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a89b512f7741a2c62204694e46b2f84f930be55c89ee28d465c4f11bcf18f58ce2bb2639ce222c03ac07bf8eb0ddb3de42879368f9332cfcf93851378ae19b0dc4144581e1aad9bb4b670159b231aff3a12fc4f1a2ec9e3f6513751ff6e1bd713edce9773ce56ececcb6ea9037bf7f983416135de07c3b78;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1164275f8f0dc10f2b90a9feeed9b9ed6019b9e66277accee34064590e052e94d705d5db01e8a6a72d0b146ada887be54d60318f7f6d9cf284455383a6bbe6a4d3252ecdf077625087edb9ddcdf817f219e0fff0f41373ddd42e6f85afd5e1db61246a680f37013781f56b4f0293a2dc1374eb19061f0d3dd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10141a276a998330d72af8b109c3959951e5eb06430de7c86ce7c57ea2ff93231ce65acbd7abf081b461623d5b8f42fd3c8244ede92e28e9ce3edc2d47913691c36e47363ecc5cc64a6e28303d8994e9360aa60adbb164cd5ced39325d7117a4ec184cc5f0787372e7df6df44b1594df298a1f69b572c9352;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ecbef9bbd7cb27d8f34a7f05f28432b4eaf311fa20eaf0c268436347ee8500d4a906ae797d792f9e516d59dc3b6b5f624d9613efcd8afabb0313bffd01e890d2b87f63e44c68110c66938add4961cbac9003491f7bba146779968f275f6f06c40f896898a3b254b50c09b1b4e1ea9d2c313cc7ec5a07e61;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74f5309f8980eb05ab49d177cd55b1b47f29a9451a844b58611b34e8945579de2a485f007778622edd8d9a9eab2928c17e0408ef057639d31e267b896844a98a64d5400e16ddb385257e3053db3bc7d79791aa85392809bfb397c1ab81dca1c0c284dd71beacb5622513d5ca2a7863c7d65bdb669a37ed45;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd80db648629fde12c7d76404f4098d90c72709cedf43fb76ef10b88ac878356510a18a670e5bbe78d04f22746e4033a2c075cc1f36333e0107dde9bf885a9e48894339e6efc9cc8d37ee36fe4a5a2364502e5427f08c390314a231e432ec63dd71ff61d292a99517f64d046fcab5855b60dc941778982d80;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7414e9021e43e49bdc1a99f485f4585c519b1fac4ffbf4e452d766e1f5d952b850f540ce22e3e889258a222ea0c6d6e6237ee70cc3acaad01ad387a9f6c16335040c270c7704fc93e6cffd333e524a6f3061ccdc8d42c111652b7a164bb2fe12fd1d01891137f8c91eb3c983670a074403b085e74a0a12d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16cddaba4c566ed8d3bb31418b42dcf7831f439b8f86b5ae26ab7cd66d2995a915035c8d86cbe4fb603178ce24e2041ee4b0e6ec6f8f5c60ecb5ffcb090e94bb781dc8569da4a32d5324fa39ac14cf71956f648b1965897fa48eacb1db77c315b0c0833652e06b92b036ab8c0520a66fdbd39ebae40eb72f9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafa5bed8474257c7fdbb1e6ab94c99cbc4ddc43bbb5d933d715e4526d29a810eff8a7f33d8c63625a2e468cdf193b41868104b0fcc8666724a9c035bbbca6b5c5c55e594153d83d87b52c60c4fc41ca42de6d076175db391c4298391f0db833d58e99bd4121a7888d66df0d6d40ad617de5ba929b1768297;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfbf18be60b6305e02e2c0db196954009adadccb74b150ab256a97eeafe35df01778a590016046485615a52a3e786e6bb69ebeb3557e14cb6a6dea8dd3d0735de20b2ed7b520ebb5849f68fcc7576c942ac5e402311e16690e08a6d3eac5c13452299f032d5e502237d3cd3f193da0e301271053794c4e80a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f491679e01812c85cef969ca4f79fce7c9cf95400ae862e9e189ccf65de7736f4095e1df0d37f63dbead2026f0ce3932399ccfe33fda6024d1b21683154594522bec07582d771207efbc5e3c1939822527b20d1847bec386f4b66037d51204557818fa9993267c1e231251acc72e6ce149a657ad1e52715;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc3eb39cc49bfa1de9445b03fb9aadb1396423a7d11450ab82dd25cad17525a2603e55169cacf66e77551a33e2b753fc8f3ea06e9ceb7610d0f1fd64d96e1c203f8d784cf89d4a68954ca4eef5c1515c1008b1b9e80ac96fde85d7c3ad6dfe02cf618340f3cb7b5acd8158a200a15acf0154676c25e830e5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a1d2e531b932668eb1edc1988a642a3a1dee240e3f3ed78580401517186da7e539e4dfe0507cbc019afd6c7638baa370ddc73804183dc0d643883ddcff7af7e1de979f90e45db7365994a24489c2481bf6493206e85d849a33fded1e7948eef7a5f18b10cb7e6d95cd6d09902f9ce4f6f211340095a6985;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eba8ab15c2bc61acbe6e471a96a39e50779bf424fe189cf8d9843883d0334a6783bb14f2bc8f78032d8cdaddd9b38f4946edc704e66cceed549fc6ec1c00447b0d7a4cdf680dbc6c46d77ed0fe268643d57a19e5211214cb1a0862711274d4a15b130e0372262841f1f8c43ea529b0ed3e5d67fb794dc489;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5977e91151d085c5564aad6fb85bf6542f3fdc2c3955940ba68e9b1814a1140e8a2c90f96ba1c1f0a243d74fa628f93a6bd67b0172a175f01974d6407765dfdf6f8238d17cf790f6accf68acdf80cceef5d0ed3db123fb473cdafd7c0658e7de9d6aa5c2042c7d39a003bb7c7a792f60a1317754dcf50b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d5a7f1c60621bfe07e0dae2d534ba4d56e12bc91ef022b26d5aee49b119a7dc2ee90648e995281238707c19c9611b3ddc49d5c3201da54c8decf49deb927dae2e73a4b238d8b76b4c5c9053777538f77b600e43ca36c220cf4003f7a748a0cd79d95aed2b1c3e1511f1409dc84fcce55a1fbd1939f6513c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15cf08e12dbb2a24589980360369df36444abd277e21ba1a9974ac666be5e54333b8c191a8947ba72350a0dc186c7057b6b84350b6a6bca5f7773ce4d7212db36de3faf42ccef127aeefb1c09cacca839a01f15d006bb92a8242ffb25cb9b2e24291e02a70a911a4e31219e086a0015d651d8dfb32d08262e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b42ad52d4daa547bec110c118ebc15a4d4087022ebf7e4091541f33be0896f520078fee702eefb6036c3f1e2434bfab170353895060c7d00176312c688a97dbe4e58980824346a93e1f2fd44095f27844b047b1ececa82cba7ff7f16e24bccfdd06191c75afea989a81103a663405ca1953ce5d49dec912;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67fdff5d0cbee85fae64831ad3e036abb8d75ef994f1c5ac2d76b2ef599aefbec0f29c100cf1839a39341c1e08eefa8bd31f612c258a797012e69c5408c7cb4799fd6e893f73270c99fb8a1eaa593b7471eaa27b07989516952e823158b395bbd76b6b6c3aea3ff252ea455ca395c58e2eed0eab08209ebf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103330c55eb8e7e0217c23c05761f12b49261a554de6f16dedefbf67b538b0691810255a2d96499290f9178a7946ea32cc5d95f97f88acf50120b4aaddc995fff30ac04e87a2bd754de12a2fd73e8aa646dc3ffecf389dff574e26eb71bdaa9d0fbbb1c4c1c43fd805e75a4e532d9e584a6bb8ff5b2fe0041;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd93ea5407d9ad80e825bf0970dbb5fd87cc3afe20c7e5fb85ec1094cdc31363b7c3ac6ff9d8d6c3bb2a6e58a1c30e2183c1309afa8bf97dac733d43b8bec4928f0c2f9256ade2caf9d77e024e33a1e3d6b57369a06b341c8ff9bb12bf44957cb021c0fee1464db18f3887ad9f68ec24794701662be864713;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14981539dd8a796979d16fa3e27e62ebee28881817c94739d382411cd174e07c041a31a0349265fc3a02034204ef6a0ddaccf9e5c85a93c70b5a553150e5c0e3f724c7ae2b62a37506fd121faa69a3cf142aab3fd11adeb6902d02b5db9175d0a7d59be7132514469ae6b398a0867530008ab4a98ae1de3a4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c2fc8a69eddb8a9ae466a519e49d1316f7b34cd877df54db0827aced6ba51c248934da67b25843123f14061214795c72b08a515e7aed019773f01667526c2390c6af5642facba23038191e0ce57e0287e257e0a65f9113ee827fe5e5b549ebe73c27a2e451b62f7691d8a9255e957511b1a018aeb83d20a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha805c029842689b60c3049780ee9ff4493b9bb30ccc50cff8d5080f5567235cbbc5c70480fdcb0f518ce7fc306fa73256a59bf875fa992ac0e51638385b46957023874eca828e60abaa841730445ffa1302d1f907d6dec005469e553280cb9593a023330876e47b1d139b909cfcaab0392f66c3831e1d3c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126ac04b23745b001bc65f59aedf0a997fb3b57b3700c87f869ecd2add137d86ba97ebb96eda0ccbfbd065d0ccf874a7ae65ae690506c8c8a3883f9fe0a20c83c33ea0e0b5617b9ac19dd0add79460ee1cb33b5786bfe441d5bcef309ef77245e1c3bad3ba6f14bd8c841b59838662c86c189e90ca40d46a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3a6849c4ab4090e546d80e1bcc971ecdf3d72a49228d4b912c2c7ee4f22d42ae5868c7725ad0b0a2d84b4bdd0f1ed1c6da9fbada065ae6597aa3527f67323d0d326609318f667a99cd6bc254b2d62fec2ac8586c5c4d85e1ffc24902b4ff6703f3d0c6187b75a03a146b9b80514bef493c0b49610d7b7f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19964227baba72d3084ec622f1cb307109de5c59d32512fc6d98ce357775e84c5db60b394ebbb4e676526a4e9d4a3224950dd1c4873fcf507e73677d0149c1ecf63061aa015a2cccc898fc49585d5562f5bf0b54fab94b3e7b60694872a9aea1dbc99d89ab40ec04bcd71ba054cebadbba59ebf4e4b737be7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8485677c03e162abd243f52de6f285037382cb90ba0d67f2c54aa31e49abb3c76d5b3df152592cdb7aaa4329ee342c0a9ae8ed93e74c97c51862dd6eb82e69c68377f876f7af7e1b38f161ad971970344d51a2c0c14dfe867840e4337e4c8f64ed3f573b7035a0f323f020aae2095b5f4c7fc80632377c2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b0900b3072448dd1f9257f9b2f5236ac4e1edd88a3af7cfbccf18a91ee2ac0c34629296e38288e35b983ca0b0187a18e30f008f948d2241d40ff7b37f5a300c184e2c90465eb88de77107a6bd1e8be60712d4a0ebe44f2a592cc227def14671625b0ad52b5a3621e359149ed8b2ebbfb817df25b786e42e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d41b08700139f73f16ad36d8fc6d4ae196959b9a4a5cd0502c051626b4b46ca2575b58ad45608114970de1ef42109f837987ebf6b42292027815994000d9b2ed4ec9ae71f07f18f8fc3f01437b46bb29585e5eebb7548a8a99ba5fc5411687c568519900bee590c835ed903de371616de9692fde4ee0479;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfe64e6aeff20397c52d4f5278cd08a1aa8080c904f11c584f2a9f8a1af32ae07164fc8a8ee1aee9cf7dbe55681a5e08a3bb5465ace7f9b85f479f63675ad8d42eb46272ea443750fb96cdbe13a370b1657f478d8aa1f536c7254608453718b4a743c985aa70bdd4dd1c902bc381009cb0e5ac74a30c6240;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eff600edcf5a938aae04f4510db091ad132fc198b5c53cd1f5a69f0e0d93c865e74df7fa7520d843db6b2559c63e26ec34e1d786d981d9a18a4ff443c29b7c63fdb6d44216e07e4488adac75f43f9ecf73dc208653ef42c38b1fb5b539369491127e972211e32ebf98b3d8372097881808842dcc9cc9e794;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43586bcffb7cfe596d5bd06d94f149de6d100ff8d5e85aa2b904308b7bf5ac235e7ed7ab7c77836f9ca892f63b1504ac67a497d6d6794cc4301cf6980ab4e4bc173236d6fa56ce827e11c6ba055ca12e4423832ce2445a1b4a07c13c12afc99ab5d3bb6a1134779c3ca3174a3f063f5d6c6ef99e5633fa04;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1849c60eeaa80b98cd456f17dd01a6ffc4e2f4ad2bfb365dda1cefa507fc9323e61c58a64d92cbc3c8030342f933fb8e8422bc070de8ca9cd25da34793f76aa664437fc896b0a6ca4f9ff881115f61fa5078abc489727a29a66b86a0decc57a0337a0d0cd7d0eef62ce0ba5b56e13f472c9a77274bae9acf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c670b042ab1e57124e88c154e7f1a8a438921b5faeaaa71f5890bad0b0539961dfdf1e647a58114a278bcebcb06a904fe9fb71e94ecebc2f7a898907b34fd5058a56c19217cd977a49b8d98b6fe75c6f5e1e474a839a8c7a22b738ab7d6073f89dd13f9f677e684cf177f8a12d69059447dee66f66528a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5596bd46870d96b7d864b7d1e91a9b73c12dd45dbbb1bb5b7be497fe5a3c4499925d4cedc2f26059dd78c955d70b937f45ecdbe449dbbe881505be69da6f4dcb9945e52e95154ec004b3e83f3beb2c1b361a5b61c039fe84c44c131af9f4d8efbf22e6e574430408b28f8f11d0ef82bfe3bdf8ceded80941;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha503b34e3a975c9ca0bbdb8ec1d4e9303452fed3c58274c25c968bc254c027d30396f9fdd1dc3063df87fb81e217e7cbd6c4d9ee5e9b3b51a3300dc951171a68a53b9018b04681c9664f1a675173c564b1a8cb70614d0647da239f5e6297ed2f1f031928209443ab16a8d646c24f9d74c7a5090501b1d6e3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6df1af9ac7425579721c059afc423e920b00d048d615e676d4c36ddfc8655f724281e00bbd623ea914247af161fc6b34d8ac3d3f991cf7ab5e750bbe001acd846b9d0a74b2dc8c870d004227afa30db1f13df5f369d408198c1c7a39bbf6afa6b9a04aa5910fee3d630dfc9f783fcc22b3051f3a8b11154;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bad27c5145d1b988461840c5e4f77b6a2a4d60cb66f997e5a59aa62f65666fc50c9c6d48e77aaec88a7dab72c8a41fa11ad80151f98e67838e74982c2b57dc06d4a1d8f3b0c8cc2123b66d026fd81509ca446a0c5401ea752c91148d5cbe31697505e9f76e1553ecd3685ca9b5d3d6696548c0b5f6706c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182103cdd3e43272bce1a8ada3b9280e128ef6ee4731260580a154cc1c3ade9f43d00ab6262ec842b0cdddbc07f7049247ce370eb1845ce7661a5c19f0983b3e1be228b81c8f0944a2ce7d8f9d40d5e8839286739286dbd43be2494293d62fa1cc9a03caa7f407607718d753579d1d4320eb96d7f0c7eb63c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h101982668218156e7f3c98a62e139b6f77a3c25e548d15430c6d939bc8d2d15745d24ebc9fcd4dfba7918c47950ae7f097e0aa61ba7db305d8f130960ca41e396e7a84f5615aa726d3d4cc262b75444e60b7e40dcba92a757b06e8ed85c766a046fc093978d145f1a084f22aa5dbcd3884a01dc1cd95194bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e92575b5c007d4176d496088402d7e6c621ab628900128b7b1739545c305385f4c114a0cc0170b7cb9e76f2b23fe6d2738ca7a94b6e83bb7437e311386bcfae3444735f3e708b7d97765558aa9362e876acb127ce5f03c1839702e7a9040542902b2942b9b5db0683372b4eac099fbf988cea9f1260fd5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1640f6e9f65e995f82b2c7ce3c5f6b1cefb8aaae053795e915bdce42e5933fe1b39a3ab07299cab9d4ed4569e35c213685ea21692f223b52fe249b70b3d58bbfcbcfda8550e9dcd8417dad231534ea124e1484ada402ada87212994ccc871bbeeb6cfc27c57d366c72e24c1711e746679b24efc42ef244dca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13274c6a75ec6051e87233df875439730f0fc5695ab1b28e5309d3b8d70587367de42e442db3851862b03a7f6032d1f7ead742d2089854e82ca83cbd558ed65749575193bc8c7d7a1d35b7c7702da2349dd5214ed2e3631653dfb7c59ed6ddfb767e691db319d578935fc2e5e3a8019c5f9233ca9185e4496;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5c519d2086dd38e4837c5e9bc29d18147540bffbff158a2962265bc4af9f362a0930fe871a88f3dc7ebac37e0e34a2cb60682e1719a1d07b5b90e63d6b20654ca2013cb4ee0737154ff31f4ceaed1de6cb870b26dd33111af44cfe95e1e79c9428ebb1c293234c079cdd9ea90e566211be668b1e238b8b4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc3299210e6c0409ef617cfb0dbb72a8fde31b2621b24f49d445b9940f7178b7507eac154aca5d6016094c6f8a4c541c73695f7cfa531117acd9488db24e31ec43f02b844df07f497d03d3c3c16965dd7668866ed33b7b0dfd3b531cf6834d4efccc500a0fde2bd53286ad914a19fb338a85d9c6cd6b5d00;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127eb78528cc4050b50889af49d862461c39c5715572d8b24c522631cc79c88be364d13bfc11898e4742814be189ac29632a6a4a100a2ed8b7ade04a564d44090c64a3e5f82bfeccdf95a3fa3713452878c13060ff2059539bc0219c40c941f7f81f8a5eeffa6f3b63ba12df296ce85672bbe7e2169d167fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19923ecb705fcf35e7ebcb34ccfa9977ec32d3deebf17e3c9b4396b45df70a365187b37fca44a6cea1626fff8aeec8d42775a34d93d417c08952f89a65944725643c0c17e4236bde1307b0053dd11f478f0c3e297cd3d4905af4e6fddf72823f2641863f7a1e3a163b97a66aa3639aaf99000b0507073ce94;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c46eef7301eab8cf80149a41c66c0303cfb85ae51361f4d08373ca8d5fdc1aef5f10f4fe61c420de6273b46a62c5b47e06467ec1d45852648851ec6b82225c1d3f4a1b0821f347a479ff4efcbda094566a0278b8708739e7c5bb921b5358054c14afb7455924fe1a7faeffbf4c8286f28979c1889fb21854;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1304739b23199cf62d2b9be74b214e2eb9cf0c8f2a210f81e54495d0490a0ef48f07a01fe027f055a2bcac1efe349c2d5649ccd49b3a69daaae88eff30eb29454058d08b4a190cf62742f20de86890751757898b410979da650c25c9f8dcb9c904fd4743342c61bd373c79fd647778fc2a2b768b1b43144ee;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3b5698b768492df48b82256798d9df8612eefbe5458cb2b0954f155050e4af3e4987683dc3c43dcaa8d1fcd6ac5965f005c4a79d5f3075087a47df3b1a8ee1c0857b459354578447947fa133cf62e6c6e5a45b5e147451fefef6d135de1cef730af09788615ee59e892d280bfbe59c41f97ac2a2b5df3e1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f36058627b3ddbe5695578e56bc310918db636fd2742cec4591d851d1b37f522919f807219e200b807252f28e25771dafe986705fb22fda47bd2d533dcd41b94c1431534ccfdb0bd1e807c3af9364d2a62fa8e5d1feb62b81720aa80d15a37170482d8f79e3c438eed73688c3085a7f5a1235c409a4b131a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h248acb0fca54ceacff969b6f7521b1785f1d6fbdadb58d197fd24c3d41c46989e8ccd3ee37254b2aaa5cc23c529ef415a15e9b55526ad4ae728b4ff7b2c72cec44a89224ba3e7d40000ee4505bb97d76836dc5fa322a62ce91a0c7fc5f6e23ca8f543bae65f47df2d80d8885f1b08fa8c788684cb2c00cb8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4884e01c93a37ecd5730a286fed5e903d112314ef618f2cc2d28c8b0faa7749ea9027859faa3b696cdd05961b2d46d5751f86bfb6bff0f00439cff6792333fca34fbd90145bd2e5d3c7ea9a326b206f1052a9c27496f4a15c4861a2e9d2ee21740edf9b597695a90c0271231165e8ac6c1dc18c99ebc7f1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173b8b1b19954aeb415baca4e9420f720b83163129a52ebfdc87a84c87ba9085710bb2e87cf0ef6190da68e398e022b78aa83fa8fa1fd3090c156cc61ef35a94f8c2c806068a5cc4fba3a3477533148fe622bcfe17dc4f6f8493dcbd1b212a2a233f7cac6334513bb6aa6d8f0218b47baf2235d4c1408cd20;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e8db0925b7a151063f001f1ba47559804a40b059d6375c7194eda0389dfeba054e765aff7ab029016b7cb140ec9e57cc6d4ec28c9db7f4b57ae03ed179f8e8c5f8e96415909a4d23d32ca0bdf84edaa4847536b00cb135b7792304355a494618474c9f4384b5535f54145d2b368b4ab73a44e2bcb4ce988;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hccd517bf331013fc28c341ac8dbd02a08f97e5180bd03c54d910a3f6dc072acc81d23188dbfae80654a067b4fcbe8bf546ce19701ef9552a6e85dbbc01be81a17a96702ffb485cbcb84646cb670a76f4007fcc5291990bd43e97de70f2957a016423fbd8db2883aaca617225e1709c260f44ca2d4a86a235;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b00732e639badeaee5e4460a12111179e2cfe15bfd87792918aed79f1d7f4b43538bcb0451a8bca849055f39c077c5a22818b00c010467df4fc8667b7701f1a5ce91901e83e5c9ddfaa6f76dcb4b0bb795b7a88f94520cacd3ac2725adc44cbbe2b795eea04a92373034e5a1be8e7fb57d0c54df751f3614;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa50a69e814bd7ed6c66bf54dabc9e4c017dd60b7d9349e1ef29176e441d8d1f517ed78aa5b9167b68ac611676007700c59f0babdb28c54fcd843a1a822a47f050b04848c0a7cb17c00e18a62987199d7095b9fbd85e3f168f7c17d05ec8e4ac4d55caf67f3e33fb88d118fde89b4d13b82c5804bbb4a4f2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c4ec2717c1a78f22c1d9a40f58ace7da7700138a4a61b5eea9752c4f4958acc7e1e7ed70b351e4c84c310556466b58a3cc53c51f2ab7e6c089ad2f5ad0780c2df49f8d6729482aa0b5a9262301c91044bd4e7993ac4202803b9957505c64562396e502a44b5d0f66406d63ee2a4be9f6ebdbf91b4068ab6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10463fec7a79cc35b3bd3f0c858c8c1f59f095d4c0cadf076c9a947a90cf7df1c6d68291b387451ddf77e1fa46cf76eca2e31a0149551250b859ed292fb9fd53bfdd90263e043d558046f6038fb4374a5cab333ce43c1175a9f15aa131709130cb635cadecf00a45376099239f7a8b006575b0f432f27bab7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99e9033b0d874d5fa393612d07eefb48e68aec1c08e4cc5f8ad0b26e2cc2b86d98d1efdecde2fbc5139fb1b35460088333ec0125c57b486fe79935e44764f2b1c3f94c68bbacf8056abe665ba032d1b2002f562e56f77fc3c05f64e4c0fb58efd9fb4b0e6a483af3d54a835ea57b1926182007735cd75fbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h947a806d2b2565dde634bf82a2e453fa4e15452115a5f7131453d1c2ee52f87c6ba47967eeb3d394ac2bb1314a53b07f5d54bf5834ba196346ad33490edfc7d98fb82415ccfbb6c6bf735bfbab10bff2fda44abdd66ccec8edae0d6591b9a5de224fe0c5a768b5658770a2d92297a45939a35ca95e6d6268;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb183084607afdf9399551b1f1fdcae69412a5c9393636d893930b55aff861232207b19fa0d29f4ee53cabcdc16e1737e4e1e727e5bd0dfe05fb933c8013e2943d6747949ea917cdd4e577685a15fe59c7dfb906cf70a6b0e17c8418fdcb2c31c798bc60b931235a68fd26b3471c450016d368fcb38be334f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14279c38f45d222bc412a83f3f596e959e0a64f137631a556ab08647919f531cebff290fa16056586b9d43287b91632255ac2dd389352466af19536fad2ec0cd946d33c197a761f34b2f23dcae146ad75d1ef7fdd9a1cf25a7d6523706fa88c9058bb43646987a1b494b520ce79056a8fdde592059a9d3e2f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9ba19b312fa6cf2d923f5097876222c1dba18bc174fa639da275427fcbf6da46ba9b90b57647cfa138da46847ce17fc5a662c01e60738dd511f4510c72a7fae265e2f291d7132cc8a7d5d97ae662fb4caf6a2aa0909bad740de09ac57c8463f14fb5f1de58cc3ae2493256b4d72446ebce2b558852e9352d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefffed0c20d89e7b130ced04a13672feb8e5fd6705920c24f69ee26eb51cbeacfe1324ea1a9e13fa58f12dc817a2dea2ab40cd424c1867086d8b3f8e9b67c915816cccfecfe0d9a5db934355f0ff452e317a5f257d4376ff03fb13ea55b210f8e58628ed902240cb713edca704d7fe05b02ffdc71e9dbe2a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57cc2623e41d2657270b1e70c4384f8b477f7bd5c74142cd52d2798b172eb3029f8b6d90c14c67bf21334b804375761d0bdffd7722e4f64107fc7f705ca5f1e74cf941d7fd975d16eeb04df29f8ac9d0c0d8114b4f422eb12532780208f67517b2e7b45ebbd11a632f803748d3f4a260ed600b02c7d85828;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bf1c9b049644f843899768a4417a3287ab5b73cd4ea9b2b795557195d753901d68b468243b70d054597d9c53a577585d1cec7284f23eca6737af406bc578122bc141a5d0d0cc9fc85e5299031a5b9cffa3055fb642a9b4db2ae53c86e443b0dd34eb0c6da833ab74932ba744498e8923643b3047dc83beb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heef4ae440e2791c8a52cbb33eeaa7953598cab7e7c46c3f138cc89d94650d5092345186727939723fe21e9ece694b53fde8fb2f44b97a0467f11df09a5f8a069bb90316de9ba4078aa149c6af06a6bfc2ab94f84806f4f28047d3df900ead55834ae1e830021b0dde3b67264ae68a5ef278a7dab91301663;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7e4c27bed53a9a41de0fd0ec95e2199168d1149523aad027f7e9814eb3ec64861bdfa515aef6f20182dc6f274be1d98144d06b37712a7c27fe792c3081f87868e5927176de0808161afb807ec8089484546133518b2c2611ff7e83be79c54d2a35ffdc04ebec2c7b8371d0f1e88da81b8a13806ae114321;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a3beb6ca5b93614bd28c1c9a065fde91faffb5646d8bd836ef4ae584cb8333d0fd1fab3718502c3266d732704ac7b0342c731417d5dae73473e644b5bcfd3c2522c16e86da71d90efdc9584367d836ccec174d4f90f4ca1af5f73c9154e61b0d7616cf846250d591b3f6b401befb0fc5384a0d81bf3f1b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f2e1e0176579e0b77f237cba089fdb24bfb00b456b9269f47cfe4e6c3b9d3fece2dc27903f4a998fa13a316dcb52f7ce3717b3ef7b169b9d1509b5da5057a95245d62e420120c120a313c37f46ea9d6ea07a7169f82b5e4f2ac128199a28b4900fc8ce3747bf1cccca0d9f47b697c62eba50c6c86a35b86;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f78673adba28f50bc2215062d97b5b1637b8d4d706d40dac2ae838667f51841f326aa689b96cd9b247e2bafdccde20bcf1742e457852944b3d47a205135127d2105b49844b080614144dad7a6f2e3363b879a1b89a290c6dda9f28e54f184ba804cb5861e8dc2a863037916ce12dda03e399f45aff003336;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b13c5cb602fdf4187f720ba04bec0a8bb217efc8a99908ebd93886119af8edf95402213b9dc497914a9452ae869d640f6cc726e2210fa00f9b35030cd8b5f16546fe30b057090815905270a4ebfaa61070e08844d369103c86283958152e8f6b3170d6f0432d3bbc24cc9cfbcfaa3f8c7a91f44076572ae0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f185413c64e4b7e60a089d9541875b45989aa033a042cf98d1ec4723ed82ed39bf966fb00c23fd1832494e887c275281c384ae357bd3293df83fb946fa1fdc15c5187f4505ca322e7cb0859b2ef398ee2a0b62ee45b3ca0dea1bc0f91472484ebc20aebdeafbf32fc3090c84be17a27a42733f9af76ef12;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he09471973b08f57afd7d80d72babe4e290007019d072ef26b9f7cf65e5125154832fb26d6039d5b970f3f35af343902409f732bb6d4e7802bc4b67191e76735463f6b22a7589f665f5a89dd833e3db541e0226fa0204327c7e95881409d573a0feead44ed9877fef689893745fd83eed709569fe48283963;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd5d516027b83207c581f8f11e22c74e94351f94692655ad4af1a5896e4a70bfeb7de3a514e4935cdb59c672b1c82f61b339be444bc9f4a73888a5a477a3436a12e64072e5071a3ae29069f2202b9a2e5bf643bbedea0db5a44413ff1261c7cf7a864468b1bafee4c200c6aa856e68674a5abfbd8a8a1b63;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c24abee71e9fc6230201c5f2504f5da65abe4e922bb2d57eea869c6bd5e6e1993e43c23fc3b31d347407a892c01db707fad81f96d85838d6c26f776386e014120b10f11a0835f79f9fd03a6c6abd01fd49c844f4b99d735366dd402347b0cec8ebfc9096d296227ccc5fa92fee707b627895fa5dc9b6025;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77931668d4849689a7cd490d0cfb6aa6c1d84c94c59baf3cd603faf605de799b0153a156f9fc3ed1bb166fbc5bcd9ee9a149f7135f0900785c3c17786f12a40196c1af5ff17156c88c1ac0f68852a0933108c9fa5233b2690fa47c7f8a3f230b6b32ebb634a2acde5e7c0552ad49e001ee2ca845ad1205d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d159a842e26cc03b29e888cb276c5e7a723cc8e9892965b63fd29809640d1cc6ecdfc7b3678f2b0a9ab6c88aac19e6bdcd519478459d5d252d26e45955085e0b906cb0065618c277c3323e36e638f50a463d2067b952872378ae4d79f4650773277f6fea6b8642909e7281574a71b264594a917c0d4ca673;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111ad131f757bd75a26cb90933baae1d06bbcfa627593bf5fc4a2bfa8c3c940da12b987ec385c53db8c4ac52bf5497b93665cfddc82413cd901dd3ee281f7df845ad528f4ee44f73912a11f91e76b434680f16a3aceceb12d417ed5c9d5b1e5907c876e811bf16cadc687ccdfd4344f133e3cb58b10f47646;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1404137a703ef2b30145faf074228975b025b86741af5ccb6b5a7fec4e02d48e3197716cb3e8869d9cfe6ccaf75b39a68aec176ff9255ee8f326c5c74c91c6f6ab6986cb7ee7afda58d924b11efc0c78af2e003386b4416a44d0e6c3cd57fe1b2a3480be4a0b80698bda42062e36703e84550f686c4b5e050;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed82d4d9c239b210ae02e17de666cb94132855ac12050245dfd44fe77b54cff6cc4193b7a3602abbed29eb6ee69cf5b95e996f1ceaf629fe7d15e06332067fa38472b3b0e3ef1638ded25aa4f216155470123b82440dff65e7e3f6e8becd650780338e5aec6c32441794bdfd5c51a21fac09444f06f8811f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e9aecd4b322218c478b54b36e42dc1855ad0de53cfdea96c15f0602b2d725cc37f9ad2273db6df5a084e402fc56dcaf8174e267cdc72b89bf05430cf34f56e1a224c0c97db0ca02ce259f0db109776979f20b0f8868648e9ec76a547312a37092fa93636e5d060100d7aef5509ddd809b4d82e634131a7b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h699cfac6d81099c0c3c2006d1a9337c9795be8d8b5713f65a2a56814d6450dac3fdf73d88d276f21b935d24e90ac16addb2eaf019c0a22acc9219e993d1af1cd403a202ab3195116e7f4f2f4f4075e873be949411070541c0a58017918cf8f6e2769347f941a3aaadbc7edfccaf87fe15c5f4248033b1afe;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h406b8e8d22fe9164f9b743f9a70eceefe652f9f6b32ae3ffcf7f95fc5ec2d6643f7368bcdf84a6c811a375262db75e0b918067411f424d0ccc732bf86d5f6e4e9c526fe46d711b8f3d1d12e5f15b9f1cc943b3d3f2a1be9e5f7d3bd57a08a79b35c67ef756b59c59b4f9189601a07b589d6cde6c71ddab66;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19644cd63919ee37003b934a435edda2f4b92f146efbd94d029fde834a0c864810eb1ab6465dc4d29c6d8568ff7c92378177d0e27734abffff97522c1c1ece2414d5241af61a3592017478315eefc5746e0a45f2eaaf47c7218907f55ca5aa6c4876514bd9b9cf9babd2ac2bf7a573615cc633453c1543538;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd06660974f37939680a1066071b3b9f5582c60b2eec6f8ae9331c412d442ca81f26a34c3c44d244e95dbc49ae312e2e15bd8562791d9892eacf3bd5ee5714d2805287940e4ec225aa58299c32f367ad2a43756da5d5caf02d89f953b2f65c4ccee5a79cde4ea6433aef04a7fa86df53efdd451e8bd179297;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2ecc69aebec2319614f2abaaf340a87605bf1161c9e2e3605e7b2f6d26a0b85e1954163b71d7376791bb20b7e0ef51a2d88209440e4a17d8d00056a1e2861ce85b5fcea36a477a3914e4e3af494ae85461546694e8e5b00fa30b17bab45ec56aa390703f7eb07664ea60a9d6a897616cbcebc90bf2b899d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2f8e0d8b703701d065b4e1ea6102ac748f735fe6a41ffaa7a8ecf2fd0baa1c218760bd0ce14495463ebeabdc668a6cd0f1f6395c2487db80844fd9184d50335389d30f338fe663c801514873545a2db49c342f3dc26e161135591a9f157d262863b3f2b4365a0324a58760c8c194b7240f9786446ca4c15;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1272c431176c35c854a0080fd52f1d2e580065f722d69ffda2555b845a0a90b29ad319f115719399f79ea3a29c6c287711ade50bc46c4f7a22479030329752e0c2fd097bbe54141b28b9e8b8ac0b05735704d0b5336a06480dc6f2a2777edce468a6e096f7676da4d39e42409b795fc81385fb3327f038681;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48178d1f127020fcdc2a5cbf6c8136bcd8104bbdca6bd6a207c8c3ad60f047b3231e730cc01dd1a86ce6f197fc6827262c1084b2bfe7ecc9ef79d345b9f34654a3745072c08bef917ed6824de4af897123ffc07500e8e502ec79c0fb2de14d935349c879d4f14af9fb472915a1b3008ee9c6c9466a7ce7a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127eec096042cfc07e67c70be3c44c10e88b7c25135130654804c435e3ac8ef0c7c0b8b0a51d1451e2ac4187e60b42854b0a0560cda9dcf232393e8bb8d0aade10f257c2801555b1db9211cb5672acb3b782845610e6e79059dd30ed903d8d532c1564169f5b8729fd4ab9aa39db76fce7f1908a8427593ff;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcdaa5e832ad735fb11479a34570647051321b677ce4023dc9c580615436b8cd0c00c3c1badb2b963b2d3625a53a7f9b6e38fe55b1b0486d171a1b3d63ae597deb265f810593ec0b008b8d38f5a468ada4218f492178db549e4296c8c01d51a86cee38806cafe7c256420adc76a758585d91f9465ec582a9f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181739b14532a1eba930258672460e2e87f13eb581b95be3b51d1f995ca174c664e2719266e11527866913ad112e934e3329a5f6d27af339950dc39e092d06ed0460ab0bdd93ebebb2e6dc53962f1657a41e54fb9d2cbe5eae8fde5b641ad00bc7dad88f1ff5698a5d07f19fd80cf51481da1869a244e6fcd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h935e6e5e137945949a0c3b8c3921cf45fb59ded8dbf4b48484cd6723e1f08226a187ac5ac408732e728b3ea8b2083546b90876fe4078a58c3643fb0d714f212a6591230ca3d0c75db7f30168963a0564f2128127717e94a7278e89a5e059dee6bdd9b8afbc1f9458f788448326650651fbf1456f44aa9129;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h218fd1852011c70912d0979266c72aa24d4d877a46eb8e7e2558b1817f95a7cba39a68c35772b177a99a2a3965c338dad7ef1be37cc29968574c60a80a4948ab5067fbeee1fcddd0fc6e8899b3b21e0401820b3ca84d51e4874aa66d81db08fc6104eea3a9c6a86dc0e1ba8cb95e3b54de0038ebf2d5993b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd127f81208362223e1d068449c7d9ef2ab5b5b156286e8f27d1fa21720409adac07f903a6c1c5ca017a4cf75b69b18a9a00b91c894c3c0cc91e9424830efcac07d7beebfbf62315ea7203239874e471f13804f67c9ee9f06182ebc6e005e281c91f51ee0c3e7915d4a0da03c74114f1f63f207cdbede6879;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c093b7fa126743146afdc0557fc9d2ce94c7dd54a53488507a680bfdaecc777e17d8a77e12f763202d27d670b75efe329297f927e7b1f30123e304524d48dfe4859d93ab2a0bdda63efdf44b0621d9884c6578028d62f35b9de79a96fcca387b3800b6cb739818b3a80fccc300042c805b7992f6b5f2915;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171dea8f1162a2b522c8e57d0b032893821f4c568ea73e2c07da2daee9cb4417253d97c309d75e6d60ed83cb9c570bf5ce9b4c85800080f3e0b2235a87216f74be649c8f52e1e3b2dfdfff8cf0440159d9a8b6eceb01597e4a5f301cea326b3cbdcab076153141890357f0912b700f977900591bc2e9e1d4b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1275664de87dc37dc29e8d29b139fc1db66adc0261cf37246573d6778d69082a83305f6da59d187bc9a5e5ee644790fbc9a149c140c3e520e68992f5555629f9af0c5683025c609e494f9941975dcc3230a3fd7cdf094585c18d329d8dd49516a2e2ce93b4648b684712c929fdc2e77031b22b755727fb900;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1301113169c41e8b6d87b76458e693c77b03c78872178d9322f569957adc9287b3328f507b7bb8be6c56b425c61a87191edaf9d3a436e61ba54846abf64460db3624f7d99bc811916b0601ff2f1157a6f4a9cf2e03427d6202fcca9f96d931c919cac8f620acf3c22a31c84a1fa2723fd59ea0bfbd52ddf7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161ff3b88b7ad0ebf34e08012c832bc0c930a88008c462b3e8e0e0744b974a985705db8c3f14ab896b9e740f5e4d0430c3e4998bcf0f4657a8112beee0b65033d0c00b224d407d18c821cb9f5f3cbb26081a28c27021c361b45faedc5723b67df8e3f7430d87bd4bde9c19c4fe241d19cfa7f2d5d013348ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2a58b55d82f2763e1c88808cf16cb09bca6bcacd22c2764b29483e704d38b0c43c738d793becbe524fd9a699dad60a094ed9c5187cd6373c531ceedd14ff1a4e631781b58a134789284451af9fe10807109394e50a4679ef3c2064578dbc8591edd94095764e4e5a03fe31019184dceb014ed1bd8b44dd4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e92e689040ce2e98e1400a6c378dd3af4df7b1d4e8be37c67df39caadbe6874621d70f3340d96e986a25c7b30d20722969df34efb1a12f4e5d8d4775bccb3a5113e37aef5049c8c7e7ec6d7ba38ad3fb80c986fee554778a74ab8953541515ab523074171454ab1ca42cf181bae66bc49296bd2f34d2f35;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1080d633d044ae9a483069ce7783b84caf108857a2ceffe3a2b565d091cf9c644ef244ab91cb2d52b7a99953ec0336b8de3ed9548720b145394f7ed5a5c4c9b66b63e1a5bcbddc8d58b8ac47459862c96e7de5dfd7899a513a0e731dfe0f1b2aafdb4252bceb559872e8f115523acf1a594a1e0fd0dbbd92f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9441a9dc51e785312d6b4b1ea74abd5867b135eb155f900a62442c4a5d099e1c25162ffeac9e84cbed9581beb1bd1c682b0234126d964c79a9bd5c4d5e1f69635ba103b872513f63268b9845f9242820e87ef43c74ed436014301532b0c6127d15e7ece2a505121d3b2fe1dbf660dad11d6729ffc1cf73d2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9d8ec3b9c0054d901afe5f6d9f1aed525b9fee99f285b5156c69eb40232747065a7b2b995a32a98b10407a480d26fe9feb60e428a2bf4c01af2fcf6c540d6e3fe93b806a349f2a41ff0a551e708119b38c4dbf8b0201be5f9f9ec54c541f3403799d52e48ba9c253d495efb0f9b5969b1eddd809c642c53;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b07552d04b164a4403ec253e6758243c1c7b4c6494ca373cceaa65e4242c9bb7c383a5c876b722dd33bc16b3ecad0c697ed70474136311c73ac73fd3546ae4131d9300d612bc232342be7b1cf4f17be999f3bbcd13fe91b68bc55a13e16e81826e7bf089bd8027cafa3216080ac89056ad40eb4737a34649;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151c95bf07fd6173dfe0ad3074f7db33f63889a592a67b79030fc3365c6302ffc19d90c93117ba050726ea23c6cfd6a72fda929421030323dd02d855ef43b8e1f91f8cbd997ee9e049cc71633af12c171cafb5aa0c23db3c497095b86d5b0a4b2bb5a23a9c3e09f37648e3831ea766c5425014ab3cfa4c498;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9b5012b22899b72e58c5a0aee846e84ef95efd9a42c76ce6041a2db96f661354dff8536c257212cf7ce19ec243fda726fe7570b3e2d0833ed08fa47017478ef56b11801cce45e28cd22f0a323c5faf99576f7a6171891bb82f67544a34538ad6058105b4712ce10159f8b356299e86f16b63326f5be9294;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b5c605018a4169ca860f439cebbb4c25b7d96472291670dc8a1f7f15590b64df0775c50ffd366e893eecc74acd4e5881b6e7dacb327567851b26e4d5f64953ba50cbc539eeb9e93e1f94536b934e7834179dc2122731b123dd64830e9fb7840ee5c6f794211a7294d426a2e3adda91dc72a4bf88e755359;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6a6dc2c12f275e49aba817928ba9e715e8d006298ff63b4752817aec3c4715ba38cbc1f731669c6c2d3d9be508e759da6de2e9d6de62a81a41a4db315812e186dd8b7f33f5fe202eb5ec114633fce73400c19ab604def8ae3a8f861477b4e5a72b8659567588cc40e405adee4961258a6a084bb4975e790;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6128bdcf77bf6cff4a2c2c6e5f5e577c57905f63be2b4f30844520f6abe3c4ec3acf3f66ab8370569a030f66650057cc7e710e7e18530431d913b341a272805566929b05daa942809ea46259c2bdb627c10b8a3570bc1b5a271d03453392d1ab6ff30d50949a1ad3e730827b86d0b2edc81085ea218a661;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h419b922c525f6de9eb74fe4438f6af6829c63436550b883d06d8ba5007f8a4338ae1337a3943ec77c7279338e9f59a625472d42be827a69f0d8e4effef951d7b43578f96f09f01158c8517b707207493644a9cae3c2ba28a469b66b34963c7e0f11d58567169be61b8c6899301e051121d6f180ae9b1488e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h30bf6f3c152a368ad99cd971f2e851401a5fd6b60364eaa0298b4c087ed12898dbf82da86776c3e48c34e29f5a432e847cb2abffc6b649c83377982b216a1501d77792bbef5719ed235e6abb4dc49041e4427c02489288c73e0b78f27b6bf526b712d366cd48c2be51e92ef60d1bfe62a934ab4bd8bb1b8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169924052b46db59843edca1f53621f87dc8ee28195e88c960e9ab9d2931104767c402ff232fe07a33868e8fdb279ce7f643dc140c3d155603f48d166966e1cd9909a1e0b8fe98a1f53e7830e266aadef0e5fe047523473b99a2ab4a2f50607b947c8b86ba3bf8825fa52f47bd801d2fbd4b9f2737e2742fd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe9575cd69d8ce2388f53acccde01ef9922a6d06e8bc74b670cc5363f7819d13fb43acb10eaf9a248e8eff626be29bbeb8ff0b9428d180fa657a493ad18448f4e81373635c4c10fcf8458be7222241ec14b426109ae46cf0ee888dda50e7dc32bc85af3c62b5d1a88794ec64a0723e373df1b04e93ae32b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7621d893924d4ab5bbb409a130cbbc9b5208269cef6abf0ebb3b62c928edd79a22a143b0519b70697a0eb84af851badf7deec1b976a39551b548d3351b36280b3eb7fab87b0538178aaaad85ec5c75af6b3d4b4ce4bbbf1cd4ece61bc9ae3e23e3d92f0a8f681db574ea8946f51282404b23c1d3bbe34d26;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f05b5ab9ce385ce44e18d3e53fcb575e3d0c81312e7b493348baaa1719a6e374ce4741f4892b31575991ed331c7d859d4e0db8a1b6a8d5e03daaaa9460272cfe12e9c5270687cdcf240e1e531d742a92313ad82733f05ff2e90ff6d6c29df896edde4962618a433451dabb2adf79a8760f59a8c57b1b862;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefb14d8b798c448578e70cde8b7e9463b6f0358da6c8f710d0cff25c11d7b79f44702cfc7f12c8fcc0f377fd465464c67ad9b43b6d008449d3b5175a23c8ecd60811dc92b54657ae095cd7a065226f9577801b4385c02f48f793e6425792723cabeabd6a77f362a6c7caf472531f5988fd4ab6b4eeba0556;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2283df6a222511ccb06678e29355f02a119dac24462719d8ed053b0fd3b4454ca5c19f1a6af66cc6e544764deeade37fcb86a2b028e11fc64ee41871610c92a2d97d2fcd5a716414b37d480723cf80f9fb19238172650d798c0ccbbd703a0a6f79231515d9441166f6095dfc1417f60d248a61f82253f10;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5e9683e2ad5b0b9fa782a7363425a0add46f5fe8e2a94dba4f79127b6646a9e6dd9392b00bad7316858a3ac2f742f85265e01c1ad9dea5c6702c9ad8b48cadc444e79b26918bdce6932ed05b076d69ef91bf54536017bc1037e9408d00776f98f169a596a7a7856a55f9493dad4a9c6fb0b2dcd870ebb5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcaa1e7f69449652e4e5288032b2b20315c0e84ca4075f5461be5dd08d609c5de1140a865edd95206dc5cc713443afeed9d361cc5dc7ade9a4f41dbb5b583105acf220d0e529dec083105aace1dcd58c4875d49f9723b77fe1297e99814035aa87a6c898350e56fd0cf9734fd7e4fa62cc5e752f1e04f6e0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a408d2f69ee1905b581d5a9605875686113a7deaf34fb0b55974d0a9702e74fc0887a4af09b758c5908a53964146e2a85a647d79a188f882530bd5cc228a50026811b9b118c8e4e06cd30f58a34bee6e2704a9f287dd07279ed4cad9cbd68ac5e1575b8ca4c45e5273fc2bef2250c92da07fb3b8814219b8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13681a86b302e78d6073278ba7a5b87e7fd99ba79c5ba5d109ac1ff45bf6d91ebcf459e906c6b766fd991cd45a42e609ec52c188517732636d83a4662f9f366eacea4b05b5001772c5dc031630345c754ed9dc449394eb5efef3864940bf29d3f6a5019d44f6fcedecfe38f15658d9c51d4fdefd6d2159a4f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fe7169aaa75f8ae51401161c0b6a02fe1448ec2145db5cbb27800e43d48dcfdc6f2492842b8a580d50ebc538b0b1377dec6bf899a6d376c5fa30d56d523485597b522e88cfba3f6c1791fed69686eecdff020ff6f79c29f11484ad72ad3e10f2874762d5ca225ef2f7040000a42a47b8ba07cbf11c8cbe0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4a880d90d604ea6672b7fbb30504c0785a2b403bfc2fdc06eed32c03ec2eaea2abf00363fbc01d05eeeec12f8d1e2db8bc0f8be8789294523516dcf7767a3479e632f2c078c85945e3a1ea646437d2ef2de03a7dd2c078f4e769e1ea29ba2d79c265c123644343482be75a1a9561daf5b0ec17835ebd3b3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc137e479d7b5b049b746cd3c5f1ac38b6b71a66ed68b3d4f8bd9ce828e3ba80d62b2e83c3cadfa6fa8a5d6a8caae3f0e35b4faa0670d5a1bf1c8532f6af0c1a408658d48f395012e08a25a7a962b06665c2f30775faa0953b22513481542f577c2284d3ef3ed8919583aa629f7dc26f92cc6eddd054388f5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149f56d84a76ec281c6674cf686a74662deed69d1943e1e662487a6610fb9902ca29e27c8adf836419a294e0dc3a45d56fffce9a1be56dd38e355a1e8d140dcc50881ca1e1cf62f0f58ff56a66bae63292c59d472d3ab50b23e847f41ddc6f4ad2743e4c0ced41762f7fa8981c692ccd72b9a297f2df6b85d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116a8bcff5425904631c28194bae0ac4e0f7dc1406697cbe2e5dfd7e3041a4d5467b5010320c1f2168f41c55844f47dda3d17d4eeac6f63a586215c5b703ae87a16a309533f2a2a022c26408f4190b5d28a25263fd55ad20466b2a3a20f246fcc8a7c1f93327891d01231dfb57d1f1e9a0d0e4d721ee6e6b1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1776f1c02066a531d5efe4bdfa8a0358e16ddbb07773ac4d556c8889b3fe5c1f99fcdd129eb28b61ae84fcf5b652a08de6a14e8dca184065369d50067728392a0b25db401227540a8af2ffbb1c13f6584eb4c03f0f1bb7e168b3f85a2f84c13b4926622c262eb90ceacc8e169234aecb6a23fb28856b67a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he545500f890375c7d6a818ce700850be62128ddc0b2ebe136e6fdb7c8ad22f92732e89b92bcb9764aa4055c23ee6d26782acbee3c497f2c2427cda60d800763f53725013c09b8179c9e1a7fa79e6b98dd2b2d2913975f727b6eec3ad7faf7cd1eb63d50024c48567ba35757be9bd24097427e4926b988ab1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf035c85364708717f642f01fd33e73d70674e4fb72a5a4a83833505dd2c931b02befeb462b8e80799e73aab9f6828ccc9ef9dec56cd2c92cd08eb5fede7e14371d81a4da0e28187b83aee30be0f52ec13dc7c0dad9f0f93df1b2096570254329d6d12743b26a898a6d1422ff4d7950bb86f4018cf3493f3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2c056739329976877e514af1bfc368d8b6d24097366fc300c512c477069a0907e7a3a5161bad83547277fdaae3c338629ca5b3e7efee2a67bb8520586453e37d402cf49364217b8104efd5d8bca7254d948037231ae20d64326c13d1c2091115e2084af2d20b0641a3a66cca18f52cd79e8f4c716ecbf5d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163ebad7be83329d54d82605148c4bdf285138e1b636d550ee1bc0b5e35ddf90570f388f952bb5efea42120d2b99aec856968aa9d0d22db4d0a022d2ee64b3734c98905d8be7acb5bfe8af3bef3d190f233be314b31578de2454470e420a55dde75d510cfcdd3566ff523008b7a8c3536a1f6fbd966c1e4b0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27eb70993e467281c77260bd20b280b7ca9839a304e8a8a95afd0e37b508112d340d79fe2bea12f23b959f6ad61b3044489a59f4779bb4244e7cde268f9ab27eecfd276f47fdda9f33c887667c691140607e245cee513658114e737dbbc573f9a18d2af9b7a72f5f16b01fd911cd98ae509e283818385a84;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d7cb84806d4abcfd60d7512821ff79052aff8973332ab5fb2ee4223943a3a3252da161a3de59295c5c5de00ee63a3cd5eb772bcbe1edb17a7c0d2e14fa1ff406d0b0b021f5171d920d654473e2a5845cd334c2612f59164aff1ffca8649f66814d66deecf07381b4178c8530dac708b32c0abedc1ce632;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168929dd13debea096019e0becff100c3c4424ef625018ee7a6e6b5a1daadf92751e942bd8b12a464128339a1932332d8d4027d39643e2a5981e236aeeec3b34bf1103c38f61ed8aca4122cf5b36ecb3238b9d0197af337a5c98f23b0ab968729555969230f8f4f47164468eaef2fdf06b66b53d22e0e8879;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc89eb6583419cbc82fc0237f2c2cdf5ac7bcc8a5d18f49b230fdaf1be17d13f442e5946ece2b160e86347f2719e1d80be4ea1da5dd0e1b08eca1adcfc3a5e55c7d2d8e9e35462e8422b4f778831efede2975c198017ebd6c83e43c615715c911bda2f57f8e0c679c97baf3bc957d07a0c6fb22d652affef5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc517956101dc4039f0519c58c7ac87d16c2b1ac095adc6fa8aef55e260fa98b4317a2fb0326832548f435dbf7c04304834d8f2447c49bc5f3fc843f09ce992a57d10a84ab3991edb64b21d8a21adad609b0d00b1ebab64fe6c1bfbfb0f3cbd25af8a10d5fc775540831a7ca6592a13d8a0343e834a07c2e7;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e81d1c80c2c060f8d09a38d352d202d3283b1ea4d6ee09ce642d43610bd048acf6ff8f188406f087cb0ad03d741859a9b12ff901626c9f43c9d38fe0301df02982b791fe03d76fc7b2abcbcf116deb34e20fb6684d25e8f87e666da95db3513e28e99c95fbfe4a1abe96f74b2d3970215208151ddd1f970;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13072417ee04c7d21500fff1d464519cb91dfe0eb7998722a48db6d2cb806ac87946b1cad55baab10f341e3c8a8dec335b327000e346508a5f19ba6344fe83fabe1cd0e2430741a756850e0c60fe88f2e50c5672449780a48d830cb88cf01c86c30de1ae5ad88cd3b01205a8d496276dc0b502c77b7999122;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0f19a719bfa6f5970d229d11ef1660626c93d91eec176b0be0671a0c2dab9783c7ec7cd392700459a16903f3ca5b82e3ac57fd5125c5e68b12052e564e4af003a0a8e5e527dd9e459fe528bd9a6c25d3f123b396f8ae69e4109c30b3ae5951e8adb8a1357f9a8665534580aecb2bd319aa70bad823c8fbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6e79888cb18984592041f17b513b3736fca91a5b0f2d810ce68f09dd4e8b919f2bc1e845ccfbe0cb04a30f0afbed6aefd9d44eb43e54fa76c404daeac148a1e82c58804e1cfdd2e54c8db8cce67edefbd227cc806d24056dd214791a54974f58f84f3aeb972a8b6e97c0b6012c60c2e4b5296d9c6191971;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb98ffc9349d26ddefd24188bd6e8d5a7a2b0812ee8950ba5a378c79952d28bc8834d0707c871a804b5a8286da4ba6cdf804a2cad1ca9e5abe7edc45c28608b671ae6c7bd78ffb74c5e0acfea0dbd200efa90e37c674e8c515326af9607e0c6d3fb3570cf06ecd0227ec373ab08788dfc3a37c4d2dfc375a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e688210a022a952ab3a5620a64a96cc08a6748a6e52a8aa0f05553ff96f4cf3d57af625d72b22e462a4f5c15276967cd8d8ff474021af9ae3c179a0d7f0473b3102c640edc4402e2e9110fa1b83ddf3c3770219267360b44af638bcaf1b9184aa7872921209421aa94f6c360f54491f87af572ad780df6b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6bb734b55f831435e04ecf6908934d17f75e7b6eaf6e36e57842b24f4ae0e9094e3eec42329f4a26ec06366a78eea747aae155f8b60a441f3ab5b537954fd754284a31ba1816ca623d700745d1f645ce9ad81be8ba11704d8e7bec8de5dcc8a28c91349edc38801720ebd1bcaaf7d6197367fc12aa2bd51;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9bf86d819cccff5e9e57e991e016a8b7dbe500829150ed38e51d6a5c183ab0ed8bd08bae3175f112303fff695a6471fa068f3b3cf0a87b8a21cab92ae34d40a3ed456d62580c9125978fdeadb381e929aa646fd4b575d17ee99fa615ff5481efa2d19b50ab3106132fd8dd5eb2f17d9d96f389cc584d779d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9efbedf5af50ac87aac68bf87ada6e224bc0404adbf074febad36d6d870fb66d356d86e7fa7bca9ff2b247352950482c4633dc8a6975ccbd9851cab4a4dd9508bcec863ee19776be60a9709cffc8ef0e7c7e9b0eb158de8a9c708b5bd42a0f2342f05b6ca2b97b46dbfc76929b9962e3dc25841c29cf662;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bcb41bbc71d8ff258ac623e1e72f6f387f101c4128c82e16a6d7ee34785e7259de4bbe2ae811810ba577851864e229639ed6cb8fb78a4437596923a17b364e761fe685671a359176385e7c9cd505c73e323a22c7714b29abad5dd5026650171f05806b630cc6113ffa90bdee36607ffbb14a084efe95306;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hada81090cd983e895b11a8318208ca8bc357f10c629d9d3bed6e50d3fc9c5f1521c088e4c65061a7d2748cfaa673cffa7a5372948648c5351210fab55b5abaa8dc82e9e56d981e13bdedb184477c48b64aa6582f912859466c87ad396b3008d02899099775b7fa9764292fbb2a24dbe8793cd652029fe205;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5d27bad849f4bd144dd480109e9b79e396f81c4e7cb3edd548b9891b400245af74799b21482985987c894ad52e7f18e97339f96e4db7a0ecc36617a1cee90fa17a0a5270abcf1a2bd48a5ff1764c7e004234a0455f0a952fcc575d78786e2ce218c3c9ee3ba28c9a38e769ce54df41179441d66e06c1474;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12721d84e231acc70eb318f35072cea681de0a7bebba7229692dacf2df5f89f54957e59edad16a96dfaf2eddeab9cb931e9f2501618c38ccae03bdd2db9e99e6d2df65dc47b2a8db275c7f214d40032f652f8faa547354d64d8b62959c42b84345b5fce068f25fde71d77c16661a6b4c49ec031a1a8dd125;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b662c266284864c6533d98b031222d33b00b37cb3e4f6e22b7779f53851a61642d677853b84a89f00440c9ca7df5a7d54395b14c28a13fa00c19339bbcd4ad42a1e559a4a7c87e0952723818b07aaf4a395bf6121fc448074d5614bb7c8af5282b8eaf64e8a2556f221c999d8746d5cb553e892285779bc;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h911d6985a264cfc8a96f28360d683a6212ef121cfb979ce7081ed1122fd165ec62d4848bc1bd6c63eb03edd01f382b16d19e69e17b47dccfa91c01c0ad7c067775514caf956d67bbe403080df8bf7159e702b6b3504b1b52ccce60fc07cd5b4b169175137dab2b182e117c6b132951c295c62ad221910838;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ea86fdcba8fa59b2b5a0cb59200f455606d803bb33612fb9b3cbd34862c11dd9584ae78109f9fb49568eeaf398042c7e01f703b3f09ac99943aff41d7c68a19284d9aebe6eb84dec7e8183707347998b3c7a33ae3a1fa41160473bb570143d67fe890a8a592dca011b9e15abc62381a848648ac474c687c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h325638b5380e7c491e08d31fde443eaeba9db188671c4e26603908d58e6193aa8f1bc1f6b457df750986b34a8e068b8a4a3ac1cd3282382d717b5a4d85d1cd0b28e7963c5485517177fd600b4ef4be7d51f244c704b393be1370d749c43058e2411d8b0f767ea0052abd48ae50cb36bc292151f71e4cc066;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17472bc81a8346880755c0b88cd8e5a2369520bee1d0150f56f22cb9324c15f05328749366ba732be80904c602df3a1d913bae200a03bf6b753390e066af3ac024a0b8f632f6286b0b6ea458674cbbd0c70c9ce52b82528e2f806e2da49bfe2faa47cc6922fec098afa940c650107383a1dfc6c8461420870;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122e1bcb9a5e011d85a453e7da96d413a00dd5fb6dead8d3464772a896d128fc8d2781cd64db0e8f7b374212fe0c9ed5496f0f88cd4ca59f034d7815e3f4f1565d13856bb43b181fbbcbf2c507e9bc4adf5d3514f94128237b638e3b639eb5c934b4147c8001353933ac6f7343b8b405bd2a79496f2ee1c6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1528ea6f14fd0a20ff797a715bbbed370ab027dbc96d4a92efa533f1580ababe9ef402e335ff77ea953b777e9be3868a78df79dab12926aeb9f28064b198b25e9222191a788ec45f2b31b3bbee83bb0160a611b9041e3ff47e106a4f73d1d0b29739c8ff8335fcce2803d0d3e45d290c168cf5bbba27ffbb9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a629b6f836ebc7a5eb0ee84183fe224a428a48fe450a01fb95c35d131f2023638833f4319094ae76bf30822c9a7348ba9c63ea2f2ecb63ba47f9135dcd93c23552ad6f956d2fa61be7a9361cbe495cdb2bc651d3b636fddb2e7caa61fc4d01a7ca644cee00b03a5b011f69d16b8a5b2c228a41f7d6893bf;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e75e898bee65dac7081c82e5bb3761356f2742f14e6db5697f0ca3571607dbb383433de6fbe5e7d16e490327d187949c9bfef0667a47672b3e969edbc019ef41ddc9fe69f8c1e8ccb5dc54a7cca08126e1bf64fbc3a203e8971352602735de61273c323f6554cacc4eb143dc1819de30db7af1a27dada623;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a6b05d8760eeb3920d478061a50e70697e8db64804379edb33a482ae0b4e1034fbfe859c749d1abb71ca834faa6061b092768c90cca385e2ed7b02be3fde58014d9991e59b0d9178774da82080c4b323ca5e5d3503eedb7988e0e5df0307f8988e1eebe532ccaaa950c7e3a42d2360a4b99a27920aa1840;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1350fcb04be187959818aa01cfd6913763c79ab65faa219ccbf42cbadd1f25aec163375086e3d67e1809c15bf2b19d713db12487017a67f18906338fef3741dee9c141c51ec2b5321a771860bf50d4aebe216b0eb6597f262f3d784f1eaad9f52683927884f0591d85c6388365cea55252ee667608e48614e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad0cb08bb452ff32b9aedc1aa644df54a13124bd7353792d29d01d4b45390e21c930203aa535dbbb69f05485f3ae32bc8d0f7b428e2d57c2b60ebff1d95f39002372d5625d3290de2ca4d4ccd394366f51ef29741ca1f704425bd8beefb52f1e0fc9337c45d36230b811320e7f49db0abc5bf19bd195aa2c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa6ee3f9a341da94b2864a46957796c5ea4f4b70acdc6416fe4814e7f9d01e12ea869be6539bc673804ec557bb674efa5c78e83b6b57d6f3b072b5ae05efd07059ddf54eed1d907818f05107f2455ef3fbd9aa40c2d64502abadd92a8e55fdb48d74957ed9a80780c8408d50b0ee790cb8714bd4c47a4560;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77807a1856f7d4d49f47f3b0f34c5bc182ea90e5c30c6213acf0a726f325d17b7fe99ad7155e49219573dfda8ba4e6354070c13cbc69dfaa53d45e37d9b48a99281d064421c80d212ceb39f1879a2e23ac1153cf68f556e0bb5e6736793c51b5a878626c96269de1bc799dea2b5ac9b02d11ebd30fd5ee8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd10836d17322c11454b8bdcc41eaffb572f486e0b86e5dd0b136bf395755e8cc7bfab88efe7e7fe653abc5776a38ed5c8035e4fb3645bb81a520a729a9ec3c86648a9c07dc98448ef0096226261e2cc7505c36785f51cc9fdef7ff38b0d83df8a4026eaec638088c8a733e0e63fb70c2b969b688de1036;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e35a201844b3ec3b78f791f54476a7116d9695d515d07ddd3dddd41189a38cd09a663d358fa22517dca3c32f2487d8ea27d21dae7263d2c38c4fafec9dfdd5c9c3bf38a975e369d828e334f7670e61fde45ce610659698e5238e790540f4fa1930ec255595e28bedb6326cb8899a2e297734813d4b5451e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40d9b0c6251e0ed53676e9871faad8018654e9fb125215f3f4547d5db967f694b4495f711585567f06dc0ffc1c35feef39258a6a921d0e7ca7006a0d84e269e42c4adb6a1cb3f747d0c32a4a3867f8c44917cc31c7e3a6de6b0351abbc780df3878395e73c2a3e70ba79fc9663269fc358b92b6a5f1f1f8d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b7daa893f00a021b9a56d9efd2a74d1b10c1e8df2f09f9cc6e197c293bb9c21c2824daf1456eccc29b707ec3d0c05e192d6abf2449dd66639d17437ada197aab5523bda88e62a039d53ded833fda1ce7194b13405bef52ece5a150e8a8e191ca3f1f5dc71bfe799fab17cb16496d926cb3f4bdbc9536c9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa9f615f99fdbd89e6a2b2ce4f1f3c19f90bc559f9ba7226a72b23758da9fae194694be6256c8fcbbe53d1099cc0941c4981afeae85175716f0a2462ff40092712a822fca521ce49c497a34fa91ae36e86cac428031b938bf48fc148f06d96c5f6ca5d3b18783e3cf77c8e2b7ec95f50676b209b99d77960;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32420d13a230a99e8c218ee624c19f6453f8eb481e7ab7c06621fc1d89c708744657346ede20d0b993f3576280b3c813498d3341860d345c6cc6cfa968034578af8d508cee902e5ce87ead2c214ad0ab96ef1a8401be7ea9550da3dac236cf935a3f6a825e49ea3cab1582bd9935e8193f49b153d5a57e9e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9e75596c4ea5261ec7bb5a64d45f660e536dfa8eb6d16fad3a10fa3d854bde70884c621525b40209912fb10523f5c2ea3fd22c5a75cf4ca51fe04f6b2b1ad799d9dfe70d8506d8b6f6342f7a95c48efdcef154947e2b45a1941d6622553073fe388132a6d8602d3829c32eed472adad05abdc3e0714392a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4fb9ab9a475e58731d612cf24b19e64b336b3faaecf974587121db645b217ec82b8a605c7e704bf3a4f3f74c2935292c914f16bbeba909f1e720bc4d71643e2be9c8157de975774bcb0b03aefd99a1c4e6150f5162fc403ad405a748a747b08278a8bb5f8cb6969948b9699e40d3cbe5ab12818e1da1cbb;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157273e072cd2e29dc405fabb36ea83d7f0707e9738b1e513e9a5d3d6181d8f8a80b172b3464241b26c380ac58be4749015fe7d837a0483c44e8547e5333b78a45b5f2acf012eae1bff4a318d60b846ac60edb04f52f633769413d1dca803e13855cc56984f72b325f32a6a0b854cda94c4aad5d61d4f485b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29f6b49b59048ab13c0593da7c06b696046dd00334844da36a6c649cb8aee2ecfad01596bfce7d1b2fa04089b24da1cc70a7d8646aa0c3dd509215685ac5f32b1864a902a5d425d470ee2ff993ffdbdb5792c26082dcfb45ff8880b72513d7f06cd4b940fd9cc7e2b877c8060d9eaf06b3e17b5aed247424;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1940282cbfe07501dc52f7809a01e06bbbb848d175cdfa63b7c61e4f54dfe9575018b89a934b015ed98429cf837374ac0955550735a294181fffd1191b14b1b433b98434a63f34f8f2203fcade46781b78ce0875bfb7a6c7061274f313cfdb59c1e952219c5610732831f127e58f3e1f638c846f3807a0050;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7de191f70bb1a1bed84af5e3a9d3e217e74c8909c73ab95ab28d2f0a845da94f073b67afdd5085eddf206311554924a9675e1e5dd124902fb9736ae119b109f8292c21753692fd97b41cbda31e40165fba1c21a7e5fd5e3e69d310ff3c83603c4cdcd19321d606e521a11b143f959ce5cce5d89c28712c16;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he06910f45aed7e37367c06f3c7d75021c65b8c7cab73d46d849ebb3ad5ced54a10bc0acbdb19cd18c7acbb6ae1a9a4fdab11891c68c4f324b4e3f28829191283f62beee33bf2562fa5adc584431dac56b6031f6da5812890c82df40bfbf9471b8005f42adccacad10df900e0400a18ae146112221a8c15a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8999b75bb0bbf707f78d1e36acf767c8d9106f69ac63fbf1e4e3c20e30a15ee889aae968218d7411c0c9243021efa8f3f339d01735c12b6908ef8905ee4bf53cb2ee819ce9a191bbb9896b5520bc166a85740471a3a2d194a2583894b81b2827032956fc089211d3cd80386671b34e141d89f860ad3aa279;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17985b766941aebc723e2fac625d81fe512809d391b96cd1b91717a6f214c54db4d36d7d4f7fe2cce0daab50d3db9d270df09dfc3eeb1d936837c3c6aca22ba6bd832e0dcad1248a2f75d285776b47739b18c62ab0f992937e051bbebaaf87597a84500af9c354f2bfdec20fe2df991a7da7c8eb05d45bb9b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d7b400c4b8f7c73322eb9af40d4f689c857e5ca8657ac685dbacdb4a6df10ccf29aa4187caaaeecfdec96b9f6c771dcf81cbe1dc3df9e892695a7cfe47bcf40128d05b33981dde26ba161ad30079cb60e42777a17c60395a13404fc54e7221852ac767a3193ab6535a1b235ce63097681002d158ba21f49;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68231d0a943241871a46748c5083dbe7ffb5e88411915e658ef568d17819a3b9016479788429b12780239addfb1356690ef226f395ebbdce91c69f8f42c1202fbc19bdf15ebf94ca9b707a743faae54ad87f659294f6077dc26b1ff30b51524d99ba895e10f1c439feab5b3bae24c459ebb43b6ba69ccc8e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6b9c3c3a78410242fe9044e4a2c694494f6d74f4cc782a86544d33eee176a58f05fbcfffe269f8964c037a72f958549e502fab031020cca1706157ea231eace9720d7138f1267f14b228065c49f7ee5a8490da1bccb3c048784cdac0383b5a3703655ab1205bb907768ff27042f8b458c05d213cff1579d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1822c0834c8bb85024c3a9016253b06b17d97efe01b58ec35a1f27977e6bbb4ab646775c0f404de08fb9aaea91d59f0ca870437941259d2f430124eb5f5d8454ef3663e002ad5c89c575597abe906a75b29d153b02071356e21052adf3cb33d96418af20ded775e33112892039526216b381bbaf8edd9998a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8ab8ddc58db437cb170c543ee2ab5ac575bc15e484aec3d9bc5d5418bcfbbc3b204fb348d54eb4fff8e7db5a053b9b594fc37e6d809f0ab4fec528a2d9490faf8348569c072e4706bf68da97c3a4d5c5c5e446e957ad670972dd22e830baec6b621e7179710682ceb6250a12d05f14426f47d8c8979ad64;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58c4ef7c09bd345fa073b4451f040147a195c56cc0ce691fa3e08d0b13406b433264396bb97ad6f8d4707a2babd1d34353e40059681f0dcaecb6aecd8c04e3841d5adfa8868f65bc474ab14d89dbe40bb10bfe8d69620f35667f18eec8644a4c4d6f28415a7aa85e7920c93cb31ca674577c9e5b16654e0b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14be4a152f92318cec79d79e540c9ab0d6eb19be617fbd1b57c6dd176c49c38117e052010acd215596024a287127a23bd7ad819f51641ce3cdc60ab8aa9f50e9cd8b1b0583a6a51c80d5a08e91102db26c4f91e9963241ea2a031c7f5c005bd93f3deb784112a3575915f9b4ad9e322b42d0ba7406f41a48a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165acfa68fec17969832b894cdb77d4c6696d5c29f44c3253f01def6bf55ab90e5744e5b470b1296f16eb464b01fa665f3719133e432255e836415d6ab63a87700422766592d6ace46f21ab780bda6c9cae54da76fcb887911ccf4093463723b9a5dc102a74f7b81bba03d838f2e9a4e2fd802c97f03e513e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12af063cf890922392cf3c25031b27e61b871ef00d4bebc0dbd5dbba8b2dab2c50b6b09f2cf2c2aa690f722b91b45c0d6e6d98b2b6b11e13faf5b58e83fb17dc56389e1fd73a6544633219ce89a5b8bc6c2d8a165528f77832479731ac5b78ad2a43849a4bc0f1add79b9c9138f109cb355aa6dc6e912975d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173a8e0291a6168e2ace9b44499e8c93191a789c1b5848fe7e945a54c793f76f4ab36ce138ade7eab2d488088e417641fcce8a34830db361752f7668add657bd290c45cd05a0b8b13138c3b81529d604345758b3fa4d8aeb11704628902fd8c4aa24e2f1f1018e886c80bf1aad3f1997fd5eac3a72a484a69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ababd40cd139cef111418b300da915ebb6c942b8b12b4fdab16aa2f1b04472298cc03b9995bddae90908bc9ba3e5be968d35026cb20c93d5ef5820d3ca8f01e3fe64e60e94de2f68c8ce000a8ac584cafcf8228991c40fe83a1b84bd0a3ae0899576be14a85ce5db81c494b0fd4d6037d6914768ed3ae22;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e5ef4b31d99601bc272dc39dfb29a5dd7187deaae9b1a6ada794961dde0caade1051ca866726723d56c0e55e95a329aa596b4d1d2fff7519cd02dd736eef9424c42c9beb6329f15262dd6b108a56c9b70d1234db704937ff624ebbe52b6926bbf17e524a543546294886809c32475ca3b8797184fa35627;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16534dd57d95cb3618d2155d76885ccf7beaa260686980fc6bf006fa8abbabac23986a2cbdb2568ef42cbf85a2cd6f9c3b951282d89889d8005f0f7d8af26731b15d4e0bee0ca680635dbea8ec3d16574b2e80479622f346711956a255cdc55b6147eed2383ec5eea2680d2dcd4af0e2e1b9a3168811c04ce;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12eafee102e1379bd4557cf9b92d9726c6edaf2d8b4d73a874a489e7edb7ebbbdcc48fdae603b865867a6443134e187cb8927f513ce867929b7cd79bf3b4548f526386eae11ccd3d6445f2988a6f1b88546a9c3ea7c43f3bcdb34683a4c803a510e10c9aa65b02fc0f027cef6fbde14a240c15398492036ba;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0f4745a13dee7556b2f354f000b20876c2bfdb302e699f4860fe0801cad409ca2335ab48066702e63616ba56c409a1040bae98f38561083704a03201a725aa67354a5e71a882bf3f04144cac27841f0df4e5ee5e0ed51e21ab283d2cc9315ec0a10b419491455362155c5d98e7ed0765622d29169dcb0cd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8c79483a37430b97ec61d660f91d9bb89a852d7a24fb6ddbf93aad6b874d062311dee9bacd5a9e5d66d5fba0bb781f62a5192d017e02cf335f7aed920e72016c6d8792989713087f6406dff8392fec0be008460d73c7e1112c40b0c589b6557a79a03e85894af1dc8d42f21f493809c2ada93fa111eb6d5;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5787006d69f09a3aaa8bb33cddb2a9b2518615f83528f3b248cfa748edd4d4a8683d1463fa866303bb857044a4af8c37c6b91ab99e1619e5d4656fddd3261384b7d35074c72eb8161fc9a8a63eb3b6f48a9d18dcb1497353c232883648845d89647abc2f6eb1502cccd27140bbf9904a3dfe81e3601fe5c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a63ba2ac632d2eef4eab4a4d8078c7d04ac2d036fc2d5c116f5cdc5a04aa8478e4f45540a1b56692151411fdaaab1243a5d6b55e74955e86432bf34772cfe57533f25a1903c36faea19dde0ce62310be8e95f98fb8360650fab4acc9d0577d600c50571024c0d8cd94ac6e46ec3137365865990cf7fb31f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dceffb810c4dd24c7c341a5d9b9ffb3be860f556a82e52cc81372d7c65516878924ad12b728e96f65bed6a1ddf91fc05b176c84b50ab1e4a395219e3fae4dfb2703117c73d0129f36ac9289047fa4342c76f32d331c9556e111e3824694dc688718b9294ee7f86caf64e70f9bd34443dad8f26d0242cad47;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1286187b90c5fad13d2a8249b6e14fb5530d17d6f9e25b0b354f6c82aa2c4980fa89a804ae87af579b5d4eedcb74e3086d73b69cfdb653d81a69b0c7df175ad592ce0bda11aebf87a9e86a4f802818416c5765391d38c5d0aab968fc02261fc44859297c8bb294e049faf02c9d73143ebaea4191de73767;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fb990283d035bc5456f3a6062e320d954b8395670fbd8ec498d1eb5c81f2ebe9cb69a9ce76c9bbe75c1bece69aa2b4183e3a1f67cd867fcb653fc0627f0b33c9835641135674303696d0df80d9b931ec7055f45db51faa02072463805dc5f3d0f234f96ca5ff94d9280531a4cbc6aa4b2dd4ff8c45aba7e;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d54ad9fe27f3011ce05004670ac4cf8fe4f9e1858a1f6a8759f9ecbaabfce569c081b4bd42c9de2add211a30284cd7394dd97e440561e74d21fe797aa7b522e57a137f5f51b09fba02b4d0d6aef3ebeda42d92852de7de94bbc0ac4f935790c700e704f7547730e4e589d508d73543e53c166aae71e66036;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5ab7afb6bca650f989d47476e5679e85dba0596e1cfa9470368552dfbdd5d239000f5112b44dde267f7fe9247dafe0afcce2e888ba9d43b9933e4f2b67c678bc8fcebb238f15c8986f3d29600a21b71cd0bf9f73c16c0a7aca31b92cad39e23d8cae15df911a84139cc8fae9befafe5485319acdb9e5378d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1308bf31c66f2192e185562234743a1d3d5e5544f2ef8eb8d8dfdff7bef2ba1ef2e2ae7a943994ffb6f70d88e51040696bf8f2708ab5061666190a3c70ec8155437e8c20e6a4eedfa2f638fa714dbeebfaab7ad4b60e16ccd13076986743e41a49bb1781d793fcfe17e27a366d43774a8db42b8c23096b3c0;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb893ea752d3866376e06ab7ce7b3b9fbccad6486786eafd5d99ba4552d13c6bfe8cbf502e6526d3597e1fa3101d8c4d30cf66c25834eba0e269676890a2a19394ed156360433435c20a9fcf8f6bc25ae1be90007aae631f807ba3e9a9dcc8f23123a960cdeab2be21bec51f1a6345a17b3c4cd857851463;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1279c3a8fea974055c0922f0eb964866abc51c2f533301d204db9efc2d3c90005e3eba3d4228ecb7fdf45583540d273cb91c36f26c39565b9a243adb570d05af1d9fe1316d4c3158edc9cf1916a7fac6644df03ddbeb6079aab5fb83ff5971ffb84d99813e894f8230a56e82a4036c9ee28f1700839ea6999;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74d7068898ed01f2f343ea9c1475c0b6805a0c036cd41cf42a96303977eda28bb6dbd9cd1ed8311da78a0f085583d947a6302c5547256ced28fa1c2b0b56c28c90c22b847c2d735ed9bbe813d8dbc34d462db894392e769e4155aa50d9b12be5a5b83c6e32667eb975362683a6265c909373192a7428554a;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa29f1ab3fbc73a3bcaef9d77a38f1a7586069f09042e4dfa61ead2c3574a938a73461f72d9362f5e2c24c37237c6bd5cc459b1b75329441f7b5a91c221d85986aac2e3fa165262fd1c9b955af369f28c8963b33f9e653e690979247f6173057d828873c6854232bdd6b9e044981c914662cd3a5b60a9f9d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e5c9710cca4d10034ce8ee5c8ef76569a8cccee10e238b5fd92866fb995b65cd7a5b70aed1250a8a06805ad2d279d19296429a1a822d7464823f2ddbb6e48248caaf97ccc4d720cbad4a8d210872eec6c507b76490029db0d24ccc2b1a60040fd6ebdfc295e99564855916fd6cc7e098215c5bcaebba7e4;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53f8afe3b860f0fce91fd4cac9867cf8d32ffed23d11fa025b1c0a023a193d50346f936bc8380aa58955269c3f2f7f3fa04e33cbfa9a54b8f995f040d5d61772411888c03d95a730c1309b871772c05ee69073c39bdc7df10ac277168bdf8468cd0a221cb723f737f952578c7cd581d5980d720693d257ac;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46df4e2f015e83c06147c11276528db2e89379d755505f45a1510ac5916435da629db3956684575dc403ee5cc498057b9cd88199ecead2c54faf92b64df5abf784be5c19a2cc4f8072d9b06750383fc7ec63070282fce9cb811993118132cef7765303e09a20acd2db3edd4e37040f7e93edcbbef223d5c1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd39e238141fbb05b074533ceeef29f7fc0d3b84359935485f610740eb1e9bb80f3b9902e83d593e3601f1f2ba15d546c039cd76efcad8686ee19aeb2712653af8a208d646d935361acf91f993fb6fd73224a99d7c0de26e34c36178261a65fe3fab50b7dfa57896181c29ade784b12b373252e1905f8823;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h765741985b471a42b302d9a392cda04d69a7a2c35d473cb6760477b800a24e03ccba51599ab4ad05906bef92d1156723757766e693ae5b4d82f4d4eb49dd13e846fd80349f1e16bcdfd34a007b53bc77af958996d6d1148c0c0e3fba0384429e05ab1a74ec8207d34c704b4959d5d7ee7b0c683e2209ea2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147e75e1f523becafe13e437747e5176fbf3e8fcd5e90cefc3201bccfb031a28f1578c7beb08e5ddc512e239a271b29af5d8b9fbe9d63283ca1d64d25bc7bdedff55c61cf32e9319ee394f87f266d8488a9f114fb8b95b0ed68e482afab7d440f41459b91879c76b67af2a68ae98f3902e1bef8228d005964;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4887715b0495020e2ff849442374fccf7bee8b2307c050f7ff2e369924f6c5428ca2702ef985215de6d822a3da4c93c7d64718eeda57f63ae5d49bae5cd1fcde1439ac02a2c9c76d2baeb0523ba89ccc2fd71a902431329d2fc3fb7544d4e534b0f8e1b5f6e8a5cd54a91e1e3632b28e010088390ddb43c;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74fc9e119d303a8ce1e443e8233ed31b61391aa5b99384670239f0ac3e73d5a0a3e57060fbc72374533a9301feedec9c3bcc36d7755bcebd51b2c85b6bd787f45595bcb2e9e503fcd38597afd051b12ba0336df06c3db8bc66a35fcc968f06daf3f1385080fd278cc0712c6b16ab079c29290a4a685dd76f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df7b298ad6019ea42c1c23ff12983bfd66ade1dedc8f77228319e493c8fc6bffef2cc83f11f5b510376c060c060e843b9636e20a67eb22beaec7c45b1d14941abe5dbd15cac30074fa9e672f36a68ed9632c3566bf67b63df411facf22743d0322acac6f40328d70812af704cc4f2ae84bbb2e711b218668;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2465ad9fdfe8f28cbd7c45f94f28e53bd5478c74c81f19edce8384ae88c02c6c18786584a17325c75c623fc3cc544f2760948e678cc9a136a0431195666c58ad0903f29c86ba0ab04facd9ccdf1a87b3be3f8e29bbd5a29bafe004389186ec505d7f249b33e7a727d534f1a824ff2e8c5aec9ff4e2f28ab2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1847151a060b9e13ca6d328ebf1b37918e88e95993e7ff276c3c13387c10d31815b42cc645c5c3440bc55c9907a49fb927822df2edf2717b1a7d42b1b0f6b97bff15d47d60301f21fb2fdc886046cbf068be7ae333361210047d5c205a45f272a661eb44c222d9c7f2633941f5330a5a3f89b290199611902;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18be1d4ef09a8777a0d31b36c1df45d93e481988146730a8e87b0dca1df6dee2307a6c542a7373c7f4fa923f24f027595e042e20e56d4d54f0c262bcb3397a91eaa58e8bfe03584ac28010bfbdada8e90f250f994de351015d213202094e3cd90ac9d448560bb901880b0d95033b8d09f70b09eb6239286d6;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1562ec18f7b097aae839a91459a784d8d662927d7b9cbab7d3b9ba5cbbd54769fd47da471887354da1140d9915cf3ad5af895367be68ffb824dc1a0a02aa03a9699d48fd236ea7dfac09e3d4f885ea3d5757716e5381f119b5339898176940e6c5efb14761a99806b2fbe51b7465be103967a3835f70736;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea1a0d7b0a45084c6b453f0445a053ef0a1e9b1f28d9318fd41b143a874c1cf45fa802cc2131d564694a7a52b05fab97e2ebcfb00b6c072a4711b6562480b1ea13f7e2a90139cd3fdbc45a2286a8c5fce0df54d08f03b5ffb7a8840b1bd6c5534c95275f744e0ab81db0661ce0c60d05af6a9fd2ffc2f4a9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca1a7bdaaa0fc4389c079295e85eeb8644bfcbdd8796aee41ac2e187212721de48e99c5dc07389840d8064439fb942b7d20b9e524a3af58fb4d6c22f15f04b75dba8feb610001d17faf89063678eac0cd69568eff146f977cf8f02ee198b9f0e14c6c5b5b4e93099684e40904ed0b30623e576f3905639b9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80ba1752bd28b9e36d9d27a8a1d25709b22eda8f591f1d9bf49c27598a0fc8243e29559b569ef4a1ed3959cf98a8386fab9d0d775225ad5683715a6625ed4cebdca7024049384fc7d4d3f23f98e59dc503a1663ef1a0ffb86dfcb39ad19e919d709e42debe9de4d98c6daa333f825e3368eef0cd57610ee9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63c4219485a40ece141284aafd4964203008bb4f2088c6df9f78e12ffba48fe7099d657d68a1869e696d34142c4ebe9d7b4e73fc5a6aedefab05d134573d736757068043ad8caa4e64811ed2031d7a1921cc1e3f9a747877909cee522782e896142506007f26bf6f9001e72fae6ea41c2f4f0eb56ecfac79;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3fb164e1071846ca5bd8da0deda4c1a5c529c6fc28818c6e4364c2d2cff5e7a46f453778e1f843bada8b1a3677791d9ac740ccc35b8d9c1e9e76fc44cdf14bc777e223525171844e686268c13f338834d7e1faee7b90892352ff4d215617cc5686b63c3d17c319a820aba821f3a92741afe52f5ff60487ca;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e65cb3de77ad87f1010a1fd487af7faf4fa7e9cc506d294f636bdcf30285cad3ab5b108218c650c103f40c8cca70ec648d330c5f94f9111e5014eedb25e333e1a3c7fc5b9db0657f98e8ad67867ab4f49ce6fea700fd33165edf3cfecc547b40fab9b3b1243b7a530dc4714467b2d90551da6faf255fb29;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20508b635aeff644b68f77399349fb9f5f5a74c5cfb0b36402f1e96821ac9c0bf18c1d28dae4311df84a81ad667cb6f2c89a9cb835ee0a1fb292519bb8d5228a794b693a58b7d521067ecdfc78f58d7780ec3fda37b8cc4bdc63df7703e8af4147d3d70e4fa836b66b6f8c3b6ff781df699ca156578902aa;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62653b31e031a5b30499270721ad1dade5e288b70693e78dfdd7e9189c7d72c793ad09d9e953503c443c54924eb5244c2180b9e60002bbd12142a9147f5871d17c9609a0722021ac98f94746bc41a86abd089be39319125e302845fbb6aa16572ddc88881fb69baf2d1149ca7d937fb482c5e73c722c0d75;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab2bb23f4e0460086267a9a12d967623f7015dddb93af7e8822b53ad25e883212cb27a1f28e78caa2a9d0beb56ec187be131e521417ba06144c313b4241a307da2605d5159f5302059718580cad3077b101124c104ba5af739c7e4b4d2d0b0a0a09b24cca969831827b1ab8e93cfa8ce2999e8828e09a941;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16afd6b00ec4a4ab0e411333eaddaa5535040e0ee5cf49127d3d7714daae7dfb7bae69c7490573557bd079b6c8ba408982494f41272dc03933bdc7f4f5a37fe13fcdfa8b729bfae99ac9c7c8fd35289637bfe005d93b8d122dfbbf8c279eb76f73f30c00062d7077416a2584775d7ea726a61ec5bcd288317;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h177bf3e106020457cdd2ef8cff5e7083cbb664b5a83066a252c6bb05d55043dcd11fa8252c745df26631c70154f8d01538b117022575e71751ea61a3e25fef699657be24e5a2a469ed39c58ed7a086b97592ecff72d9cefcbf873ef19b0d8a8ddea08d5f0be8fa93ee9f328081abc92bb3d60d4cb9ec03430;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c065f0469ed8e4b64371127285bf10913fb5ce9fc64a6b5e6382a8da51bcd01abfd81557215a6dcebf3a9212a23f3da85673a44437c42e4070e2b9618fafd3e8cf11adb5d41aedea88da6b7cb67b0691cc4c961643f06c7d5eef6e90c58f9affe042e5bd4f941867df03784295a53ab2f4ba8b641ab45bd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae67f76932528453b20c4668e5621169ceaabce7bfa6989d1410b3ff4983611ca502fa8abe1237ffa6e8027e18cdd465e184711125e4fab396e406e7d03cebb13d3f97df3b2bc16a6f76834eeb460013386a4626561d7976379b5c6e054b8fe093a6147b44fb92f14d0e20419c59e2c79664d73d6986cdf8;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ad18db3a7d55fa30c364c4893c2d263829c77a2bc81cfcb509bab7b1d28789dc972551860656c58da6f29bda669aa9df4c6e5996abfcbbf2b94f50fb65f6ea64373f1a731fb33cd567ae4b656d48ded5cffecde4f29983e947551d04b9e1be8656f261c23849ec559f97160fe51c52ef938d0abc8a8d327;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11144b5ba1abe823d09caa7417bf196b068d89bc85f17a4dc403f7d26c1c79ee37fed4ad2b5f147188ddfb0f7ad076184a55347f55ed9f08fcd4edd04c01b84cb27b7e5ddc852c091d669a4aa096a4de65aa1c1b0dadfd85c919a113b16455892c0d0945fd9ee7959422379ffbf49b0dad1da3da72a006a62;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106426b64f6891602a406b2901453faac2faf99be644807661d5f4dc5596695a56c258c63643f5a45f757f7509c4e913696c31a4a85ad63c7e57c0f9667a7bcfb9c4b67953f2b991201f71622d15dbe35b271738576cfdd999f7d40dc19f7ec6fa18d5b758ebe998dd529aff7652caf0e3cb4a6915d06f166;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1299bfea1dd8a163ce4ed34590a559c3451ea4aa3b911625d25b207d5c10bd8def9f56d331cec3a594ef7c985cc7f0e114688222ba243153f929b2f65be6f67f86b61ac10b620731e4bf79426e8ab765cce29c3529bce578083159c573f85081a4cc1b79f6b59e2f448df6a3cea4d1f91fc20be8368c4610f;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72543ca3d650ae93e49254fe5317b7ae488110edcbf2ae995cbac0c9fccd433006518b79b5144ff63627c29449a48c0e8d1e355b47982638ac46729aa1b9fcbb7a4f77f3c7088e9f220a84763fe0d572ad1a7c127e161bbdedeb058685e5d53986a4f095ab4609f49e832d972f48476a7a2c7d7da5e81110;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1857f75d6a500ff0ebc994283a257ad26b06a81c0165ef38acd38b8e7a11105e82ee8012dea46d0064116645f28afd280c970cd0eee34047f7d8d80a256c6082de174132f5005b90bc6f5f6ca5ee5ee0a69517717504a171fb48be24b482b8b91867bcc3e92529a01f96a528ad71c2a5f2a2d63ec50b82a3d;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9f11bb50292b6f16eb9983cdcdee0f0067e32363d555e8dc92a3f69dd01c65cd7fe9797c3ccd154f5ea685539bdcdf630853e45313294d4ae979a38ba607c940d62a8adb4fe414f557394dd532b70c76ced942808e55448dc7bcaa06140029b953882fcc9701296437d5002f68ba06df57d7ef3c8476da3;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d0586b683ef797c59b0afff456863d070fb925d5a3d035720f1ec0167c3f3667f4788afc6560e3843d38e2ec948bad1b1ac189a0019e614a974cd96076bed5373b68944e484145dd4c01eb1921a3ccbab088f826b4bef13eca57b049b41b50dd488cd47e3aef20d2c6b93d4b13ff76055f39243aeebbda2b;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b016049ed26a39a0e3d2c491839609004c53930de57e10fd6acbfbeaa4fffda517a5bda1214754b691c4b5fb3b1db4f07346f84349bae4adfd45a1889717fc7a004d7a7fbad343248390f79a8ff938c3f606a55d02ae0bad58e68a8e345cb39e83d15342ee54a65159e813bf0cf76a25cbe5ac2d5894dd01;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f7bba8f55ac447934b0f5dfcc8bf53c178ca8cb1fff7a422a74cb799350ee402077666d00ec4b9503be4f86d6d0f0221519412c5587739d1c0df6dc0cb654002d97e2f9d4c7e7d2044ddb8310010a5a680599daa15af7bbf5f6c8cb12deb771cb4997554e93e51637c9d7da1b87e5cd76539350b32829b2;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf4d0b2c53782df106360be3dec179441fff6b32867a6a14cdb2b0b736e8b20e6e6fe77e8c96bc151b5d4b52bf35b5b7b748c0145ce65af13924f27f234dc83aa71da973225045f29e7cca76bf789e762034e9e5917e2ee89640c2c0340e41128026f1a27e0c6853144120c956c1ccb4d3e459e8cee89111;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h936f862f5088eccac954a6f891373e16a25454d5c22d0f6a1529d14cfcc1e727689faeda69ae39c97306a2c6f39d83454ad7f2f4d089156e209d55108f69e4ddf949943dae2520537c147b3a5796c84888dbe485cf19cc954aaabda69a888562c798c2e909736299a60459599fd710b07004e5a631ad15ad;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c2ad35d181d68285c8b327f3966bff429b279aa2d3630c6dd26ad5177dace0f70787186352d97d2be7ce334d67e590304c15b33cd8dd48162403f35842f7e6c56e418e7d1fb5d595deac3c3a330110b2da2a80760b8fdda721ff21ef9325c7233ff626b439ad471b5d061af63a4683974f07e9821761d89;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h30ffeb7af5e53888ee503ee7d21cd3a1aa5869c219fa717c14270fdd7dac941eff397264ee0e1b3666df54d7a1fe25bdaee301307453dd78b13d2efd8016b208e20545748a2c5e3fcf6fe630287cd6db574b987ce5fafac568082d4c424329e7f410a432b51228586db837870b1ba0f90e860e650de96d69;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eff42c4045e5364d51f507044f7c6ff4bb6e377f80bd4331a2a7287b786c77025b9a766fd1046bd7b699c582c28e8b7f2f031a4e44a06b696ef4701c7be111919e33a9419d6bf428c76cb5c8b10f3b73048e6d0805be5514575e364527a5f8d928192e02f261228de0a0e1d08f24f3341258bd40756c3972;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h744c972df083799f2be242c1ed538836626603c21a55cac79a23daf33ac38395cc7495f6f43032ff55c2eb006cb920b7ae28531a5b7100284d6157e99fbc5d978514b02fe0055654f5f063044580d7f5785f7d058e5e27fb12b263c04b9ef3c4764aaa19de6010c87b0e93d150996be57bf2f6822f6d4382;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he4eefb6e48f189d713cf7ff32eebc9ce1fa04715d5747260b1a84ec50d68e799818df49e32319220327b676d8fd84f7b4ea5db1f20b55167fa83857c074036f5d2652f315754f1714941342d86ceef2c63608597ab94f86ce2cba20c4fb97f3fcd97858022ea7b79f2037714962ea30b5fc3193af606adc9;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68af0c1b238af204ef614f1e9c523fa5df8eca879605b7074df91e00b27b6ea7a675cdaaa9b2dd811227ea5ed9a1bf3ad843bfd906b771e3cfe7e9833f0594a6b89cb2d76466a80e113a694c6b0eeb24b3ada967df9c46945ea009f560a5b2777e21deb75cea6666de3673d768303ced2c0bd1615869e9d1;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11263c2b1df3fe8abdb963d5feae2e484af62fe0308a750c7cab0f22efd4ad1bff0607e9107b12cb7983f47ff524b65c05f28ef5f4144a205899b419a1167fcd6e8392e7516d2c41d951276822e2aca9b48ccc6447ea012fd942d001f6d447e452b05a78960cf93b1f1a05d7ae9d5fa2ed134c075b2c01bbd;
        #1
        {src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14af06df7dc64cf359c6e7d245b9609c1aa411716908fab369d529bf5dcaf7cfd98bf77c5898512d6f472119593db37db4e6ef0349ebfde4fa6e1bbe6dda22dbf26a6de67c1742a11676aa67788e2c45ca555c6489479e6f8264bc40da9b7bfffe691b503ac141d82e453a3d129fcd5ba781f05211b47b664;
        #1
        $finish();
    end
endmodule
