module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    compressor2_1_256_32 compressor2_1_256_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
        src16 <= 256'h0;
        src17 <= 256'h0;
        src18 <= 256'h0;
        src19 <= 256'h0;
        src20 <= 256'h0;
        src21 <= 256'h0;
        src22 <= 256'h0;
        src23 <= 256'h0;
        src24 <= 256'h0;
        src25 <= 256'h0;
        src26 <= 256'h0;
        src27 <= 256'h0;
        src28 <= 256'h0;
        src29 <= 256'h0;
        src30 <= 256'h0;
        src31 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor2_1_256_32(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    input [255:0]src16,
    input [255:0]src17,
    input [255:0]src18,
    input [255:0]src19,
    input [255:0]src20,
    input [255:0]src21,
    input [255:0]src22,
    input [255:0]src23,
    input [255:0]src24,
    input [255:0]src25,
    input [255:0]src26,
    input [255:0]src27,
    input [255:0]src28,
    input [255:0]src29,
    input [255:0]src30,
    input [255:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [0:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [0:0] comp_out38;
    wire [0:0] comp_out39;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39)
    );
    rowadder2_1_40 rowadder2_1inst(
        .src0({comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], 1'h0, comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, comp_out2[1], comp_out1[1], 1'h0}),
        .dst0({dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      input wire [255:0] src16,
      input wire [255:0] src17,
      input wire [255:0] src18,
      input wire [255:0] src19,
      input wire [255:0] src20,
      input wire [255:0] src21,
      input wire [255:0] src22,
      input wire [255:0] src23,
      input wire [255:0] src24,
      input wire [255:0] src25,
      input wire [255:0] src26,
      input wire [255:0] src27,
      input wire [255:0] src28,
      input wire [255:0] src29,
      input wire [255:0] src30,
      input wire [255:0] src31,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [0:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [0:0] dst38,
      output wire [0:0] dst39);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [255:0] stage0_16;
   wire [255:0] stage0_17;
   wire [255:0] stage0_18;
   wire [255:0] stage0_19;
   wire [255:0] stage0_20;
   wire [255:0] stage0_21;
   wire [255:0] stage0_22;
   wire [255:0] stage0_23;
   wire [255:0] stage0_24;
   wire [255:0] stage0_25;
   wire [255:0] stage0_26;
   wire [255:0] stage0_27;
   wire [255:0] stage0_28;
   wire [255:0] stage0_29;
   wire [255:0] stage0_30;
   wire [255:0] stage0_31;
   wire [49:0] stage1_0;
   wire [97:0] stage1_1;
   wire [91:0] stage1_2;
   wire [90:0] stage1_3;
   wire [148:0] stage1_4;
   wire [125:0] stage1_5;
   wire [95:0] stage1_6;
   wire [100:0] stage1_7;
   wire [119:0] stage1_8;
   wire [131:0] stage1_9;
   wire [96:0] stage1_10;
   wire [139:0] stage1_11;
   wire [197:0] stage1_12;
   wire [92:0] stage1_13;
   wire [113:0] stage1_14;
   wire [92:0] stage1_15;
   wire [95:0] stage1_16;
   wire [126:0] stage1_17;
   wire [150:0] stage1_18;
   wire [93:0] stage1_19;
   wire [115:0] stage1_20;
   wire [138:0] stage1_21;
   wire [93:0] stage1_22;
   wire [93:0] stage1_23;
   wire [253:0] stage1_24;
   wire [117:0] stage1_25;
   wire [236:0] stage1_26;
   wire [107:0] stage1_27;
   wire [101:0] stage1_28;
   wire [117:0] stage1_29;
   wire [96:0] stage1_30;
   wire [132:0] stage1_31;
   wire [73:0] stage1_32;
   wire [33:0] stage1_33;
   wire [23:0] stage2_0;
   wire [32:0] stage2_1;
   wire [34:0] stage2_2;
   wire [42:0] stage2_3;
   wire [73:0] stage2_4;
   wire [41:0] stage2_5;
   wire [52:0] stage2_6;
   wire [53:0] stage2_7;
   wire [55:0] stage2_8;
   wire [65:0] stage2_9;
   wire [48:0] stage2_10;
   wire [57:0] stage2_11;
   wire [74:0] stage2_12;
   wire [56:0] stage2_13;
   wire [89:0] stage2_14;
   wire [46:0] stage2_15;
   wire [40:0] stage2_16;
   wire [54:0] stage2_17;
   wire [90:0] stage2_18;
   wire [45:0] stage2_19;
   wire [125:0] stage2_20;
   wire [71:0] stage2_21;
   wire [46:0] stage2_22;
   wire [56:0] stage2_23;
   wire [63:0] stage2_24;
   wire [65:0] stage2_25;
   wire [67:0] stage2_26;
   wire [95:0] stage2_27;
   wire [71:0] stage2_28;
   wire [39:0] stage2_29;
   wire [44:0] stage2_30;
   wire [47:0] stage2_31;
   wire [43:0] stage2_32;
   wire [30:0] stage2_33;
   wire [16:0] stage2_34;
   wire [5:0] stage2_35;
   wire [5:0] stage3_0;
   wire [27:0] stage3_1;
   wire [24:0] stage3_2;
   wire [34:0] stage3_3;
   wire [35:0] stage3_4;
   wire [15:0] stage3_5;
   wire [19:0] stage3_6;
   wire [23:0] stage3_7;
   wire [26:0] stage3_8;
   wire [21:0] stage3_9;
   wire [18:0] stage3_10;
   wire [25:0] stage3_11;
   wire [31:0] stage3_12;
   wire [36:0] stage3_13;
   wire [25:0] stage3_14;
   wire [32:0] stage3_15;
   wire [26:0] stage3_16;
   wire [19:0] stage3_17;
   wire [37:0] stage3_18;
   wire [34:0] stage3_19;
   wire [36:0] stage3_20;
   wire [32:0] stage3_21;
   wire [34:0] stage3_22;
   wire [20:0] stage3_23;
   wire [23:0] stage3_24;
   wire [35:0] stage3_25;
   wire [23:0] stage3_26;
   wire [38:0] stage3_27;
   wire [44:0] stage3_28;
   wire [27:0] stage3_29;
   wire [17:0] stage3_30;
   wire [36:0] stage3_31;
   wire [19:0] stage3_32;
   wire [17:0] stage3_33;
   wire [9:0] stage3_34;
   wire [12:0] stage3_35;
   wire [2:0] stage3_36;
   wire [5:0] stage4_0;
   wire [12:0] stage4_1;
   wire [7:0] stage4_2;
   wire [11:0] stage4_3;
   wire [15:0] stage4_4;
   wire [11:0] stage4_5;
   wire [14:0] stage4_6;
   wire [14:0] stage4_7;
   wire [7:0] stage4_8;
   wire [9:0] stage4_9;
   wire [14:0] stage4_10;
   wire [10:0] stage4_11;
   wire [11:0] stage4_12;
   wire [20:0] stage4_13;
   wire [11:0] stage4_14;
   wire [16:0] stage4_15;
   wire [18:0] stage4_16;
   wire [7:0] stage4_17;
   wire [13:0] stage4_18;
   wire [13:0] stage4_19;
   wire [18:0] stage4_20;
   wire [11:0] stage4_21;
   wire [24:0] stage4_22;
   wire [10:0] stage4_23;
   wire [7:0] stage4_24;
   wire [11:0] stage4_25;
   wire [15:0] stage4_26;
   wire [16:0] stage4_27;
   wire [19:0] stage4_28;
   wire [23:0] stage4_29;
   wire [9:0] stage4_30;
   wire [16:0] stage4_31;
   wire [9:0] stage4_32;
   wire [8:0] stage4_33;
   wire [5:0] stage4_34;
   wire [11:0] stage4_35;
   wire [5:0] stage4_36;
   wire [0:0] stage4_37;
   wire [0:0] stage5_0;
   wire [3:0] stage5_1;
   wire [4:0] stage5_2;
   wire [2:0] stage5_3;
   wire [8:0] stage5_4;
   wire [5:0] stage5_5;
   wire [6:0] stage5_6;
   wire [6:0] stage5_7;
   wire [6:0] stage5_8;
   wire [12:0] stage5_9;
   wire [5:0] stage5_10;
   wire [6:0] stage5_11;
   wire [3:0] stage5_12;
   wire [7:0] stage5_13;
   wire [6:0] stage5_14;
   wire [8:0] stage5_15;
   wire [5:0] stage5_16;
   wire [7:0] stage5_17;
   wire [5:0] stage5_18;
   wire [6:0] stage5_19;
   wire [9:0] stage5_20;
   wire [5:0] stage5_21;
   wire [7:0] stage5_22;
   wire [6:0] stage5_23;
   wire [5:0] stage5_24;
   wire [2:0] stage5_25;
   wire [5:0] stage5_26;
   wire [7:0] stage5_27;
   wire [5:0] stage5_28;
   wire [6:0] stage5_29;
   wire [12:0] stage5_30;
   wire [5:0] stage5_31;
   wire [5:0] stage5_32;
   wire [5:0] stage5_33;
   wire [3:0] stage5_34;
   wire [7:0] stage5_35;
   wire [7:0] stage5_36;
   wire [1:0] stage5_37;
   wire [0:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [0:0] stage6_3;
   wire [3:0] stage6_4;
   wire [2:0] stage6_5;
   wire [2:0] stage6_6;
   wire [2:0] stage6_7;
   wire [4:0] stage6_8;
   wire [3:0] stage6_9;
   wire [5:0] stage6_10;
   wire [2:0] stage6_11;
   wire [5:0] stage6_12;
   wire [2:0] stage6_13;
   wire [3:0] stage6_14;
   wire [3:0] stage6_15;
   wire [1:0] stage6_16;
   wire [2:0] stage6_17;
   wire [4:0] stage6_18;
   wire [1:0] stage6_19;
   wire [5:0] stage6_20;
   wire [2:0] stage6_21;
   wire [5:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [2:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [2:0] stage6_28;
   wire [3:0] stage6_29;
   wire [5:0] stage6_30;
   wire [2:0] stage6_31;
   wire [2:0] stage6_32;
   wire [2:0] stage6_33;
   wire [2:0] stage6_34;
   wire [2:0] stage6_35;
   wire [3:0] stage6_36;
   wire [3:0] stage6_37;
   wire [0:0] stage6_38;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [0:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [0:0] stage7_25;
   wire [1:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [1:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [1:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [0:0] stage7_38;
   wire [0:0] stage7_39;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc135_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc135_4 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1406_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[7]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[8]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[3],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[4],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[5],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[6],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[7],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[8],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[9],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[10],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[11],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[12],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[13],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[14],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[15],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[16],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[17],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[18],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[19],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[20],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[21],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[22],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[23],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[24],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[25],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[26],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[27],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[28],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[29],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[30],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[31],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[32],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[33],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[34],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[35],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[36],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[37],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[38],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[39],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[40],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[41],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[42],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[43],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[44],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[45],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[46],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[47],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[48],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[49],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[50],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[51],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[52],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[53],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[54],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[55],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[56],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[57],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[18],stage1_4[58],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[19],stage1_4[59],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[20],stage1_4[60],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[21],stage1_4[61],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[22],stage1_4[62],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[23],stage1_4[63],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[24],stage1_4[64],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[25],stage1_4[65],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[26],stage1_4[66],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[27],stage1_4[67],stage1_3[70],stage1_2[70],stage1_1[70]}
   );
   gpc606_5 gpc71 (
      {stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[28],stage1_4[68],stage1_3[71],stage1_2[71],stage1_1[71]}
   );
   gpc606_5 gpc72 (
      {stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[29],stage1_4[69],stage1_3[72],stage1_2[72],stage1_1[72]}
   );
   gpc606_5 gpc73 (
      {stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[30],stage1_4[70],stage1_3[73],stage1_2[73],stage1_1[73]}
   );
   gpc606_5 gpc74 (
      {stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[31],stage1_4[71],stage1_3[74],stage1_2[74],stage1_1[74]}
   );
   gpc606_5 gpc75 (
      {stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[32],stage1_4[72],stage1_3[75],stage1_2[75],stage1_1[75]}
   );
   gpc606_5 gpc76 (
      {stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[33],stage1_4[73],stage1_3[76],stage1_2[76],stage1_1[76]}
   );
   gpc606_5 gpc77 (
      {stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[34],stage1_4[74],stage1_3[77],stage1_2[77],stage1_1[77]}
   );
   gpc606_5 gpc78 (
      {stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[35],stage1_4[75],stage1_3[78],stage1_2[78],stage1_1[78]}
   );
   gpc606_5 gpc79 (
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[36],stage1_4[76],stage1_3[79],stage1_2[79]}
   );
   gpc606_5 gpc80 (
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[37],stage1_4[77],stage1_3[80],stage1_2[80]}
   );
   gpc623_5 gpc81 (
      {stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage0_3[219], stage0_3[220]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[38],stage1_4[78],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225]},
      {stage0_4[18]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[39],stage1_4[79],stage1_3[82]}
   );
   gpc615_5 gpc83 (
      {stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230]},
      {stage0_4[19]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[40],stage1_4[80],stage1_3[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235]},
      {stage0_4[20]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[5],stage1_5[41],stage1_4[81],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage0_4[21]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[6],stage1_5[42],stage1_4[82],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245]},
      {stage0_4[22]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[7],stage1_5[43],stage1_4[83],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage0_4[23]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[8],stage1_5[44],stage1_4[84],stage1_3[87]}
   );
   gpc623_5 gpc88 (
      {stage0_3[251], stage0_3[252], stage0_3[253]},
      {stage0_4[24], stage0_4[25]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[9],stage1_5[45],stage1_4[85],stage1_3[88]}
   );
   gpc1163_5 gpc89 (
      {stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_6[0]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[7],stage1_6[10],stage1_5[46],stage1_4[86]}
   );
   gpc1163_5 gpc90 (
      {stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[1]},
      {stage0_7[1]},
      {stage1_8[1],stage1_7[8],stage1_6[11],stage1_5[47],stage1_4[87]}
   );
   gpc1163_5 gpc91 (
      {stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_6[2]},
      {stage0_7[2]},
      {stage1_8[2],stage1_7[9],stage1_6[12],stage1_5[48],stage1_4[88]}
   );
   gpc1163_5 gpc92 (
      {stage0_4[35], stage0_4[36], stage0_4[37]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_6[3]},
      {stage0_7[3]},
      {stage1_8[3],stage1_7[10],stage1_6[13],stage1_5[49],stage1_4[89]}
   );
   gpc1163_5 gpc93 (
      {stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_6[4]},
      {stage0_7[4]},
      {stage1_8[4],stage1_7[11],stage1_6[14],stage1_5[50],stage1_4[90]}
   );
   gpc1163_5 gpc94 (
      {stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_6[5]},
      {stage0_7[5]},
      {stage1_8[5],stage1_7[12],stage1_6[15],stage1_5[51],stage1_4[91]}
   );
   gpc606_5 gpc95 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[6],stage1_7[13],stage1_6[16],stage1_5[52],stage1_4[92]}
   );
   gpc606_5 gpc96 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[7],stage1_7[14],stage1_6[17],stage1_5[53],stage1_4[93]}
   );
   gpc606_5 gpc97 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[8],stage1_7[15],stage1_6[18],stage1_5[54],stage1_4[94]}
   );
   gpc606_5 gpc98 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[9],stage1_7[16],stage1_6[19],stage1_5[55],stage1_4[95]}
   );
   gpc606_5 gpc99 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[10],stage1_7[17],stage1_6[20],stage1_5[56],stage1_4[96]}
   );
   gpc606_5 gpc100 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[11],stage1_7[18],stage1_6[21],stage1_5[57],stage1_4[97]}
   );
   gpc606_5 gpc101 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[12],stage1_7[19],stage1_6[22],stage1_5[58],stage1_4[98]}
   );
   gpc606_5 gpc102 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[13],stage1_7[20],stage1_6[23],stage1_5[59],stage1_4[99]}
   );
   gpc606_5 gpc103 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[14],stage1_7[21],stage1_6[24],stage1_5[60],stage1_4[100]}
   );
   gpc606_5 gpc104 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[15],stage1_7[22],stage1_6[25],stage1_5[61],stage1_4[101]}
   );
   gpc606_5 gpc105 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[16],stage1_7[23],stage1_6[26],stage1_5[62],stage1_4[102]}
   );
   gpc606_5 gpc106 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[17],stage1_7[24],stage1_6[27],stage1_5[63],stage1_4[103]}
   );
   gpc606_5 gpc107 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[18],stage1_7[25],stage1_6[28],stage1_5[64],stage1_4[104]}
   );
   gpc606_5 gpc108 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[19],stage1_7[26],stage1_6[29],stage1_5[65],stage1_4[105]}
   );
   gpc606_5 gpc109 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[20],stage1_7[27],stage1_6[30],stage1_5[66],stage1_4[106]}
   );
   gpc606_5 gpc110 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[21],stage1_7[28],stage1_6[31],stage1_5[67],stage1_4[107]}
   );
   gpc606_5 gpc111 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[22],stage1_7[29],stage1_6[32],stage1_5[68],stage1_4[108]}
   );
   gpc606_5 gpc112 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[23],stage1_7[30],stage1_6[33],stage1_5[69],stage1_4[109]}
   );
   gpc606_5 gpc113 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[24],stage1_7[31],stage1_6[34],stage1_5[70],stage1_4[110]}
   );
   gpc606_5 gpc114 (
      {stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[25],stage1_7[32],stage1_6[35],stage1_5[71],stage1_4[111]}
   );
   gpc606_5 gpc115 (
      {stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[26],stage1_7[33],stage1_6[36],stage1_5[72],stage1_4[112]}
   );
   gpc606_5 gpc116 (
      {stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[27],stage1_7[34],stage1_6[37],stage1_5[73],stage1_4[113]}
   );
   gpc606_5 gpc117 (
      {stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[28],stage1_7[35],stage1_6[38],stage1_5[74],stage1_4[114]}
   );
   gpc606_5 gpc118 (
      {stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[29],stage1_7[36],stage1_6[39],stage1_5[75],stage1_4[115]}
   );
   gpc606_5 gpc119 (
      {stage0_4[188], stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[30],stage1_7[37],stage1_6[40],stage1_5[76],stage1_4[116]}
   );
   gpc606_5 gpc120 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[31],stage1_7[38],stage1_6[41],stage1_5[77],stage1_4[117]}
   );
   gpc606_5 gpc121 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[32],stage1_7[39],stage1_6[42],stage1_5[78],stage1_4[118]}
   );
   gpc606_5 gpc122 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[33],stage1_7[40],stage1_6[43],stage1_5[79],stage1_4[119]}
   );
   gpc606_5 gpc123 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[34],stage1_7[41],stage1_6[44],stage1_5[80],stage1_4[120]}
   );
   gpc606_5 gpc124 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[35],stage1_7[42],stage1_6[45],stage1_5[81],stage1_4[121]}
   );
   gpc606_5 gpc125 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[36],stage1_7[43],stage1_6[46],stage1_5[82],stage1_4[122]}
   );
   gpc606_5 gpc126 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[0],stage1_8[37],stage1_7[44],stage1_6[47],stage1_5[83]}
   );
   gpc606_5 gpc127 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[1],stage1_8[38],stage1_7[45],stage1_6[48],stage1_5[84]}
   );
   gpc606_5 gpc128 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[2],stage1_8[39],stage1_7[46],stage1_6[49],stage1_5[85]}
   );
   gpc606_5 gpc129 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[3],stage1_8[40],stage1_7[47],stage1_6[50],stage1_5[86]}
   );
   gpc606_5 gpc130 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[4],stage1_8[41],stage1_7[48],stage1_6[51],stage1_5[87]}
   );
   gpc606_5 gpc131 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[5],stage1_8[42],stage1_7[49],stage1_6[52],stage1_5[88]}
   );
   gpc606_5 gpc132 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[6],stage1_8[43],stage1_7[50],stage1_6[53],stage1_5[89]}
   );
   gpc606_5 gpc133 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[7],stage1_8[44],stage1_7[51],stage1_6[54],stage1_5[90]}
   );
   gpc606_5 gpc134 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[8],stage1_8[45],stage1_7[52],stage1_6[55],stage1_5[91]}
   );
   gpc606_5 gpc135 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[9],stage1_8[46],stage1_7[53],stage1_6[56],stage1_5[92]}
   );
   gpc606_5 gpc136 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[10],stage1_8[47],stage1_7[54],stage1_6[57],stage1_5[93]}
   );
   gpc606_5 gpc137 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[11],stage1_8[48],stage1_7[55],stage1_6[58],stage1_5[94]}
   );
   gpc606_5 gpc138 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[12],stage1_8[49],stage1_7[56],stage1_6[59],stage1_5[95]}
   );
   gpc606_5 gpc139 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[13],stage1_8[50],stage1_7[57],stage1_6[60],stage1_5[96]}
   );
   gpc606_5 gpc140 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[14],stage1_8[51],stage1_7[58],stage1_6[61],stage1_5[97]}
   );
   gpc606_5 gpc141 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[15],stage1_8[52],stage1_7[59],stage1_6[62],stage1_5[98]}
   );
   gpc606_5 gpc142 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[16],stage1_8[53],stage1_7[60],stage1_6[63],stage1_5[99]}
   );
   gpc606_5 gpc143 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[17],stage1_8[54],stage1_7[61],stage1_6[64],stage1_5[100]}
   );
   gpc606_5 gpc144 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[18],stage1_8[55],stage1_7[62],stage1_6[65],stage1_5[101]}
   );
   gpc606_5 gpc145 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[19],stage1_8[56],stage1_7[63],stage1_6[66],stage1_5[102]}
   );
   gpc606_5 gpc146 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[20],stage1_8[57],stage1_7[64],stage1_6[67],stage1_5[103]}
   );
   gpc606_5 gpc147 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[21],stage1_8[58],stage1_7[65],stage1_6[68],stage1_5[104]}
   );
   gpc606_5 gpc148 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[22],stage1_8[59],stage1_7[66],stage1_6[69],stage1_5[105]}
   );
   gpc606_5 gpc149 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[23],stage1_8[60],stage1_7[67],stage1_6[70],stage1_5[106]}
   );
   gpc606_5 gpc150 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[24],stage1_8[61],stage1_7[68],stage1_6[71],stage1_5[107]}
   );
   gpc606_5 gpc151 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[25],stage1_8[62],stage1_7[69],stage1_6[72],stage1_5[108]}
   );
   gpc606_5 gpc152 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[26],stage1_8[63],stage1_7[70],stage1_6[73],stage1_5[109]}
   );
   gpc606_5 gpc153 (
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[64],stage1_7[71],stage1_6[74]}
   );
   gpc606_5 gpc154 (
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[65],stage1_7[72],stage1_6[75]}
   );
   gpc606_5 gpc155 (
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[66],stage1_7[73],stage1_6[76]}
   );
   gpc606_5 gpc156 (
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[67],stage1_7[74],stage1_6[77]}
   );
   gpc606_5 gpc157 (
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[68],stage1_7[75],stage1_6[78]}
   );
   gpc606_5 gpc158 (
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[69],stage1_7[76],stage1_6[79]}
   );
   gpc615_5 gpc159 (
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232]},
      {stage0_7[168]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[33],stage1_8[70],stage1_7[77],stage1_6[80]}
   );
   gpc615_5 gpc160 (
      {stage0_6[233], stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237]},
      {stage0_7[169]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[34],stage1_8[71],stage1_7[78],stage1_6[81]}
   );
   gpc615_5 gpc161 (
      {stage0_6[238], stage0_6[239], stage0_6[240], stage0_6[241], stage0_6[242]},
      {stage0_7[170]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[35],stage1_8[72],stage1_7[79],stage1_6[82]}
   );
   gpc615_5 gpc162 (
      {stage0_7[171], stage0_7[172], stage0_7[173], stage0_7[174], stage0_7[175]},
      {stage0_8[54]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[9],stage1_9[36],stage1_8[73],stage1_7[80]}
   );
   gpc615_5 gpc163 (
      {stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179], stage0_7[180]},
      {stage0_8[55]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[10],stage1_9[37],stage1_8[74],stage1_7[81]}
   );
   gpc615_5 gpc164 (
      {stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage0_8[56]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[11],stage1_9[38],stage1_8[75],stage1_7[82]}
   );
   gpc615_5 gpc165 (
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190]},
      {stage0_8[57]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[12],stage1_9[39],stage1_8[76],stage1_7[83]}
   );
   gpc615_5 gpc166 (
      {stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_8[58]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[13],stage1_9[40],stage1_8[77],stage1_7[84]}
   );
   gpc615_5 gpc167 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[59]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[14],stage1_9[41],stage1_8[78],stage1_7[85]}
   );
   gpc615_5 gpc168 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[60]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[15],stage1_9[42],stage1_8[79],stage1_7[86]}
   );
   gpc615_5 gpc169 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[61]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[16],stage1_9[43],stage1_8[80],stage1_7[87]}
   );
   gpc615_5 gpc170 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[62]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[17],stage1_9[44],stage1_8[81],stage1_7[88]}
   );
   gpc615_5 gpc171 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[63]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[18],stage1_9[45],stage1_8[82],stage1_7[89]}
   );
   gpc615_5 gpc172 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[64]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[19],stage1_9[46],stage1_8[83],stage1_7[90]}
   );
   gpc615_5 gpc173 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[65]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[20],stage1_9[47],stage1_8[84],stage1_7[91]}
   );
   gpc615_5 gpc174 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[66]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[21],stage1_9[48],stage1_8[85],stage1_7[92]}
   );
   gpc615_5 gpc175 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[67]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[22],stage1_9[49],stage1_8[86],stage1_7[93]}
   );
   gpc615_5 gpc176 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[68]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[23],stage1_9[50],stage1_8[87],stage1_7[94]}
   );
   gpc615_5 gpc177 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[69]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[24],stage1_9[51],stage1_8[88],stage1_7[95]}
   );
   gpc606_5 gpc178 (
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[16],stage1_10[25],stage1_9[52],stage1_8[89]}
   );
   gpc606_5 gpc179 (
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[17],stage1_10[26],stage1_9[53],stage1_8[90]}
   );
   gpc606_5 gpc180 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[18],stage1_10[27],stage1_9[54],stage1_8[91]}
   );
   gpc606_5 gpc181 (
      {stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[19],stage1_10[28],stage1_9[55],stage1_8[92]}
   );
   gpc606_5 gpc182 (
      {stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[20],stage1_10[29],stage1_9[56],stage1_8[93]}
   );
   gpc606_5 gpc183 (
      {stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[21],stage1_10[30],stage1_9[57],stage1_8[94]}
   );
   gpc606_5 gpc184 (
      {stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[22],stage1_10[31],stage1_9[58],stage1_8[95]}
   );
   gpc606_5 gpc185 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[23],stage1_10[32],stage1_9[59],stage1_8[96]}
   );
   gpc606_5 gpc186 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[24],stage1_10[33],stage1_9[60],stage1_8[97]}
   );
   gpc606_5 gpc187 (
      {stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[25],stage1_10[34],stage1_9[61],stage1_8[98]}
   );
   gpc606_5 gpc188 (
      {stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[26],stage1_10[35],stage1_9[62],stage1_8[99]}
   );
   gpc606_5 gpc189 (
      {stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[27],stage1_10[36],stage1_9[63],stage1_8[100]}
   );
   gpc606_5 gpc190 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[28],stage1_10[37],stage1_9[64],stage1_8[101]}
   );
   gpc606_5 gpc191 (
      {stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[29],stage1_10[38],stage1_9[65],stage1_8[102]}
   );
   gpc606_5 gpc192 (
      {stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[30],stage1_10[39],stage1_9[66],stage1_8[103]}
   );
   gpc606_5 gpc193 (
      {stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[31],stage1_10[40],stage1_9[67],stage1_8[104]}
   );
   gpc606_5 gpc194 (
      {stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[32],stage1_10[41],stage1_9[68],stage1_8[105]}
   );
   gpc606_5 gpc195 (
      {stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[33],stage1_10[42],stage1_9[69],stage1_8[106]}
   );
   gpc606_5 gpc196 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[34],stage1_10[43],stage1_9[70],stage1_8[107]}
   );
   gpc606_5 gpc197 (
      {stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[35],stage1_10[44],stage1_9[71],stage1_8[108]}
   );
   gpc606_5 gpc198 (
      {stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[36],stage1_10[45],stage1_9[72],stage1_8[109]}
   );
   gpc606_5 gpc199 (
      {stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[37],stage1_10[46],stage1_9[73],stage1_8[110]}
   );
   gpc606_5 gpc200 (
      {stage0_8[202], stage0_8[203], stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[38],stage1_10[47],stage1_9[74],stage1_8[111]}
   );
   gpc606_5 gpc201 (
      {stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[39],stage1_10[48],stage1_9[75],stage1_8[112]}
   );
   gpc606_5 gpc202 (
      {stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[40],stage1_10[49],stage1_9[76],stage1_8[113]}
   );
   gpc606_5 gpc203 (
      {stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[41],stage1_10[50],stage1_9[77],stage1_8[114]}
   );
   gpc606_5 gpc204 (
      {stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[42],stage1_10[51],stage1_9[78],stage1_8[115]}
   );
   gpc606_5 gpc205 (
      {stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[43],stage1_10[52],stage1_9[79],stage1_8[116]}
   );
   gpc606_5 gpc206 (
      {stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[44],stage1_10[53],stage1_9[80],stage1_8[117]}
   );
   gpc606_5 gpc207 (
      {stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[45],stage1_10[54],stage1_9[81],stage1_8[118]}
   );
   gpc606_5 gpc208 (
      {stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[46],stage1_10[55],stage1_9[82],stage1_8[119]}
   );
   gpc606_5 gpc209 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[31],stage1_11[47],stage1_10[56],stage1_9[83]}
   );
   gpc606_5 gpc210 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[32],stage1_11[48],stage1_10[57],stage1_9[84]}
   );
   gpc606_5 gpc211 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[33],stage1_11[49],stage1_10[58],stage1_9[85]}
   );
   gpc606_5 gpc212 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[34],stage1_11[50],stage1_10[59],stage1_9[86]}
   );
   gpc606_5 gpc213 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[35],stage1_11[51],stage1_10[60],stage1_9[87]}
   );
   gpc606_5 gpc214 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[36],stage1_11[52],stage1_10[61],stage1_9[88]}
   );
   gpc606_5 gpc215 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[37],stage1_11[53],stage1_10[62],stage1_9[89]}
   );
   gpc606_5 gpc216 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[38],stage1_11[54],stage1_10[63],stage1_9[90]}
   );
   gpc606_5 gpc217 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[39],stage1_11[55],stage1_10[64],stage1_9[91]}
   );
   gpc606_5 gpc218 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[40],stage1_11[56],stage1_10[65],stage1_9[92]}
   );
   gpc606_5 gpc219 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[41],stage1_11[57],stage1_10[66],stage1_9[93]}
   );
   gpc606_5 gpc220 (
      {stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[42],stage1_11[58],stage1_10[67],stage1_9[94]}
   );
   gpc606_5 gpc221 (
      {stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[43],stage1_11[59],stage1_10[68],stage1_9[95]}
   );
   gpc606_5 gpc222 (
      {stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[44],stage1_11[60],stage1_10[69],stage1_9[96]}
   );
   gpc606_5 gpc223 (
      {stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[45],stage1_11[61],stage1_10[70],stage1_9[97]}
   );
   gpc606_5 gpc224 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[46],stage1_11[62],stage1_10[71],stage1_9[98]}
   );
   gpc606_5 gpc225 (
      {stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[47],stage1_11[63],stage1_10[72],stage1_9[99]}
   );
   gpc606_5 gpc226 (
      {stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[48],stage1_11[64],stage1_10[73],stage1_9[100]}
   );
   gpc606_5 gpc227 (
      {stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[49],stage1_11[65],stage1_10[74],stage1_9[101]}
   );
   gpc615_5 gpc228 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214]},
      {stage0_10[186]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[50],stage1_11[66],stage1_10[75],stage1_9[102]}
   );
   gpc615_5 gpc229 (
      {stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_10[187]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[51],stage1_11[67],stage1_10[76],stage1_9[103]}
   );
   gpc615_5 gpc230 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_10[188]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[52],stage1_11[68],stage1_10[77],stage1_9[104]}
   );
   gpc615_5 gpc231 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229]},
      {stage0_10[189]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[53],stage1_11[69],stage1_10[78],stage1_9[105]}
   );
   gpc615_5 gpc232 (
      {stage0_10[190], stage0_10[191], stage0_10[192], stage0_10[193], stage0_10[194]},
      {stage0_11[138]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[23],stage1_12[54],stage1_11[70],stage1_10[79]}
   );
   gpc615_5 gpc233 (
      {stage0_10[195], stage0_10[196], stage0_10[197], stage0_10[198], stage0_10[199]},
      {stage0_11[139]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[24],stage1_12[55],stage1_11[71],stage1_10[80]}
   );
   gpc615_5 gpc234 (
      {stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203], stage0_10[204]},
      {stage0_11[140]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[25],stage1_12[56],stage1_11[72],stage1_10[81]}
   );
   gpc615_5 gpc235 (
      {stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage0_11[141]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[26],stage1_12[57],stage1_11[73],stage1_10[82]}
   );
   gpc615_5 gpc236 (
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214]},
      {stage0_11[142]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[27],stage1_12[58],stage1_11[74],stage1_10[83]}
   );
   gpc615_5 gpc237 (
      {stage0_10[215], stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219]},
      {stage0_11[143]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[28],stage1_12[59],stage1_11[75],stage1_10[84]}
   );
   gpc615_5 gpc238 (
      {stage0_10[220], stage0_10[221], stage0_10[222], stage0_10[223], stage0_10[224]},
      {stage0_11[144]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[29],stage1_12[60],stage1_11[76],stage1_10[85]}
   );
   gpc615_5 gpc239 (
      {stage0_10[225], stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229]},
      {stage0_11[145]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[30],stage1_12[61],stage1_11[77],stage1_10[86]}
   );
   gpc615_5 gpc240 (
      {stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234]},
      {stage0_11[146]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[31],stage1_12[62],stage1_11[78],stage1_10[87]}
   );
   gpc615_5 gpc241 (
      {stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage0_11[147]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[32],stage1_12[63],stage1_11[79],stage1_10[88]}
   );
   gpc615_5 gpc242 (
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244]},
      {stage0_11[148]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[33],stage1_12[64],stage1_11[80],stage1_10[89]}
   );
   gpc615_5 gpc243 (
      {stage0_10[245], stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249]},
      {stage0_11[149]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[34],stage1_12[65],stage1_11[81],stage1_10[90]}
   );
   gpc615_5 gpc244 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154]},
      {stage0_12[72]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[12],stage1_13[35],stage1_12[66],stage1_11[82]}
   );
   gpc615_5 gpc245 (
      {stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage0_12[73]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[13],stage1_13[36],stage1_12[67],stage1_11[83]}
   );
   gpc615_5 gpc246 (
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_12[74]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[14],stage1_13[37],stage1_12[68],stage1_11[84]}
   );
   gpc615_5 gpc247 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169]},
      {stage0_12[75]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[15],stage1_13[38],stage1_12[69],stage1_11[85]}
   );
   gpc615_5 gpc248 (
      {stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174]},
      {stage0_12[76]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[16],stage1_13[39],stage1_12[70],stage1_11[86]}
   );
   gpc615_5 gpc249 (
      {stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage0_12[77]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[17],stage1_13[40],stage1_12[71],stage1_11[87]}
   );
   gpc615_5 gpc250 (
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184]},
      {stage0_12[78]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[18],stage1_13[41],stage1_12[72],stage1_11[88]}
   );
   gpc615_5 gpc251 (
      {stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage0_12[79]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[19],stage1_13[42],stage1_12[73],stage1_11[89]}
   );
   gpc615_5 gpc252 (
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194]},
      {stage0_12[80]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[20],stage1_13[43],stage1_12[74],stage1_11[90]}
   );
   gpc615_5 gpc253 (
      {stage0_11[195], stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199]},
      {stage0_12[81]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[21],stage1_13[44],stage1_12[75],stage1_11[91]}
   );
   gpc615_5 gpc254 (
      {stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203], stage0_11[204]},
      {stage0_12[82]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[22],stage1_13[45],stage1_12[76],stage1_11[92]}
   );
   gpc615_5 gpc255 (
      {stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage0_12[83]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[23],stage1_13[46],stage1_12[77],stage1_11[93]}
   );
   gpc117_4 gpc256 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90]},
      {stage0_13[72]},
      {stage0_14[0]},
      {stage1_15[12],stage1_14[24],stage1_13[47],stage1_12[78]}
   );
   gpc606_5 gpc257 (
      {stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96]},
      {stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6]},
      {stage1_16[0],stage1_15[13],stage1_14[25],stage1_13[48],stage1_12[79]}
   );
   gpc606_5 gpc258 (
      {stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102]},
      {stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage1_16[1],stage1_15[14],stage1_14[26],stage1_13[49],stage1_12[80]}
   );
   gpc615_5 gpc259 (
      {stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_13[73]},
      {stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18]},
      {stage1_16[2],stage1_15[15],stage1_14[27],stage1_13[50],stage1_12[81]}
   );
   gpc615_5 gpc260 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112]},
      {stage0_13[74]},
      {stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24]},
      {stage1_16[3],stage1_15[16],stage1_14[28],stage1_13[51],stage1_12[82]}
   );
   gpc615_5 gpc261 (
      {stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage0_13[75]},
      {stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30]},
      {stage1_16[4],stage1_15[17],stage1_14[29],stage1_13[52],stage1_12[83]}
   );
   gpc615_5 gpc262 (
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_13[76]},
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36]},
      {stage1_16[5],stage1_15[18],stage1_14[30],stage1_13[53],stage1_12[84]}
   );
   gpc615_5 gpc263 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_13[77]},
      {stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42]},
      {stage1_16[6],stage1_15[19],stage1_14[31],stage1_13[54],stage1_12[85]}
   );
   gpc615_5 gpc264 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132]},
      {stage0_13[78]},
      {stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47], stage0_14[48]},
      {stage1_16[7],stage1_15[20],stage1_14[32],stage1_13[55],stage1_12[86]}
   );
   gpc615_5 gpc265 (
      {stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_13[79]},
      {stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54]},
      {stage1_16[8],stage1_15[21],stage1_14[33],stage1_13[56],stage1_12[87]}
   );
   gpc615_5 gpc266 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142]},
      {stage0_13[80]},
      {stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60]},
      {stage1_16[9],stage1_15[22],stage1_14[34],stage1_13[57],stage1_12[88]}
   );
   gpc615_5 gpc267 (
      {stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage0_13[81]},
      {stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66]},
      {stage1_16[10],stage1_15[23],stage1_14[35],stage1_13[58],stage1_12[89]}
   );
   gpc606_5 gpc268 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[11],stage1_15[24],stage1_14[36],stage1_13[59]}
   );
   gpc606_5 gpc269 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[12],stage1_15[25],stage1_14[37],stage1_13[60]}
   );
   gpc606_5 gpc270 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[13],stage1_15[26],stage1_14[38],stage1_13[61]}
   );
   gpc606_5 gpc271 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[14],stage1_15[27],stage1_14[39],stage1_13[62]}
   );
   gpc615_5 gpc272 (
      {stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110]},
      {stage0_14[67]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[15],stage1_15[28],stage1_14[40],stage1_13[63]}
   );
   gpc615_5 gpc273 (
      {stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115]},
      {stage0_14[68]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[16],stage1_15[29],stage1_14[41],stage1_13[64]}
   );
   gpc615_5 gpc274 (
      {stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119], stage0_13[120]},
      {stage0_14[69]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[17],stage1_15[30],stage1_14[42],stage1_13[65]}
   );
   gpc615_5 gpc275 (
      {stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_14[70]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[18],stage1_15[31],stage1_14[43],stage1_13[66]}
   );
   gpc615_5 gpc276 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130]},
      {stage0_14[71]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[19],stage1_15[32],stage1_14[44],stage1_13[67]}
   );
   gpc615_5 gpc277 (
      {stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135]},
      {stage0_14[72]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[20],stage1_15[33],stage1_14[45],stage1_13[68]}
   );
   gpc615_5 gpc278 (
      {stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139], stage0_13[140]},
      {stage0_14[73]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[21],stage1_15[34],stage1_14[46],stage1_13[69]}
   );
   gpc615_5 gpc279 (
      {stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145]},
      {stage0_14[74]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[22],stage1_15[35],stage1_14[47],stage1_13[70]}
   );
   gpc615_5 gpc280 (
      {stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150]},
      {stage0_14[75]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[23],stage1_15[36],stage1_14[48],stage1_13[71]}
   );
   gpc615_5 gpc281 (
      {stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_14[76]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[24],stage1_15[37],stage1_14[49],stage1_13[72]}
   );
   gpc615_5 gpc282 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160]},
      {stage0_14[77]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[25],stage1_15[38],stage1_14[50],stage1_13[73]}
   );
   gpc615_5 gpc283 (
      {stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165]},
      {stage0_14[78]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[26],stage1_15[39],stage1_14[51],stage1_13[74]}
   );
   gpc615_5 gpc284 (
      {stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170]},
      {stage0_14[79]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[27],stage1_15[40],stage1_14[52],stage1_13[75]}
   );
   gpc615_5 gpc285 (
      {stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175]},
      {stage0_14[80]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[28],stage1_15[41],stage1_14[53],stage1_13[76]}
   );
   gpc615_5 gpc286 (
      {stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180]},
      {stage0_14[81]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[29],stage1_15[42],stage1_14[54],stage1_13[77]}
   );
   gpc615_5 gpc287 (
      {stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage0_14[82]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[30],stage1_15[43],stage1_14[55],stage1_13[78]}
   );
   gpc615_5 gpc288 (
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190]},
      {stage0_14[83]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[31],stage1_15[44],stage1_14[56],stage1_13[79]}
   );
   gpc615_5 gpc289 (
      {stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195]},
      {stage0_14[84]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[32],stage1_15[45],stage1_14[57],stage1_13[80]}
   );
   gpc615_5 gpc290 (
      {stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_14[85]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[33],stage1_15[46],stage1_14[58],stage1_13[81]}
   );
   gpc615_5 gpc291 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_14[86]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[34],stage1_15[47],stage1_14[59],stage1_13[82]}
   );
   gpc615_5 gpc292 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210]},
      {stage0_14[87]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[35],stage1_15[48],stage1_14[60],stage1_13[83]}
   );
   gpc615_5 gpc293 (
      {stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_14[88]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[36],stage1_15[49],stage1_14[61],stage1_13[84]}
   );
   gpc615_5 gpc294 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220]},
      {stage0_14[89]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[37],stage1_15[50],stage1_14[62],stage1_13[85]}
   );
   gpc615_5 gpc295 (
      {stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_14[90]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[38],stage1_15[51],stage1_14[63],stage1_13[86]}
   );
   gpc615_5 gpc296 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[91]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[39],stage1_15[52],stage1_14[64],stage1_13[87]}
   );
   gpc615_5 gpc297 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[92]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[40],stage1_15[53],stage1_14[65],stage1_13[88]}
   );
   gpc615_5 gpc298 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[93]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[41],stage1_15[54],stage1_14[66],stage1_13[89]}
   );
   gpc615_5 gpc299 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[94]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[42],stage1_15[55],stage1_14[67],stage1_13[90]}
   );
   gpc615_5 gpc300 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[95]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[43],stage1_15[56],stage1_14[68],stage1_13[91]}
   );
   gpc615_5 gpc301 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[96]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[44],stage1_15[57],stage1_14[69],stage1_13[92]}
   );
   gpc606_5 gpc302 (
      {stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[34],stage1_16[45],stage1_15[58],stage1_14[70]}
   );
   gpc606_5 gpc303 (
      {stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[35],stage1_16[46],stage1_15[59],stage1_14[71]}
   );
   gpc606_5 gpc304 (
      {stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113], stage0_14[114]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[36],stage1_16[47],stage1_15[60],stage1_14[72]}
   );
   gpc606_5 gpc305 (
      {stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119], stage0_14[120]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[37],stage1_16[48],stage1_15[61],stage1_14[73]}
   );
   gpc606_5 gpc306 (
      {stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[38],stage1_16[49],stage1_15[62],stage1_14[74]}
   );
   gpc606_5 gpc307 (
      {stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[39],stage1_16[50],stage1_15[63],stage1_14[75]}
   );
   gpc606_5 gpc308 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[40],stage1_16[51],stage1_15[64],stage1_14[76]}
   );
   gpc606_5 gpc309 (
      {stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143], stage0_14[144]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[41],stage1_16[52],stage1_15[65],stage1_14[77]}
   );
   gpc606_5 gpc310 (
      {stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149], stage0_14[150]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[42],stage1_16[53],stage1_15[66],stage1_14[78]}
   );
   gpc606_5 gpc311 (
      {stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[43],stage1_16[54],stage1_15[67],stage1_14[79]}
   );
   gpc606_5 gpc312 (
      {stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161], stage0_14[162]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[44],stage1_16[55],stage1_15[68],stage1_14[80]}
   );
   gpc606_5 gpc313 (
      {stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167], stage0_14[168]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[45],stage1_16[56],stage1_15[69],stage1_14[81]}
   );
   gpc606_5 gpc314 (
      {stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173], stage0_14[174]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[46],stage1_16[57],stage1_15[70],stage1_14[82]}
   );
   gpc606_5 gpc315 (
      {stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179], stage0_14[180]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[47],stage1_16[58],stage1_15[71],stage1_14[83]}
   );
   gpc606_5 gpc316 (
      {stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185], stage0_14[186]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[48],stage1_16[59],stage1_15[72],stage1_14[84]}
   );
   gpc606_5 gpc317 (
      {stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191], stage0_14[192]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[49],stage1_16[60],stage1_15[73],stage1_14[85]}
   );
   gpc606_5 gpc318 (
      {stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197], stage0_14[198]},
      {stage0_16[96], stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101]},
      {stage1_18[16],stage1_17[50],stage1_16[61],stage1_15[74],stage1_14[86]}
   );
   gpc606_5 gpc319 (
      {stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203], stage0_14[204]},
      {stage0_16[102], stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107]},
      {stage1_18[17],stage1_17[51],stage1_16[62],stage1_15[75],stage1_14[87]}
   );
   gpc606_5 gpc320 (
      {stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209], stage0_14[210]},
      {stage0_16[108], stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113]},
      {stage1_18[18],stage1_17[52],stage1_16[63],stage1_15[76],stage1_14[88]}
   );
   gpc606_5 gpc321 (
      {stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215], stage0_14[216]},
      {stage0_16[114], stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119]},
      {stage1_18[19],stage1_17[53],stage1_16[64],stage1_15[77],stage1_14[89]}
   );
   gpc606_5 gpc322 (
      {stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221], stage0_14[222]},
      {stage0_16[120], stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125]},
      {stage1_18[20],stage1_17[54],stage1_16[65],stage1_15[78],stage1_14[90]}
   );
   gpc606_5 gpc323 (
      {stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227], stage0_14[228]},
      {stage0_16[126], stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131]},
      {stage1_18[21],stage1_17[55],stage1_16[66],stage1_15[79],stage1_14[91]}
   );
   gpc606_5 gpc324 (
      {stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233], stage0_14[234]},
      {stage0_16[132], stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137]},
      {stage1_18[22],stage1_17[56],stage1_16[67],stage1_15[80],stage1_14[92]}
   );
   gpc615_5 gpc325 (
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208]},
      {stage0_16[138]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[23],stage1_17[57],stage1_16[68],stage1_15[81]}
   );
   gpc615_5 gpc326 (
      {stage0_15[209], stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213]},
      {stage0_16[139]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[24],stage1_17[58],stage1_16[69],stage1_15[82]}
   );
   gpc615_5 gpc327 (
      {stage0_15[214], stage0_15[215], stage0_15[216], stage0_15[217], stage0_15[218]},
      {stage0_16[140]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[25],stage1_17[59],stage1_16[70],stage1_15[83]}
   );
   gpc615_5 gpc328 (
      {stage0_15[219], stage0_15[220], stage0_15[221], stage0_15[222], stage0_15[223]},
      {stage0_16[141]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[26],stage1_17[60],stage1_16[71],stage1_15[84]}
   );
   gpc615_5 gpc329 (
      {stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227], stage0_15[228]},
      {stage0_16[142]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[27],stage1_17[61],stage1_16[72],stage1_15[85]}
   );
   gpc615_5 gpc330 (
      {stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage0_16[143]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[28],stage1_17[62],stage1_16[73],stage1_15[86]}
   );
   gpc615_5 gpc331 (
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238]},
      {stage0_16[144]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[29],stage1_17[63],stage1_16[74],stage1_15[87]}
   );
   gpc615_5 gpc332 (
      {stage0_15[239], stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243]},
      {stage0_16[145]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[30],stage1_17[64],stage1_16[75],stage1_15[88]}
   );
   gpc615_5 gpc333 (
      {stage0_15[244], stage0_15[245], stage0_15[246], stage0_15[247], stage0_15[248]},
      {stage0_16[146]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[31],stage1_17[65],stage1_16[76],stage1_15[89]}
   );
   gpc615_5 gpc334 (
      {stage0_15[249], stage0_15[250], stage0_15[251], stage0_15[252], stage0_15[253]},
      {stage0_16[147]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[32],stage1_17[66],stage1_16[77],stage1_15[90]}
   );
   gpc606_5 gpc335 (
      {stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151], stage0_16[152], stage0_16[153]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[10],stage1_18[33],stage1_17[67],stage1_16[78]}
   );
   gpc606_5 gpc336 (
      {stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157], stage0_16[158], stage0_16[159]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[11],stage1_18[34],stage1_17[68],stage1_16[79]}
   );
   gpc606_5 gpc337 (
      {stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163], stage0_16[164], stage0_16[165]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[12],stage1_18[35],stage1_17[69],stage1_16[80]}
   );
   gpc606_5 gpc338 (
      {stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169], stage0_16[170], stage0_16[171]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[13],stage1_18[36],stage1_17[70],stage1_16[81]}
   );
   gpc606_5 gpc339 (
      {stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175], stage0_16[176], stage0_16[177]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[14],stage1_18[37],stage1_17[71],stage1_16[82]}
   );
   gpc606_5 gpc340 (
      {stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181], stage0_16[182], stage0_16[183]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[15],stage1_18[38],stage1_17[72],stage1_16[83]}
   );
   gpc606_5 gpc341 (
      {stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188], stage0_16[189]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[16],stage1_18[39],stage1_17[73],stage1_16[84]}
   );
   gpc606_5 gpc342 (
      {stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194], stage0_16[195]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[17],stage1_18[40],stage1_17[74],stage1_16[85]}
   );
   gpc606_5 gpc343 (
      {stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199], stage0_16[200], stage0_16[201]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[18],stage1_18[41],stage1_17[75],stage1_16[86]}
   );
   gpc606_5 gpc344 (
      {stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205], stage0_16[206], stage0_16[207]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[19],stage1_18[42],stage1_17[76],stage1_16[87]}
   );
   gpc606_5 gpc345 (
      {stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211], stage0_16[212], stage0_16[213]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[20],stage1_18[43],stage1_17[77],stage1_16[88]}
   );
   gpc606_5 gpc346 (
      {stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218], stage0_16[219]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[21],stage1_18[44],stage1_17[78],stage1_16[89]}
   );
   gpc606_5 gpc347 (
      {stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224], stage0_16[225]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[22],stage1_18[45],stage1_17[79],stage1_16[90]}
   );
   gpc606_5 gpc348 (
      {stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229], stage0_16[230], stage0_16[231]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[23],stage1_18[46],stage1_17[80],stage1_16[91]}
   );
   gpc606_5 gpc349 (
      {stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235], stage0_16[236], stage0_16[237]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[24],stage1_18[47],stage1_17[81],stage1_16[92]}
   );
   gpc606_5 gpc350 (
      {stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241], stage0_16[242], stage0_16[243]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[25],stage1_18[48],stage1_17[82],stage1_16[93]}
   );
   gpc606_5 gpc351 (
      {stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248], stage0_16[249]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[26],stage1_18[49],stage1_17[83],stage1_16[94]}
   );
   gpc606_5 gpc352 (
      {stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254], stage0_16[255]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[27],stage1_18[50],stage1_17[84],stage1_16[95]}
   );
   gpc606_5 gpc353 (
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[18],stage1_19[28],stage1_18[51],stage1_17[85]}
   );
   gpc606_5 gpc354 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[19],stage1_19[29],stage1_18[52],stage1_17[86]}
   );
   gpc615_5 gpc355 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76]},
      {stage0_18[108]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[20],stage1_19[30],stage1_18[53],stage1_17[87]}
   );
   gpc615_5 gpc356 (
      {stage0_17[77], stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81]},
      {stage0_18[109]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[21],stage1_19[31],stage1_18[54],stage1_17[88]}
   );
   gpc615_5 gpc357 (
      {stage0_17[82], stage0_17[83], stage0_17[84], stage0_17[85], stage0_17[86]},
      {stage0_18[110]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[22],stage1_19[32],stage1_18[55],stage1_17[89]}
   );
   gpc615_5 gpc358 (
      {stage0_17[87], stage0_17[88], stage0_17[89], stage0_17[90], stage0_17[91]},
      {stage0_18[111]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[23],stage1_19[33],stage1_18[56],stage1_17[90]}
   );
   gpc615_5 gpc359 (
      {stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95], stage0_17[96]},
      {stage0_18[112]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[24],stage1_19[34],stage1_18[57],stage1_17[91]}
   );
   gpc615_5 gpc360 (
      {stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_18[113]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[25],stage1_19[35],stage1_18[58],stage1_17[92]}
   );
   gpc615_5 gpc361 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106]},
      {stage0_18[114]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[26],stage1_19[36],stage1_18[59],stage1_17[93]}
   );
   gpc615_5 gpc362 (
      {stage0_17[107], stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111]},
      {stage0_18[115]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[27],stage1_19[37],stage1_18[60],stage1_17[94]}
   );
   gpc615_5 gpc363 (
      {stage0_17[112], stage0_17[113], stage0_17[114], stage0_17[115], stage0_17[116]},
      {stage0_18[116]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[28],stage1_19[38],stage1_18[61],stage1_17[95]}
   );
   gpc615_5 gpc364 (
      {stage0_17[117], stage0_17[118], stage0_17[119], stage0_17[120], stage0_17[121]},
      {stage0_18[117]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[29],stage1_19[39],stage1_18[62],stage1_17[96]}
   );
   gpc615_5 gpc365 (
      {stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125], stage0_17[126]},
      {stage0_18[118]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[30],stage1_19[40],stage1_18[63],stage1_17[97]}
   );
   gpc615_5 gpc366 (
      {stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage0_18[119]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[31],stage1_19[41],stage1_18[64],stage1_17[98]}
   );
   gpc615_5 gpc367 (
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136]},
      {stage0_18[120]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[32],stage1_19[42],stage1_18[65],stage1_17[99]}
   );
   gpc615_5 gpc368 (
      {stage0_17[137], stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141]},
      {stage0_18[121]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[33],stage1_19[43],stage1_18[66],stage1_17[100]}
   );
   gpc615_5 gpc369 (
      {stage0_17[142], stage0_17[143], stage0_17[144], stage0_17[145], stage0_17[146]},
      {stage0_18[122]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[34],stage1_19[44],stage1_18[67],stage1_17[101]}
   );
   gpc615_5 gpc370 (
      {stage0_17[147], stage0_17[148], stage0_17[149], stage0_17[150], stage0_17[151]},
      {stage0_18[123]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[35],stage1_19[45],stage1_18[68],stage1_17[102]}
   );
   gpc615_5 gpc371 (
      {stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155], stage0_17[156]},
      {stage0_18[124]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[36],stage1_19[46],stage1_18[69],stage1_17[103]}
   );
   gpc615_5 gpc372 (
      {stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_18[125]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[37],stage1_19[47],stage1_18[70],stage1_17[104]}
   );
   gpc615_5 gpc373 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166]},
      {stage0_18[126]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[38],stage1_19[48],stage1_18[71],stage1_17[105]}
   );
   gpc615_5 gpc374 (
      {stage0_17[167], stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171]},
      {stage0_18[127]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[39],stage1_19[49],stage1_18[72],stage1_17[106]}
   );
   gpc615_5 gpc375 (
      {stage0_17[172], stage0_17[173], stage0_17[174], stage0_17[175], stage0_17[176]},
      {stage0_18[128]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[40],stage1_19[50],stage1_18[73],stage1_17[107]}
   );
   gpc615_5 gpc376 (
      {stage0_17[177], stage0_17[178], stage0_17[179], stage0_17[180], stage0_17[181]},
      {stage0_18[129]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[41],stage1_19[51],stage1_18[74],stage1_17[108]}
   );
   gpc615_5 gpc377 (
      {stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185], stage0_17[186]},
      {stage0_18[130]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[42],stage1_19[52],stage1_18[75],stage1_17[109]}
   );
   gpc615_5 gpc378 (
      {stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_18[131]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[43],stage1_19[53],stage1_18[76],stage1_17[110]}
   );
   gpc615_5 gpc379 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196]},
      {stage0_18[132]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[44],stage1_19[54],stage1_18[77],stage1_17[111]}
   );
   gpc615_5 gpc380 (
      {stage0_17[197], stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201]},
      {stage0_18[133]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[45],stage1_19[55],stage1_18[78],stage1_17[112]}
   );
   gpc615_5 gpc381 (
      {stage0_17[202], stage0_17[203], stage0_17[204], stage0_17[205], stage0_17[206]},
      {stage0_18[134]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[46],stage1_19[56],stage1_18[79],stage1_17[113]}
   );
   gpc615_5 gpc382 (
      {stage0_17[207], stage0_17[208], stage0_17[209], stage0_17[210], stage0_17[211]},
      {stage0_18[135]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[47],stage1_19[57],stage1_18[80],stage1_17[114]}
   );
   gpc615_5 gpc383 (
      {stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215], stage0_17[216]},
      {stage0_18[136]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[48],stage1_19[58],stage1_18[81],stage1_17[115]}
   );
   gpc615_5 gpc384 (
      {stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_18[137]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[49],stage1_19[59],stage1_18[82],stage1_17[116]}
   );
   gpc615_5 gpc385 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226]},
      {stage0_18[138]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[50],stage1_19[60],stage1_18[83],stage1_17[117]}
   );
   gpc615_5 gpc386 (
      {stage0_17[227], stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231]},
      {stage0_18[139]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[51],stage1_19[61],stage1_18[84],stage1_17[118]}
   );
   gpc615_5 gpc387 (
      {stage0_17[232], stage0_17[233], stage0_17[234], stage0_17[235], stage0_17[236]},
      {stage0_18[140]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[52],stage1_19[62],stage1_18[85],stage1_17[119]}
   );
   gpc615_5 gpc388 (
      {stage0_17[237], stage0_17[238], stage0_17[239], stage0_17[240], stage0_17[241]},
      {stage0_18[141]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[53],stage1_19[63],stage1_18[86],stage1_17[120]}
   );
   gpc615_5 gpc389 (
      {stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245], stage0_17[246]},
      {stage0_18[142]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[54],stage1_19[64],stage1_18[87],stage1_17[121]}
   );
   gpc615_5 gpc390 (
      {stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_18[143]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[55],stage1_19[65],stage1_18[88],stage1_17[122]}
   );
   gpc606_5 gpc391 (
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[38],stage1_20[56],stage1_19[66],stage1_18[89]}
   );
   gpc606_5 gpc392 (
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[39],stage1_20[57],stage1_19[67],stage1_18[90]}
   );
   gpc606_5 gpc393 (
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[40],stage1_20[58],stage1_19[68],stage1_18[91]}
   );
   gpc606_5 gpc394 (
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[41],stage1_20[59],stage1_19[69],stage1_18[92]}
   );
   gpc606_5 gpc395 (
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[42],stage1_20[60],stage1_19[70],stage1_18[93]}
   );
   gpc606_5 gpc396 (
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[43],stage1_20[61],stage1_19[71],stage1_18[94]}
   );
   gpc606_5 gpc397 (
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[44],stage1_20[62],stage1_19[72],stage1_18[95]}
   );
   gpc606_5 gpc398 (
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[45],stage1_20[63],stage1_19[73],stage1_18[96]}
   );
   gpc606_5 gpc399 (
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[46],stage1_20[64],stage1_19[74],stage1_18[97]}
   );
   gpc606_5 gpc400 (
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[47],stage1_20[65],stage1_19[75],stage1_18[98]}
   );
   gpc606_5 gpc401 (
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[10],stage1_21[48],stage1_20[66],stage1_19[76]}
   );
   gpc606_5 gpc402 (
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[11],stage1_21[49],stage1_20[67],stage1_19[77]}
   );
   gpc615_5 gpc403 (
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64]},
      {stage0_21[12]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[12],stage1_21[50],stage1_20[68]}
   );
   gpc615_5 gpc404 (
      {stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69]},
      {stage0_21[13]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[13],stage1_21[51],stage1_20[69]}
   );
   gpc615_5 gpc405 (
      {stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74]},
      {stage0_21[14]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[14],stage1_21[52],stage1_20[70]}
   );
   gpc615_5 gpc406 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79]},
      {stage0_21[15]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[15],stage1_21[53],stage1_20[71]}
   );
   gpc615_5 gpc407 (
      {stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84]},
      {stage0_21[16]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[16],stage1_21[54],stage1_20[72]}
   );
   gpc615_5 gpc408 (
      {stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage0_21[17]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[17],stage1_21[55],stage1_20[73]}
   );
   gpc615_5 gpc409 (
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94]},
      {stage0_21[18]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[18],stage1_21[56],stage1_20[74]}
   );
   gpc615_5 gpc410 (
      {stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99]},
      {stage0_21[19]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[9],stage1_22[19],stage1_21[57],stage1_20[75]}
   );
   gpc615_5 gpc411 (
      {stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_21[20]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[10],stage1_22[20],stage1_21[58],stage1_20[76]}
   );
   gpc615_5 gpc412 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109]},
      {stage0_21[21]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[11],stage1_22[21],stage1_21[59],stage1_20[77]}
   );
   gpc615_5 gpc413 (
      {stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114]},
      {stage0_21[22]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[12],stage1_22[22],stage1_21[60],stage1_20[78]}
   );
   gpc615_5 gpc414 (
      {stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage0_21[23]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[13],stage1_22[23],stage1_21[61],stage1_20[79]}
   );
   gpc615_5 gpc415 (
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124]},
      {stage0_21[24]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[14],stage1_22[24],stage1_21[62],stage1_20[80]}
   );
   gpc615_5 gpc416 (
      {stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129]},
      {stage0_21[25]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[15],stage1_22[25],stage1_21[63],stage1_20[81]}
   );
   gpc615_5 gpc417 (
      {stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134]},
      {stage0_21[26]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[16],stage1_22[26],stage1_21[64],stage1_20[82]}
   );
   gpc615_5 gpc418 (
      {stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139]},
      {stage0_21[27]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[17],stage1_22[27],stage1_21[65],stage1_20[83]}
   );
   gpc615_5 gpc419 (
      {stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144]},
      {stage0_21[28]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[18],stage1_22[28],stage1_21[66],stage1_20[84]}
   );
   gpc615_5 gpc420 (
      {stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage0_21[29]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[19],stage1_22[29],stage1_21[67],stage1_20[85]}
   );
   gpc615_5 gpc421 (
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154]},
      {stage0_21[30]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[20],stage1_22[30],stage1_21[68],stage1_20[86]}
   );
   gpc615_5 gpc422 (
      {stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159]},
      {stage0_21[31]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[21],stage1_22[31],stage1_21[69],stage1_20[87]}
   );
   gpc615_5 gpc423 (
      {stage0_20[160], stage0_20[161], stage0_20[162], stage0_20[163], stage0_20[164]},
      {stage0_21[32]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[22],stage1_22[32],stage1_21[70],stage1_20[88]}
   );
   gpc615_5 gpc424 (
      {stage0_20[165], stage0_20[166], stage0_20[167], stage0_20[168], stage0_20[169]},
      {stage0_21[33]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[23],stage1_22[33],stage1_21[71],stage1_20[89]}
   );
   gpc615_5 gpc425 (
      {stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173], stage0_20[174]},
      {stage0_21[34]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[24],stage1_22[34],stage1_21[72],stage1_20[90]}
   );
   gpc615_5 gpc426 (
      {stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage0_21[35]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[25],stage1_22[35],stage1_21[73],stage1_20[91]}
   );
   gpc615_5 gpc427 (
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184]},
      {stage0_21[36]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[26],stage1_22[36],stage1_21[74],stage1_20[92]}
   );
   gpc615_5 gpc428 (
      {stage0_20[185], stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189]},
      {stage0_21[37]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[27],stage1_22[37],stage1_21[75],stage1_20[93]}
   );
   gpc615_5 gpc429 (
      {stage0_20[190], stage0_20[191], stage0_20[192], stage0_20[193], stage0_20[194]},
      {stage0_21[38]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[28],stage1_22[38],stage1_21[76],stage1_20[94]}
   );
   gpc615_5 gpc430 (
      {stage0_20[195], stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199]},
      {stage0_21[39]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[29],stage1_22[39],stage1_21[77],stage1_20[95]}
   );
   gpc615_5 gpc431 (
      {stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203], stage0_20[204]},
      {stage0_21[40]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[30],stage1_22[40],stage1_21[78],stage1_20[96]}
   );
   gpc615_5 gpc432 (
      {stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage0_21[41]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[31],stage1_22[41],stage1_21[79],stage1_20[97]}
   );
   gpc615_5 gpc433 (
      {stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214]},
      {stage0_21[42]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[32],stage1_22[42],stage1_21[80],stage1_20[98]}
   );
   gpc615_5 gpc434 (
      {stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219]},
      {stage0_21[43]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[33],stage1_22[43],stage1_21[81],stage1_20[99]}
   );
   gpc615_5 gpc435 (
      {stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224]},
      {stage0_21[44]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[34],stage1_22[44],stage1_21[82],stage1_20[100]}
   );
   gpc615_5 gpc436 (
      {stage0_20[225], stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229]},
      {stage0_21[45]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[35],stage1_22[45],stage1_21[83],stage1_20[101]}
   );
   gpc615_5 gpc437 (
      {stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233], stage0_20[234]},
      {stage0_21[46]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[36],stage1_22[46],stage1_21[84],stage1_20[102]}
   );
   gpc615_5 gpc438 (
      {stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_21[47]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[37],stage1_22[47],stage1_21[85],stage1_20[103]}
   );
   gpc615_5 gpc439 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244]},
      {stage0_21[48]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[38],stage1_22[48],stage1_21[86],stage1_20[104]}
   );
   gpc606_5 gpc440 (
      {stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[37],stage1_23[39],stage1_22[49],stage1_21[87]}
   );
   gpc606_5 gpc441 (
      {stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59], stage0_21[60]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[38],stage1_23[40],stage1_22[50],stage1_21[88]}
   );
   gpc606_5 gpc442 (
      {stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65], stage0_21[66]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[39],stage1_23[41],stage1_22[51],stage1_21[89]}
   );
   gpc606_5 gpc443 (
      {stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[40],stage1_23[42],stage1_22[52],stage1_21[90]}
   );
   gpc606_5 gpc444 (
      {stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[41],stage1_23[43],stage1_22[53],stage1_21[91]}
   );
   gpc606_5 gpc445 (
      {stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[42],stage1_23[44],stage1_22[54],stage1_21[92]}
   );
   gpc606_5 gpc446 (
      {stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[43],stage1_23[45],stage1_22[55],stage1_21[93]}
   );
   gpc606_5 gpc447 (
      {stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95], stage0_21[96]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[44],stage1_23[46],stage1_22[56],stage1_21[94]}
   );
   gpc606_5 gpc448 (
      {stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101], stage0_21[102]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[45],stage1_23[47],stage1_22[57],stage1_21[95]}
   );
   gpc606_5 gpc449 (
      {stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107], stage0_21[108]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[46],stage1_23[48],stage1_22[58],stage1_21[96]}
   );
   gpc606_5 gpc450 (
      {stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[47],stage1_23[49],stage1_22[59],stage1_21[97]}
   );
   gpc606_5 gpc451 (
      {stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[48],stage1_23[50],stage1_22[60],stage1_21[98]}
   );
   gpc606_5 gpc452 (
      {stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125], stage0_21[126]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[49],stage1_23[51],stage1_22[61],stage1_21[99]}
   );
   gpc606_5 gpc453 (
      {stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131], stage0_21[132]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[50],stage1_23[52],stage1_22[62],stage1_21[100]}
   );
   gpc606_5 gpc454 (
      {stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137], stage0_21[138]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[51],stage1_23[53],stage1_22[63],stage1_21[101]}
   );
   gpc606_5 gpc455 (
      {stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143], stage0_21[144]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[52],stage1_23[54],stage1_22[64],stage1_21[102]}
   );
   gpc606_5 gpc456 (
      {stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149], stage0_21[150]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[53],stage1_23[55],stage1_22[65],stage1_21[103]}
   );
   gpc606_5 gpc457 (
      {stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155], stage0_21[156]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[54],stage1_23[56],stage1_22[66],stage1_21[104]}
   );
   gpc606_5 gpc458 (
      {stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161], stage0_21[162]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[55],stage1_23[57],stage1_22[67],stage1_21[105]}
   );
   gpc606_5 gpc459 (
      {stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167], stage0_21[168]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[56],stage1_23[58],stage1_22[68],stage1_21[106]}
   );
   gpc606_5 gpc460 (
      {stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173], stage0_21[174]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[57],stage1_23[59],stage1_22[69],stage1_21[107]}
   );
   gpc606_5 gpc461 (
      {stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179], stage0_21[180]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[58],stage1_23[60],stage1_22[70],stage1_21[108]}
   );
   gpc606_5 gpc462 (
      {stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185], stage0_21[186]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[59],stage1_23[61],stage1_22[71],stage1_21[109]}
   );
   gpc606_5 gpc463 (
      {stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191], stage0_21[192]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[60],stage1_23[62],stage1_22[72],stage1_21[110]}
   );
   gpc606_5 gpc464 (
      {stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197], stage0_21[198]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[61],stage1_23[63],stage1_22[73],stage1_21[111]}
   );
   gpc606_5 gpc465 (
      {stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203], stage0_21[204]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[62],stage1_23[64],stage1_22[74],stage1_21[112]}
   );
   gpc606_5 gpc466 (
      {stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209], stage0_21[210]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[63],stage1_23[65],stage1_22[75],stage1_21[113]}
   );
   gpc606_5 gpc467 (
      {stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215], stage0_21[216]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[64],stage1_23[66],stage1_22[76],stage1_21[114]}
   );
   gpc606_5 gpc468 (
      {stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221], stage0_21[222]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[65],stage1_23[67],stage1_22[77],stage1_21[115]}
   );
   gpc606_5 gpc469 (
      {stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227], stage0_21[228]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[66],stage1_23[68],stage1_22[78],stage1_21[116]}
   );
   gpc606_5 gpc470 (
      {stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233], stage0_21[234]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[67],stage1_23[69],stage1_22[79],stage1_21[117]}
   );
   gpc606_5 gpc471 (
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[31],stage1_24[68],stage1_23[70],stage1_22[80]}
   );
   gpc606_5 gpc472 (
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[32],stage1_24[69],stage1_23[71],stage1_22[81]}
   );
   gpc606_5 gpc473 (
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[33],stage1_24[70],stage1_23[72],stage1_22[82]}
   );
   gpc606_5 gpc474 (
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[34],stage1_24[71],stage1_23[73],stage1_22[83]}
   );
   gpc606_5 gpc475 (
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[4],stage1_25[35],stage1_24[72],stage1_23[74]}
   );
   gpc606_5 gpc476 (
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[5],stage1_25[36],stage1_24[73],stage1_23[75]}
   );
   gpc606_5 gpc477 (
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[6],stage1_25[37],stage1_24[74],stage1_23[76]}
   );
   gpc606_5 gpc478 (
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[7],stage1_25[38],stage1_24[75],stage1_23[77]}
   );
   gpc606_5 gpc479 (
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[8],stage1_25[39],stage1_24[76],stage1_23[78]}
   );
   gpc606_5 gpc480 (
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[9],stage1_25[40],stage1_24[77],stage1_23[79]}
   );
   gpc606_5 gpc481 (
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[10],stage1_25[41],stage1_24[78],stage1_23[80]}
   );
   gpc606_5 gpc482 (
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[11],stage1_25[42],stage1_24[79],stage1_23[81]}
   );
   gpc606_5 gpc483 (
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[12],stage1_25[43],stage1_24[80],stage1_23[82]}
   );
   gpc606_5 gpc484 (
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[13],stage1_25[44],stage1_24[81],stage1_23[83]}
   );
   gpc606_5 gpc485 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[14],stage1_25[45],stage1_24[82]}
   );
   gpc606_5 gpc486 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[15],stage1_25[46],stage1_24[83]}
   );
   gpc606_5 gpc487 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[16],stage1_25[47],stage1_24[84]}
   );
   gpc606_5 gpc488 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[17],stage1_25[48],stage1_24[85]}
   );
   gpc606_5 gpc489 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[18],stage1_25[49],stage1_24[86]}
   );
   gpc606_5 gpc490 (
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[19],stage1_25[50],stage1_24[87]}
   );
   gpc606_5 gpc491 (
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[16],stage1_26[20],stage1_25[51],stage1_24[88]}
   );
   gpc606_5 gpc492 (
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[17],stage1_26[21],stage1_25[52],stage1_24[89]}
   );
   gpc606_5 gpc493 (
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[18],stage1_26[22],stage1_25[53],stage1_24[90]}
   );
   gpc606_5 gpc494 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[19],stage1_26[23],stage1_25[54],stage1_24[91]}
   );
   gpc606_5 gpc495 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[20],stage1_26[24],stage1_25[55],stage1_24[92]}
   );
   gpc606_5 gpc496 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[21],stage1_26[25],stage1_25[56],stage1_24[93]}
   );
   gpc606_5 gpc497 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[12],stage1_27[22],stage1_26[26],stage1_25[57]}
   );
   gpc606_5 gpc498 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[13],stage1_27[23],stage1_26[27],stage1_25[58]}
   );
   gpc606_5 gpc499 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[14],stage1_27[24],stage1_26[28],stage1_25[59]}
   );
   gpc606_5 gpc500 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[15],stage1_27[25],stage1_26[29],stage1_25[60]}
   );
   gpc606_5 gpc501 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[16],stage1_27[26],stage1_26[30],stage1_25[61]}
   );
   gpc606_5 gpc502 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[17],stage1_27[27],stage1_26[31],stage1_25[62]}
   );
   gpc606_5 gpc503 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[18],stage1_27[28],stage1_26[32],stage1_25[63]}
   );
   gpc606_5 gpc504 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[19],stage1_27[29],stage1_26[33],stage1_25[64]}
   );
   gpc606_5 gpc505 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[20],stage1_27[30],stage1_26[34],stage1_25[65]}
   );
   gpc606_5 gpc506 (
      {stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[21],stage1_27[31],stage1_26[35],stage1_25[66]}
   );
   gpc606_5 gpc507 (
      {stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[22],stage1_27[32],stage1_26[36],stage1_25[67]}
   );
   gpc606_5 gpc508 (
      {stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[23],stage1_27[33],stage1_26[37],stage1_25[68]}
   );
   gpc606_5 gpc509 (
      {stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[24],stage1_27[34],stage1_26[38],stage1_25[69]}
   );
   gpc606_5 gpc510 (
      {stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[25],stage1_27[35],stage1_26[39],stage1_25[70]}
   );
   gpc606_5 gpc511 (
      {stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[26],stage1_27[36],stage1_26[40],stage1_25[71]}
   );
   gpc606_5 gpc512 (
      {stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[27],stage1_27[37],stage1_26[41],stage1_25[72]}
   );
   gpc606_5 gpc513 (
      {stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[28],stage1_27[38],stage1_26[42],stage1_25[73]}
   );
   gpc606_5 gpc514 (
      {stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[29],stage1_27[39],stage1_26[43],stage1_25[74]}
   );
   gpc606_5 gpc515 (
      {stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[30],stage1_27[40],stage1_26[44],stage1_25[75]}
   );
   gpc606_5 gpc516 (
      {stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[31],stage1_27[41],stage1_26[45],stage1_25[76]}
   );
   gpc606_5 gpc517 (
      {stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[32],stage1_27[42],stage1_26[46],stage1_25[77]}
   );
   gpc606_5 gpc518 (
      {stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[33],stage1_27[43],stage1_26[47],stage1_25[78]}
   );
   gpc606_5 gpc519 (
      {stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[34],stage1_27[44],stage1_26[48],stage1_25[79]}
   );
   gpc606_5 gpc520 (
      {stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[35],stage1_27[45],stage1_26[49],stage1_25[80]}
   );
   gpc606_5 gpc521 (
      {stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[36],stage1_27[46],stage1_26[50],stage1_25[81]}
   );
   gpc606_5 gpc522 (
      {stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[37],stage1_27[47],stage1_26[51],stage1_25[82]}
   );
   gpc606_5 gpc523 (
      {stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[38],stage1_27[48],stage1_26[52],stage1_25[83]}
   );
   gpc606_5 gpc524 (
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[27],stage1_28[39],stage1_27[49]}
   );
   gpc606_5 gpc525 (
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[1],stage1_29[28],stage1_28[40],stage1_27[50]}
   );
   gpc606_5 gpc526 (
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[2],stage1_29[29],stage1_28[41],stage1_27[51]}
   );
   gpc606_5 gpc527 (
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[3],stage1_29[30],stage1_28[42],stage1_27[52]}
   );
   gpc606_5 gpc528 (
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[4],stage1_29[31],stage1_28[43],stage1_27[53]}
   );
   gpc606_5 gpc529 (
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[5],stage1_29[32],stage1_28[44],stage1_27[54]}
   );
   gpc606_5 gpc530 (
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[6],stage1_29[33],stage1_28[45],stage1_27[55]}
   );
   gpc606_5 gpc531 (
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[7],stage1_30[7],stage1_29[34],stage1_28[46]}
   );
   gpc606_5 gpc532 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[8],stage1_30[8],stage1_29[35],stage1_28[47]}
   );
   gpc606_5 gpc533 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[9],stage1_30[9],stage1_29[36],stage1_28[48]}
   );
   gpc606_5 gpc534 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[10],stage1_30[10],stage1_29[37],stage1_28[49]}
   );
   gpc606_5 gpc535 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[11],stage1_30[11],stage1_29[38],stage1_28[50]}
   );
   gpc606_5 gpc536 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[12],stage1_30[12],stage1_29[39],stage1_28[51]}
   );
   gpc606_5 gpc537 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[13],stage1_30[13],stage1_29[40],stage1_28[52]}
   );
   gpc606_5 gpc538 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[14],stage1_30[14],stage1_29[41],stage1_28[53]}
   );
   gpc606_5 gpc539 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[15],stage1_30[15],stage1_29[42],stage1_28[54]}
   );
   gpc606_5 gpc540 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[16],stage1_30[16],stage1_29[43],stage1_28[55]}
   );
   gpc606_5 gpc541 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[17],stage1_30[17],stage1_29[44],stage1_28[56]}
   );
   gpc606_5 gpc542 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[18],stage1_30[18],stage1_29[45],stage1_28[57]}
   );
   gpc606_5 gpc543 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[19],stage1_30[19],stage1_29[46],stage1_28[58]}
   );
   gpc606_5 gpc544 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[20],stage1_30[20],stage1_29[47],stage1_28[59]}
   );
   gpc606_5 gpc545 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[21],stage1_30[21],stage1_29[48],stage1_28[60]}
   );
   gpc606_5 gpc546 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[22],stage1_30[22],stage1_29[49],stage1_28[61]}
   );
   gpc606_5 gpc547 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[23],stage1_30[23],stage1_29[50],stage1_28[62]}
   );
   gpc606_5 gpc548 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[24],stage1_30[24],stage1_29[51],stage1_28[63]}
   );
   gpc606_5 gpc549 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[25],stage1_30[25],stage1_29[52],stage1_28[64]}
   );
   gpc606_5 gpc550 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[26],stage1_30[26],stage1_29[53],stage1_28[65]}
   );
   gpc606_5 gpc551 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[27],stage1_30[27],stage1_29[54],stage1_28[66]}
   );
   gpc606_5 gpc552 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[28],stage1_30[28],stage1_29[55],stage1_28[67]}
   );
   gpc606_5 gpc553 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[29],stage1_30[29],stage1_29[56],stage1_28[68]}
   );
   gpc606_5 gpc554 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[30],stage1_30[30],stage1_29[57],stage1_28[69]}
   );
   gpc606_5 gpc555 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[31],stage1_30[31],stage1_29[58],stage1_28[70]}
   );
   gpc606_5 gpc556 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[32],stage1_30[32],stage1_29[59],stage1_28[71]}
   );
   gpc606_5 gpc557 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[33],stage1_30[33],stage1_29[60],stage1_28[72]}
   );
   gpc606_5 gpc558 (
      {stage0_28[162], stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[34],stage1_30[34],stage1_29[61],stage1_28[73]}
   );
   gpc606_5 gpc559 (
      {stage0_28[168], stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[35],stage1_30[35],stage1_29[62],stage1_28[74]}
   );
   gpc606_5 gpc560 (
      {stage0_28[174], stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[36],stage1_30[36],stage1_29[63],stage1_28[75]}
   );
   gpc606_5 gpc561 (
      {stage0_28[180], stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[37],stage1_30[37],stage1_29[64],stage1_28[76]}
   );
   gpc606_5 gpc562 (
      {stage0_28[186], stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[38],stage1_30[38],stage1_29[65],stage1_28[77]}
   );
   gpc606_5 gpc563 (
      {stage0_28[192], stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[39],stage1_30[39],stage1_29[66],stage1_28[78]}
   );
   gpc606_5 gpc564 (
      {stage0_28[198], stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[40],stage1_30[40],stage1_29[67],stage1_28[79]}
   );
   gpc606_5 gpc565 (
      {stage0_28[204], stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[41],stage1_30[41],stage1_29[68],stage1_28[80]}
   );
   gpc606_5 gpc566 (
      {stage0_28[210], stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[42],stage1_30[42],stage1_29[69],stage1_28[81]}
   );
   gpc606_5 gpc567 (
      {stage0_28[216], stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[43],stage1_30[43],stage1_29[70],stage1_28[82]}
   );
   gpc606_5 gpc568 (
      {stage0_28[222], stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[44],stage1_30[44],stage1_29[71],stage1_28[83]}
   );
   gpc606_5 gpc569 (
      {stage0_28[228], stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[45],stage1_30[45],stage1_29[72],stage1_28[84]}
   );
   gpc606_5 gpc570 (
      {stage0_28[234], stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[46],stage1_30[46],stage1_29[73],stage1_28[85]}
   );
   gpc606_5 gpc571 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[40],stage1_31[47],stage1_30[47],stage1_29[74]}
   );
   gpc606_5 gpc572 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[41],stage1_31[48],stage1_30[48],stage1_29[75]}
   );
   gpc606_5 gpc573 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[42],stage1_31[49],stage1_30[49],stage1_29[76]}
   );
   gpc606_5 gpc574 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[43],stage1_31[50],stage1_30[50],stage1_29[77]}
   );
   gpc606_5 gpc575 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[44],stage1_31[51],stage1_30[51],stage1_29[78]}
   );
   gpc606_5 gpc576 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[45],stage1_31[52],stage1_30[52],stage1_29[79]}
   );
   gpc606_5 gpc577 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[46],stage1_31[53],stage1_30[53],stage1_29[80]}
   );
   gpc606_5 gpc578 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[47],stage1_31[54],stage1_30[54],stage1_29[81]}
   );
   gpc606_5 gpc579 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[48],stage1_31[55],stage1_30[55],stage1_29[82]}
   );
   gpc606_5 gpc580 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[49],stage1_31[56],stage1_30[56],stage1_29[83]}
   );
   gpc606_5 gpc581 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[50],stage1_31[57],stage1_30[57],stage1_29[84]}
   );
   gpc606_5 gpc582 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[51],stage1_31[58],stage1_30[58],stage1_29[85]}
   );
   gpc606_5 gpc583 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[52],stage1_31[59],stage1_30[59],stage1_29[86]}
   );
   gpc606_5 gpc584 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[53],stage1_31[60],stage1_30[60],stage1_29[87]}
   );
   gpc606_5 gpc585 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[54],stage1_31[61],stage1_30[61],stage1_29[88]}
   );
   gpc606_5 gpc586 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[55],stage1_31[62],stage1_30[62],stage1_29[89]}
   );
   gpc606_5 gpc587 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[56],stage1_31[63],stage1_30[63],stage1_29[90]}
   );
   gpc606_5 gpc588 (
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[57],stage1_31[64],stage1_30[64],stage1_29[91]}
   );
   gpc606_5 gpc589 (
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[58],stage1_31[65],stage1_30[65],stage1_29[92]}
   );
   gpc606_5 gpc590 (
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[59],stage1_31[66],stage1_30[66],stage1_29[93]}
   );
   gpc606_5 gpc591 (
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[60],stage1_31[67],stage1_30[67],stage1_29[94]}
   );
   gpc606_5 gpc592 (
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[61],stage1_31[68],stage1_30[68],stage1_29[95]}
   );
   gpc606_5 gpc593 (
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[62],stage1_31[69],stage1_30[69],stage1_29[96]}
   );
   gpc606_5 gpc594 (
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[63],stage1_31[70],stage1_30[70],stage1_29[97]}
   );
   gpc606_5 gpc595 (
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[64],stage1_31[71],stage1_30[71],stage1_29[98]}
   );
   gpc606_5 gpc596 (
      {stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[65],stage1_31[72],stage1_30[72],stage1_29[99]}
   );
   gpc606_5 gpc597 (
      {stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[66],stage1_31[73],stage1_30[73],stage1_29[100]}
   );
   gpc606_5 gpc598 (
      {stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[67],stage1_31[74],stage1_30[74],stage1_29[101]}
   );
   gpc606_5 gpc599 (
      {stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[68],stage1_31[75],stage1_30[75],stage1_29[102]}
   );
   gpc606_5 gpc600 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[69],stage1_31[76],stage1_30[76],stage1_29[103]}
   );
   gpc606_5 gpc601 (
      {stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[70],stage1_31[77],stage1_30[77],stage1_29[104]}
   );
   gpc606_5 gpc602 (
      {stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[71],stage1_31[78],stage1_30[78],stage1_29[105]}
   );
   gpc606_5 gpc603 (
      {stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[72],stage1_31[79],stage1_30[79],stage1_29[106]}
   );
   gpc606_5 gpc604 (
      {stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[73],stage1_31[80],stage1_30[80],stage1_29[107]}
   );
   gpc1_1 gpc605 (
      {stage0_0[249]},
      {stage1_0[43]}
   );
   gpc1_1 gpc606 (
      {stage0_0[250]},
      {stage1_0[44]}
   );
   gpc1_1 gpc607 (
      {stage0_0[251]},
      {stage1_0[45]}
   );
   gpc1_1 gpc608 (
      {stage0_0[252]},
      {stage1_0[46]}
   );
   gpc1_1 gpc609 (
      {stage0_0[253]},
      {stage1_0[47]}
   );
   gpc1_1 gpc610 (
      {stage0_0[254]},
      {stage1_0[48]}
   );
   gpc1_1 gpc611 (
      {stage0_0[255]},
      {stage1_0[49]}
   );
   gpc1_1 gpc612 (
      {stage0_1[237]},
      {stage1_1[79]}
   );
   gpc1_1 gpc613 (
      {stage0_1[238]},
      {stage1_1[80]}
   );
   gpc1_1 gpc614 (
      {stage0_1[239]},
      {stage1_1[81]}
   );
   gpc1_1 gpc615 (
      {stage0_1[240]},
      {stage1_1[82]}
   );
   gpc1_1 gpc616 (
      {stage0_1[241]},
      {stage1_1[83]}
   );
   gpc1_1 gpc617 (
      {stage0_1[242]},
      {stage1_1[84]}
   );
   gpc1_1 gpc618 (
      {stage0_1[243]},
      {stage1_1[85]}
   );
   gpc1_1 gpc619 (
      {stage0_1[244]},
      {stage1_1[86]}
   );
   gpc1_1 gpc620 (
      {stage0_1[245]},
      {stage1_1[87]}
   );
   gpc1_1 gpc621 (
      {stage0_1[246]},
      {stage1_1[88]}
   );
   gpc1_1 gpc622 (
      {stage0_1[247]},
      {stage1_1[89]}
   );
   gpc1_1 gpc623 (
      {stage0_1[248]},
      {stage1_1[90]}
   );
   gpc1_1 gpc624 (
      {stage0_1[249]},
      {stage1_1[91]}
   );
   gpc1_1 gpc625 (
      {stage0_1[250]},
      {stage1_1[92]}
   );
   gpc1_1 gpc626 (
      {stage0_1[251]},
      {stage1_1[93]}
   );
   gpc1_1 gpc627 (
      {stage0_1[252]},
      {stage1_1[94]}
   );
   gpc1_1 gpc628 (
      {stage0_1[253]},
      {stage1_1[95]}
   );
   gpc1_1 gpc629 (
      {stage0_1[254]},
      {stage1_1[96]}
   );
   gpc1_1 gpc630 (
      {stage0_1[255]},
      {stage1_1[97]}
   );
   gpc1_1 gpc631 (
      {stage0_2[246]},
      {stage1_2[82]}
   );
   gpc1_1 gpc632 (
      {stage0_2[247]},
      {stage1_2[83]}
   );
   gpc1_1 gpc633 (
      {stage0_2[248]},
      {stage1_2[84]}
   );
   gpc1_1 gpc634 (
      {stage0_2[249]},
      {stage1_2[85]}
   );
   gpc1_1 gpc635 (
      {stage0_2[250]},
      {stage1_2[86]}
   );
   gpc1_1 gpc636 (
      {stage0_2[251]},
      {stage1_2[87]}
   );
   gpc1_1 gpc637 (
      {stage0_2[252]},
      {stage1_2[88]}
   );
   gpc1_1 gpc638 (
      {stage0_2[253]},
      {stage1_2[89]}
   );
   gpc1_1 gpc639 (
      {stage0_2[254]},
      {stage1_2[90]}
   );
   gpc1_1 gpc640 (
      {stage0_2[255]},
      {stage1_2[91]}
   );
   gpc1_1 gpc641 (
      {stage0_3[254]},
      {stage1_3[89]}
   );
   gpc1_1 gpc642 (
      {stage0_3[255]},
      {stage1_3[90]}
   );
   gpc1_1 gpc643 (
      {stage0_4[230]},
      {stage1_4[123]}
   );
   gpc1_1 gpc644 (
      {stage0_4[231]},
      {stage1_4[124]}
   );
   gpc1_1 gpc645 (
      {stage0_4[232]},
      {stage1_4[125]}
   );
   gpc1_1 gpc646 (
      {stage0_4[233]},
      {stage1_4[126]}
   );
   gpc1_1 gpc647 (
      {stage0_4[234]},
      {stage1_4[127]}
   );
   gpc1_1 gpc648 (
      {stage0_4[235]},
      {stage1_4[128]}
   );
   gpc1_1 gpc649 (
      {stage0_4[236]},
      {stage1_4[129]}
   );
   gpc1_1 gpc650 (
      {stage0_4[237]},
      {stage1_4[130]}
   );
   gpc1_1 gpc651 (
      {stage0_4[238]},
      {stage1_4[131]}
   );
   gpc1_1 gpc652 (
      {stage0_4[239]},
      {stage1_4[132]}
   );
   gpc1_1 gpc653 (
      {stage0_4[240]},
      {stage1_4[133]}
   );
   gpc1_1 gpc654 (
      {stage0_4[241]},
      {stage1_4[134]}
   );
   gpc1_1 gpc655 (
      {stage0_4[242]},
      {stage1_4[135]}
   );
   gpc1_1 gpc656 (
      {stage0_4[243]},
      {stage1_4[136]}
   );
   gpc1_1 gpc657 (
      {stage0_4[244]},
      {stage1_4[137]}
   );
   gpc1_1 gpc658 (
      {stage0_4[245]},
      {stage1_4[138]}
   );
   gpc1_1 gpc659 (
      {stage0_4[246]},
      {stage1_4[139]}
   );
   gpc1_1 gpc660 (
      {stage0_4[247]},
      {stage1_4[140]}
   );
   gpc1_1 gpc661 (
      {stage0_4[248]},
      {stage1_4[141]}
   );
   gpc1_1 gpc662 (
      {stage0_4[249]},
      {stage1_4[142]}
   );
   gpc1_1 gpc663 (
      {stage0_4[250]},
      {stage1_4[143]}
   );
   gpc1_1 gpc664 (
      {stage0_4[251]},
      {stage1_4[144]}
   );
   gpc1_1 gpc665 (
      {stage0_4[252]},
      {stage1_4[145]}
   );
   gpc1_1 gpc666 (
      {stage0_4[253]},
      {stage1_4[146]}
   );
   gpc1_1 gpc667 (
      {stage0_4[254]},
      {stage1_4[147]}
   );
   gpc1_1 gpc668 (
      {stage0_4[255]},
      {stage1_4[148]}
   );
   gpc1_1 gpc669 (
      {stage0_5[240]},
      {stage1_5[110]}
   );
   gpc1_1 gpc670 (
      {stage0_5[241]},
      {stage1_5[111]}
   );
   gpc1_1 gpc671 (
      {stage0_5[242]},
      {stage1_5[112]}
   );
   gpc1_1 gpc672 (
      {stage0_5[243]},
      {stage1_5[113]}
   );
   gpc1_1 gpc673 (
      {stage0_5[244]},
      {stage1_5[114]}
   );
   gpc1_1 gpc674 (
      {stage0_5[245]},
      {stage1_5[115]}
   );
   gpc1_1 gpc675 (
      {stage0_5[246]},
      {stage1_5[116]}
   );
   gpc1_1 gpc676 (
      {stage0_5[247]},
      {stage1_5[117]}
   );
   gpc1_1 gpc677 (
      {stage0_5[248]},
      {stage1_5[118]}
   );
   gpc1_1 gpc678 (
      {stage0_5[249]},
      {stage1_5[119]}
   );
   gpc1_1 gpc679 (
      {stage0_5[250]},
      {stage1_5[120]}
   );
   gpc1_1 gpc680 (
      {stage0_5[251]},
      {stage1_5[121]}
   );
   gpc1_1 gpc681 (
      {stage0_5[252]},
      {stage1_5[122]}
   );
   gpc1_1 gpc682 (
      {stage0_5[253]},
      {stage1_5[123]}
   );
   gpc1_1 gpc683 (
      {stage0_5[254]},
      {stage1_5[124]}
   );
   gpc1_1 gpc684 (
      {stage0_5[255]},
      {stage1_5[125]}
   );
   gpc1_1 gpc685 (
      {stage0_6[243]},
      {stage1_6[83]}
   );
   gpc1_1 gpc686 (
      {stage0_6[244]},
      {stage1_6[84]}
   );
   gpc1_1 gpc687 (
      {stage0_6[245]},
      {stage1_6[85]}
   );
   gpc1_1 gpc688 (
      {stage0_6[246]},
      {stage1_6[86]}
   );
   gpc1_1 gpc689 (
      {stage0_6[247]},
      {stage1_6[87]}
   );
   gpc1_1 gpc690 (
      {stage0_6[248]},
      {stage1_6[88]}
   );
   gpc1_1 gpc691 (
      {stage0_6[249]},
      {stage1_6[89]}
   );
   gpc1_1 gpc692 (
      {stage0_6[250]},
      {stage1_6[90]}
   );
   gpc1_1 gpc693 (
      {stage0_6[251]},
      {stage1_6[91]}
   );
   gpc1_1 gpc694 (
      {stage0_6[252]},
      {stage1_6[92]}
   );
   gpc1_1 gpc695 (
      {stage0_6[253]},
      {stage1_6[93]}
   );
   gpc1_1 gpc696 (
      {stage0_6[254]},
      {stage1_6[94]}
   );
   gpc1_1 gpc697 (
      {stage0_6[255]},
      {stage1_6[95]}
   );
   gpc1_1 gpc698 (
      {stage0_7[251]},
      {stage1_7[96]}
   );
   gpc1_1 gpc699 (
      {stage0_7[252]},
      {stage1_7[97]}
   );
   gpc1_1 gpc700 (
      {stage0_7[253]},
      {stage1_7[98]}
   );
   gpc1_1 gpc701 (
      {stage0_7[254]},
      {stage1_7[99]}
   );
   gpc1_1 gpc702 (
      {stage0_7[255]},
      {stage1_7[100]}
   );
   gpc1_1 gpc703 (
      {stage0_9[230]},
      {stage1_9[106]}
   );
   gpc1_1 gpc704 (
      {stage0_9[231]},
      {stage1_9[107]}
   );
   gpc1_1 gpc705 (
      {stage0_9[232]},
      {stage1_9[108]}
   );
   gpc1_1 gpc706 (
      {stage0_9[233]},
      {stage1_9[109]}
   );
   gpc1_1 gpc707 (
      {stage0_9[234]},
      {stage1_9[110]}
   );
   gpc1_1 gpc708 (
      {stage0_9[235]},
      {stage1_9[111]}
   );
   gpc1_1 gpc709 (
      {stage0_9[236]},
      {stage1_9[112]}
   );
   gpc1_1 gpc710 (
      {stage0_9[237]},
      {stage1_9[113]}
   );
   gpc1_1 gpc711 (
      {stage0_9[238]},
      {stage1_9[114]}
   );
   gpc1_1 gpc712 (
      {stage0_9[239]},
      {stage1_9[115]}
   );
   gpc1_1 gpc713 (
      {stage0_9[240]},
      {stage1_9[116]}
   );
   gpc1_1 gpc714 (
      {stage0_9[241]},
      {stage1_9[117]}
   );
   gpc1_1 gpc715 (
      {stage0_9[242]},
      {stage1_9[118]}
   );
   gpc1_1 gpc716 (
      {stage0_9[243]},
      {stage1_9[119]}
   );
   gpc1_1 gpc717 (
      {stage0_9[244]},
      {stage1_9[120]}
   );
   gpc1_1 gpc718 (
      {stage0_9[245]},
      {stage1_9[121]}
   );
   gpc1_1 gpc719 (
      {stage0_9[246]},
      {stage1_9[122]}
   );
   gpc1_1 gpc720 (
      {stage0_9[247]},
      {stage1_9[123]}
   );
   gpc1_1 gpc721 (
      {stage0_9[248]},
      {stage1_9[124]}
   );
   gpc1_1 gpc722 (
      {stage0_9[249]},
      {stage1_9[125]}
   );
   gpc1_1 gpc723 (
      {stage0_9[250]},
      {stage1_9[126]}
   );
   gpc1_1 gpc724 (
      {stage0_9[251]},
      {stage1_9[127]}
   );
   gpc1_1 gpc725 (
      {stage0_9[252]},
      {stage1_9[128]}
   );
   gpc1_1 gpc726 (
      {stage0_9[253]},
      {stage1_9[129]}
   );
   gpc1_1 gpc727 (
      {stage0_9[254]},
      {stage1_9[130]}
   );
   gpc1_1 gpc728 (
      {stage0_9[255]},
      {stage1_9[131]}
   );
   gpc1_1 gpc729 (
      {stage0_10[250]},
      {stage1_10[91]}
   );
   gpc1_1 gpc730 (
      {stage0_10[251]},
      {stage1_10[92]}
   );
   gpc1_1 gpc731 (
      {stage0_10[252]},
      {stage1_10[93]}
   );
   gpc1_1 gpc732 (
      {stage0_10[253]},
      {stage1_10[94]}
   );
   gpc1_1 gpc733 (
      {stage0_10[254]},
      {stage1_10[95]}
   );
   gpc1_1 gpc734 (
      {stage0_10[255]},
      {stage1_10[96]}
   );
   gpc1_1 gpc735 (
      {stage0_11[210]},
      {stage1_11[94]}
   );
   gpc1_1 gpc736 (
      {stage0_11[211]},
      {stage1_11[95]}
   );
   gpc1_1 gpc737 (
      {stage0_11[212]},
      {stage1_11[96]}
   );
   gpc1_1 gpc738 (
      {stage0_11[213]},
      {stage1_11[97]}
   );
   gpc1_1 gpc739 (
      {stage0_11[214]},
      {stage1_11[98]}
   );
   gpc1_1 gpc740 (
      {stage0_11[215]},
      {stage1_11[99]}
   );
   gpc1_1 gpc741 (
      {stage0_11[216]},
      {stage1_11[100]}
   );
   gpc1_1 gpc742 (
      {stage0_11[217]},
      {stage1_11[101]}
   );
   gpc1_1 gpc743 (
      {stage0_11[218]},
      {stage1_11[102]}
   );
   gpc1_1 gpc744 (
      {stage0_11[219]},
      {stage1_11[103]}
   );
   gpc1_1 gpc745 (
      {stage0_11[220]},
      {stage1_11[104]}
   );
   gpc1_1 gpc746 (
      {stage0_11[221]},
      {stage1_11[105]}
   );
   gpc1_1 gpc747 (
      {stage0_11[222]},
      {stage1_11[106]}
   );
   gpc1_1 gpc748 (
      {stage0_11[223]},
      {stage1_11[107]}
   );
   gpc1_1 gpc749 (
      {stage0_11[224]},
      {stage1_11[108]}
   );
   gpc1_1 gpc750 (
      {stage0_11[225]},
      {stage1_11[109]}
   );
   gpc1_1 gpc751 (
      {stage0_11[226]},
      {stage1_11[110]}
   );
   gpc1_1 gpc752 (
      {stage0_11[227]},
      {stage1_11[111]}
   );
   gpc1_1 gpc753 (
      {stage0_11[228]},
      {stage1_11[112]}
   );
   gpc1_1 gpc754 (
      {stage0_11[229]},
      {stage1_11[113]}
   );
   gpc1_1 gpc755 (
      {stage0_11[230]},
      {stage1_11[114]}
   );
   gpc1_1 gpc756 (
      {stage0_11[231]},
      {stage1_11[115]}
   );
   gpc1_1 gpc757 (
      {stage0_11[232]},
      {stage1_11[116]}
   );
   gpc1_1 gpc758 (
      {stage0_11[233]},
      {stage1_11[117]}
   );
   gpc1_1 gpc759 (
      {stage0_11[234]},
      {stage1_11[118]}
   );
   gpc1_1 gpc760 (
      {stage0_11[235]},
      {stage1_11[119]}
   );
   gpc1_1 gpc761 (
      {stage0_11[236]},
      {stage1_11[120]}
   );
   gpc1_1 gpc762 (
      {stage0_11[237]},
      {stage1_11[121]}
   );
   gpc1_1 gpc763 (
      {stage0_11[238]},
      {stage1_11[122]}
   );
   gpc1_1 gpc764 (
      {stage0_11[239]},
      {stage1_11[123]}
   );
   gpc1_1 gpc765 (
      {stage0_11[240]},
      {stage1_11[124]}
   );
   gpc1_1 gpc766 (
      {stage0_11[241]},
      {stage1_11[125]}
   );
   gpc1_1 gpc767 (
      {stage0_11[242]},
      {stage1_11[126]}
   );
   gpc1_1 gpc768 (
      {stage0_11[243]},
      {stage1_11[127]}
   );
   gpc1_1 gpc769 (
      {stage0_11[244]},
      {stage1_11[128]}
   );
   gpc1_1 gpc770 (
      {stage0_11[245]},
      {stage1_11[129]}
   );
   gpc1_1 gpc771 (
      {stage0_11[246]},
      {stage1_11[130]}
   );
   gpc1_1 gpc772 (
      {stage0_11[247]},
      {stage1_11[131]}
   );
   gpc1_1 gpc773 (
      {stage0_11[248]},
      {stage1_11[132]}
   );
   gpc1_1 gpc774 (
      {stage0_11[249]},
      {stage1_11[133]}
   );
   gpc1_1 gpc775 (
      {stage0_11[250]},
      {stage1_11[134]}
   );
   gpc1_1 gpc776 (
      {stage0_11[251]},
      {stage1_11[135]}
   );
   gpc1_1 gpc777 (
      {stage0_11[252]},
      {stage1_11[136]}
   );
   gpc1_1 gpc778 (
      {stage0_11[253]},
      {stage1_11[137]}
   );
   gpc1_1 gpc779 (
      {stage0_11[254]},
      {stage1_11[138]}
   );
   gpc1_1 gpc780 (
      {stage0_11[255]},
      {stage1_11[139]}
   );
   gpc1_1 gpc781 (
      {stage0_12[148]},
      {stage1_12[90]}
   );
   gpc1_1 gpc782 (
      {stage0_12[149]},
      {stage1_12[91]}
   );
   gpc1_1 gpc783 (
      {stage0_12[150]},
      {stage1_12[92]}
   );
   gpc1_1 gpc784 (
      {stage0_12[151]},
      {stage1_12[93]}
   );
   gpc1_1 gpc785 (
      {stage0_12[152]},
      {stage1_12[94]}
   );
   gpc1_1 gpc786 (
      {stage0_12[153]},
      {stage1_12[95]}
   );
   gpc1_1 gpc787 (
      {stage0_12[154]},
      {stage1_12[96]}
   );
   gpc1_1 gpc788 (
      {stage0_12[155]},
      {stage1_12[97]}
   );
   gpc1_1 gpc789 (
      {stage0_12[156]},
      {stage1_12[98]}
   );
   gpc1_1 gpc790 (
      {stage0_12[157]},
      {stage1_12[99]}
   );
   gpc1_1 gpc791 (
      {stage0_12[158]},
      {stage1_12[100]}
   );
   gpc1_1 gpc792 (
      {stage0_12[159]},
      {stage1_12[101]}
   );
   gpc1_1 gpc793 (
      {stage0_12[160]},
      {stage1_12[102]}
   );
   gpc1_1 gpc794 (
      {stage0_12[161]},
      {stage1_12[103]}
   );
   gpc1_1 gpc795 (
      {stage0_12[162]},
      {stage1_12[104]}
   );
   gpc1_1 gpc796 (
      {stage0_12[163]},
      {stage1_12[105]}
   );
   gpc1_1 gpc797 (
      {stage0_12[164]},
      {stage1_12[106]}
   );
   gpc1_1 gpc798 (
      {stage0_12[165]},
      {stage1_12[107]}
   );
   gpc1_1 gpc799 (
      {stage0_12[166]},
      {stage1_12[108]}
   );
   gpc1_1 gpc800 (
      {stage0_12[167]},
      {stage1_12[109]}
   );
   gpc1_1 gpc801 (
      {stage0_12[168]},
      {stage1_12[110]}
   );
   gpc1_1 gpc802 (
      {stage0_12[169]},
      {stage1_12[111]}
   );
   gpc1_1 gpc803 (
      {stage0_12[170]},
      {stage1_12[112]}
   );
   gpc1_1 gpc804 (
      {stage0_12[171]},
      {stage1_12[113]}
   );
   gpc1_1 gpc805 (
      {stage0_12[172]},
      {stage1_12[114]}
   );
   gpc1_1 gpc806 (
      {stage0_12[173]},
      {stage1_12[115]}
   );
   gpc1_1 gpc807 (
      {stage0_12[174]},
      {stage1_12[116]}
   );
   gpc1_1 gpc808 (
      {stage0_12[175]},
      {stage1_12[117]}
   );
   gpc1_1 gpc809 (
      {stage0_12[176]},
      {stage1_12[118]}
   );
   gpc1_1 gpc810 (
      {stage0_12[177]},
      {stage1_12[119]}
   );
   gpc1_1 gpc811 (
      {stage0_12[178]},
      {stage1_12[120]}
   );
   gpc1_1 gpc812 (
      {stage0_12[179]},
      {stage1_12[121]}
   );
   gpc1_1 gpc813 (
      {stage0_12[180]},
      {stage1_12[122]}
   );
   gpc1_1 gpc814 (
      {stage0_12[181]},
      {stage1_12[123]}
   );
   gpc1_1 gpc815 (
      {stage0_12[182]},
      {stage1_12[124]}
   );
   gpc1_1 gpc816 (
      {stage0_12[183]},
      {stage1_12[125]}
   );
   gpc1_1 gpc817 (
      {stage0_12[184]},
      {stage1_12[126]}
   );
   gpc1_1 gpc818 (
      {stage0_12[185]},
      {stage1_12[127]}
   );
   gpc1_1 gpc819 (
      {stage0_12[186]},
      {stage1_12[128]}
   );
   gpc1_1 gpc820 (
      {stage0_12[187]},
      {stage1_12[129]}
   );
   gpc1_1 gpc821 (
      {stage0_12[188]},
      {stage1_12[130]}
   );
   gpc1_1 gpc822 (
      {stage0_12[189]},
      {stage1_12[131]}
   );
   gpc1_1 gpc823 (
      {stage0_12[190]},
      {stage1_12[132]}
   );
   gpc1_1 gpc824 (
      {stage0_12[191]},
      {stage1_12[133]}
   );
   gpc1_1 gpc825 (
      {stage0_12[192]},
      {stage1_12[134]}
   );
   gpc1_1 gpc826 (
      {stage0_12[193]},
      {stage1_12[135]}
   );
   gpc1_1 gpc827 (
      {stage0_12[194]},
      {stage1_12[136]}
   );
   gpc1_1 gpc828 (
      {stage0_12[195]},
      {stage1_12[137]}
   );
   gpc1_1 gpc829 (
      {stage0_12[196]},
      {stage1_12[138]}
   );
   gpc1_1 gpc830 (
      {stage0_12[197]},
      {stage1_12[139]}
   );
   gpc1_1 gpc831 (
      {stage0_12[198]},
      {stage1_12[140]}
   );
   gpc1_1 gpc832 (
      {stage0_12[199]},
      {stage1_12[141]}
   );
   gpc1_1 gpc833 (
      {stage0_12[200]},
      {stage1_12[142]}
   );
   gpc1_1 gpc834 (
      {stage0_12[201]},
      {stage1_12[143]}
   );
   gpc1_1 gpc835 (
      {stage0_12[202]},
      {stage1_12[144]}
   );
   gpc1_1 gpc836 (
      {stage0_12[203]},
      {stage1_12[145]}
   );
   gpc1_1 gpc837 (
      {stage0_12[204]},
      {stage1_12[146]}
   );
   gpc1_1 gpc838 (
      {stage0_12[205]},
      {stage1_12[147]}
   );
   gpc1_1 gpc839 (
      {stage0_12[206]},
      {stage1_12[148]}
   );
   gpc1_1 gpc840 (
      {stage0_12[207]},
      {stage1_12[149]}
   );
   gpc1_1 gpc841 (
      {stage0_12[208]},
      {stage1_12[150]}
   );
   gpc1_1 gpc842 (
      {stage0_12[209]},
      {stage1_12[151]}
   );
   gpc1_1 gpc843 (
      {stage0_12[210]},
      {stage1_12[152]}
   );
   gpc1_1 gpc844 (
      {stage0_12[211]},
      {stage1_12[153]}
   );
   gpc1_1 gpc845 (
      {stage0_12[212]},
      {stage1_12[154]}
   );
   gpc1_1 gpc846 (
      {stage0_12[213]},
      {stage1_12[155]}
   );
   gpc1_1 gpc847 (
      {stage0_12[214]},
      {stage1_12[156]}
   );
   gpc1_1 gpc848 (
      {stage0_12[215]},
      {stage1_12[157]}
   );
   gpc1_1 gpc849 (
      {stage0_12[216]},
      {stage1_12[158]}
   );
   gpc1_1 gpc850 (
      {stage0_12[217]},
      {stage1_12[159]}
   );
   gpc1_1 gpc851 (
      {stage0_12[218]},
      {stage1_12[160]}
   );
   gpc1_1 gpc852 (
      {stage0_12[219]},
      {stage1_12[161]}
   );
   gpc1_1 gpc853 (
      {stage0_12[220]},
      {stage1_12[162]}
   );
   gpc1_1 gpc854 (
      {stage0_12[221]},
      {stage1_12[163]}
   );
   gpc1_1 gpc855 (
      {stage0_12[222]},
      {stage1_12[164]}
   );
   gpc1_1 gpc856 (
      {stage0_12[223]},
      {stage1_12[165]}
   );
   gpc1_1 gpc857 (
      {stage0_12[224]},
      {stage1_12[166]}
   );
   gpc1_1 gpc858 (
      {stage0_12[225]},
      {stage1_12[167]}
   );
   gpc1_1 gpc859 (
      {stage0_12[226]},
      {stage1_12[168]}
   );
   gpc1_1 gpc860 (
      {stage0_12[227]},
      {stage1_12[169]}
   );
   gpc1_1 gpc861 (
      {stage0_12[228]},
      {stage1_12[170]}
   );
   gpc1_1 gpc862 (
      {stage0_12[229]},
      {stage1_12[171]}
   );
   gpc1_1 gpc863 (
      {stage0_12[230]},
      {stage1_12[172]}
   );
   gpc1_1 gpc864 (
      {stage0_12[231]},
      {stage1_12[173]}
   );
   gpc1_1 gpc865 (
      {stage0_12[232]},
      {stage1_12[174]}
   );
   gpc1_1 gpc866 (
      {stage0_12[233]},
      {stage1_12[175]}
   );
   gpc1_1 gpc867 (
      {stage0_12[234]},
      {stage1_12[176]}
   );
   gpc1_1 gpc868 (
      {stage0_12[235]},
      {stage1_12[177]}
   );
   gpc1_1 gpc869 (
      {stage0_12[236]},
      {stage1_12[178]}
   );
   gpc1_1 gpc870 (
      {stage0_12[237]},
      {stage1_12[179]}
   );
   gpc1_1 gpc871 (
      {stage0_12[238]},
      {stage1_12[180]}
   );
   gpc1_1 gpc872 (
      {stage0_12[239]},
      {stage1_12[181]}
   );
   gpc1_1 gpc873 (
      {stage0_12[240]},
      {stage1_12[182]}
   );
   gpc1_1 gpc874 (
      {stage0_12[241]},
      {stage1_12[183]}
   );
   gpc1_1 gpc875 (
      {stage0_12[242]},
      {stage1_12[184]}
   );
   gpc1_1 gpc876 (
      {stage0_12[243]},
      {stage1_12[185]}
   );
   gpc1_1 gpc877 (
      {stage0_12[244]},
      {stage1_12[186]}
   );
   gpc1_1 gpc878 (
      {stage0_12[245]},
      {stage1_12[187]}
   );
   gpc1_1 gpc879 (
      {stage0_12[246]},
      {stage1_12[188]}
   );
   gpc1_1 gpc880 (
      {stage0_12[247]},
      {stage1_12[189]}
   );
   gpc1_1 gpc881 (
      {stage0_12[248]},
      {stage1_12[190]}
   );
   gpc1_1 gpc882 (
      {stage0_12[249]},
      {stage1_12[191]}
   );
   gpc1_1 gpc883 (
      {stage0_12[250]},
      {stage1_12[192]}
   );
   gpc1_1 gpc884 (
      {stage0_12[251]},
      {stage1_12[193]}
   );
   gpc1_1 gpc885 (
      {stage0_12[252]},
      {stage1_12[194]}
   );
   gpc1_1 gpc886 (
      {stage0_12[253]},
      {stage1_12[195]}
   );
   gpc1_1 gpc887 (
      {stage0_12[254]},
      {stage1_12[196]}
   );
   gpc1_1 gpc888 (
      {stage0_12[255]},
      {stage1_12[197]}
   );
   gpc1_1 gpc889 (
      {stage0_14[235]},
      {stage1_14[93]}
   );
   gpc1_1 gpc890 (
      {stage0_14[236]},
      {stage1_14[94]}
   );
   gpc1_1 gpc891 (
      {stage0_14[237]},
      {stage1_14[95]}
   );
   gpc1_1 gpc892 (
      {stage0_14[238]},
      {stage1_14[96]}
   );
   gpc1_1 gpc893 (
      {stage0_14[239]},
      {stage1_14[97]}
   );
   gpc1_1 gpc894 (
      {stage0_14[240]},
      {stage1_14[98]}
   );
   gpc1_1 gpc895 (
      {stage0_14[241]},
      {stage1_14[99]}
   );
   gpc1_1 gpc896 (
      {stage0_14[242]},
      {stage1_14[100]}
   );
   gpc1_1 gpc897 (
      {stage0_14[243]},
      {stage1_14[101]}
   );
   gpc1_1 gpc898 (
      {stage0_14[244]},
      {stage1_14[102]}
   );
   gpc1_1 gpc899 (
      {stage0_14[245]},
      {stage1_14[103]}
   );
   gpc1_1 gpc900 (
      {stage0_14[246]},
      {stage1_14[104]}
   );
   gpc1_1 gpc901 (
      {stage0_14[247]},
      {stage1_14[105]}
   );
   gpc1_1 gpc902 (
      {stage0_14[248]},
      {stage1_14[106]}
   );
   gpc1_1 gpc903 (
      {stage0_14[249]},
      {stage1_14[107]}
   );
   gpc1_1 gpc904 (
      {stage0_14[250]},
      {stage1_14[108]}
   );
   gpc1_1 gpc905 (
      {stage0_14[251]},
      {stage1_14[109]}
   );
   gpc1_1 gpc906 (
      {stage0_14[252]},
      {stage1_14[110]}
   );
   gpc1_1 gpc907 (
      {stage0_14[253]},
      {stage1_14[111]}
   );
   gpc1_1 gpc908 (
      {stage0_14[254]},
      {stage1_14[112]}
   );
   gpc1_1 gpc909 (
      {stage0_14[255]},
      {stage1_14[113]}
   );
   gpc1_1 gpc910 (
      {stage0_15[254]},
      {stage1_15[91]}
   );
   gpc1_1 gpc911 (
      {stage0_15[255]},
      {stage1_15[92]}
   );
   gpc1_1 gpc912 (
      {stage0_17[252]},
      {stage1_17[123]}
   );
   gpc1_1 gpc913 (
      {stage0_17[253]},
      {stage1_17[124]}
   );
   gpc1_1 gpc914 (
      {stage0_17[254]},
      {stage1_17[125]}
   );
   gpc1_1 gpc915 (
      {stage0_17[255]},
      {stage1_17[126]}
   );
   gpc1_1 gpc916 (
      {stage0_18[204]},
      {stage1_18[99]}
   );
   gpc1_1 gpc917 (
      {stage0_18[205]},
      {stage1_18[100]}
   );
   gpc1_1 gpc918 (
      {stage0_18[206]},
      {stage1_18[101]}
   );
   gpc1_1 gpc919 (
      {stage0_18[207]},
      {stage1_18[102]}
   );
   gpc1_1 gpc920 (
      {stage0_18[208]},
      {stage1_18[103]}
   );
   gpc1_1 gpc921 (
      {stage0_18[209]},
      {stage1_18[104]}
   );
   gpc1_1 gpc922 (
      {stage0_18[210]},
      {stage1_18[105]}
   );
   gpc1_1 gpc923 (
      {stage0_18[211]},
      {stage1_18[106]}
   );
   gpc1_1 gpc924 (
      {stage0_18[212]},
      {stage1_18[107]}
   );
   gpc1_1 gpc925 (
      {stage0_18[213]},
      {stage1_18[108]}
   );
   gpc1_1 gpc926 (
      {stage0_18[214]},
      {stage1_18[109]}
   );
   gpc1_1 gpc927 (
      {stage0_18[215]},
      {stage1_18[110]}
   );
   gpc1_1 gpc928 (
      {stage0_18[216]},
      {stage1_18[111]}
   );
   gpc1_1 gpc929 (
      {stage0_18[217]},
      {stage1_18[112]}
   );
   gpc1_1 gpc930 (
      {stage0_18[218]},
      {stage1_18[113]}
   );
   gpc1_1 gpc931 (
      {stage0_18[219]},
      {stage1_18[114]}
   );
   gpc1_1 gpc932 (
      {stage0_18[220]},
      {stage1_18[115]}
   );
   gpc1_1 gpc933 (
      {stage0_18[221]},
      {stage1_18[116]}
   );
   gpc1_1 gpc934 (
      {stage0_18[222]},
      {stage1_18[117]}
   );
   gpc1_1 gpc935 (
      {stage0_18[223]},
      {stage1_18[118]}
   );
   gpc1_1 gpc936 (
      {stage0_18[224]},
      {stage1_18[119]}
   );
   gpc1_1 gpc937 (
      {stage0_18[225]},
      {stage1_18[120]}
   );
   gpc1_1 gpc938 (
      {stage0_18[226]},
      {stage1_18[121]}
   );
   gpc1_1 gpc939 (
      {stage0_18[227]},
      {stage1_18[122]}
   );
   gpc1_1 gpc940 (
      {stage0_18[228]},
      {stage1_18[123]}
   );
   gpc1_1 gpc941 (
      {stage0_18[229]},
      {stage1_18[124]}
   );
   gpc1_1 gpc942 (
      {stage0_18[230]},
      {stage1_18[125]}
   );
   gpc1_1 gpc943 (
      {stage0_18[231]},
      {stage1_18[126]}
   );
   gpc1_1 gpc944 (
      {stage0_18[232]},
      {stage1_18[127]}
   );
   gpc1_1 gpc945 (
      {stage0_18[233]},
      {stage1_18[128]}
   );
   gpc1_1 gpc946 (
      {stage0_18[234]},
      {stage1_18[129]}
   );
   gpc1_1 gpc947 (
      {stage0_18[235]},
      {stage1_18[130]}
   );
   gpc1_1 gpc948 (
      {stage0_18[236]},
      {stage1_18[131]}
   );
   gpc1_1 gpc949 (
      {stage0_18[237]},
      {stage1_18[132]}
   );
   gpc1_1 gpc950 (
      {stage0_18[238]},
      {stage1_18[133]}
   );
   gpc1_1 gpc951 (
      {stage0_18[239]},
      {stage1_18[134]}
   );
   gpc1_1 gpc952 (
      {stage0_18[240]},
      {stage1_18[135]}
   );
   gpc1_1 gpc953 (
      {stage0_18[241]},
      {stage1_18[136]}
   );
   gpc1_1 gpc954 (
      {stage0_18[242]},
      {stage1_18[137]}
   );
   gpc1_1 gpc955 (
      {stage0_18[243]},
      {stage1_18[138]}
   );
   gpc1_1 gpc956 (
      {stage0_18[244]},
      {stage1_18[139]}
   );
   gpc1_1 gpc957 (
      {stage0_18[245]},
      {stage1_18[140]}
   );
   gpc1_1 gpc958 (
      {stage0_18[246]},
      {stage1_18[141]}
   );
   gpc1_1 gpc959 (
      {stage0_18[247]},
      {stage1_18[142]}
   );
   gpc1_1 gpc960 (
      {stage0_18[248]},
      {stage1_18[143]}
   );
   gpc1_1 gpc961 (
      {stage0_18[249]},
      {stage1_18[144]}
   );
   gpc1_1 gpc962 (
      {stage0_18[250]},
      {stage1_18[145]}
   );
   gpc1_1 gpc963 (
      {stage0_18[251]},
      {stage1_18[146]}
   );
   gpc1_1 gpc964 (
      {stage0_18[252]},
      {stage1_18[147]}
   );
   gpc1_1 gpc965 (
      {stage0_18[253]},
      {stage1_18[148]}
   );
   gpc1_1 gpc966 (
      {stage0_18[254]},
      {stage1_18[149]}
   );
   gpc1_1 gpc967 (
      {stage0_18[255]},
      {stage1_18[150]}
   );
   gpc1_1 gpc968 (
      {stage0_19[240]},
      {stage1_19[78]}
   );
   gpc1_1 gpc969 (
      {stage0_19[241]},
      {stage1_19[79]}
   );
   gpc1_1 gpc970 (
      {stage0_19[242]},
      {stage1_19[80]}
   );
   gpc1_1 gpc971 (
      {stage0_19[243]},
      {stage1_19[81]}
   );
   gpc1_1 gpc972 (
      {stage0_19[244]},
      {stage1_19[82]}
   );
   gpc1_1 gpc973 (
      {stage0_19[245]},
      {stage1_19[83]}
   );
   gpc1_1 gpc974 (
      {stage0_19[246]},
      {stage1_19[84]}
   );
   gpc1_1 gpc975 (
      {stage0_19[247]},
      {stage1_19[85]}
   );
   gpc1_1 gpc976 (
      {stage0_19[248]},
      {stage1_19[86]}
   );
   gpc1_1 gpc977 (
      {stage0_19[249]},
      {stage1_19[87]}
   );
   gpc1_1 gpc978 (
      {stage0_19[250]},
      {stage1_19[88]}
   );
   gpc1_1 gpc979 (
      {stage0_19[251]},
      {stage1_19[89]}
   );
   gpc1_1 gpc980 (
      {stage0_19[252]},
      {stage1_19[90]}
   );
   gpc1_1 gpc981 (
      {stage0_19[253]},
      {stage1_19[91]}
   );
   gpc1_1 gpc982 (
      {stage0_19[254]},
      {stage1_19[92]}
   );
   gpc1_1 gpc983 (
      {stage0_19[255]},
      {stage1_19[93]}
   );
   gpc1_1 gpc984 (
      {stage0_20[245]},
      {stage1_20[105]}
   );
   gpc1_1 gpc985 (
      {stage0_20[246]},
      {stage1_20[106]}
   );
   gpc1_1 gpc986 (
      {stage0_20[247]},
      {stage1_20[107]}
   );
   gpc1_1 gpc987 (
      {stage0_20[248]},
      {stage1_20[108]}
   );
   gpc1_1 gpc988 (
      {stage0_20[249]},
      {stage1_20[109]}
   );
   gpc1_1 gpc989 (
      {stage0_20[250]},
      {stage1_20[110]}
   );
   gpc1_1 gpc990 (
      {stage0_20[251]},
      {stage1_20[111]}
   );
   gpc1_1 gpc991 (
      {stage0_20[252]},
      {stage1_20[112]}
   );
   gpc1_1 gpc992 (
      {stage0_20[253]},
      {stage1_20[113]}
   );
   gpc1_1 gpc993 (
      {stage0_20[254]},
      {stage1_20[114]}
   );
   gpc1_1 gpc994 (
      {stage0_20[255]},
      {stage1_20[115]}
   );
   gpc1_1 gpc995 (
      {stage0_21[235]},
      {stage1_21[118]}
   );
   gpc1_1 gpc996 (
      {stage0_21[236]},
      {stage1_21[119]}
   );
   gpc1_1 gpc997 (
      {stage0_21[237]},
      {stage1_21[120]}
   );
   gpc1_1 gpc998 (
      {stage0_21[238]},
      {stage1_21[121]}
   );
   gpc1_1 gpc999 (
      {stage0_21[239]},
      {stage1_21[122]}
   );
   gpc1_1 gpc1000 (
      {stage0_21[240]},
      {stage1_21[123]}
   );
   gpc1_1 gpc1001 (
      {stage0_21[241]},
      {stage1_21[124]}
   );
   gpc1_1 gpc1002 (
      {stage0_21[242]},
      {stage1_21[125]}
   );
   gpc1_1 gpc1003 (
      {stage0_21[243]},
      {stage1_21[126]}
   );
   gpc1_1 gpc1004 (
      {stage0_21[244]},
      {stage1_21[127]}
   );
   gpc1_1 gpc1005 (
      {stage0_21[245]},
      {stage1_21[128]}
   );
   gpc1_1 gpc1006 (
      {stage0_21[246]},
      {stage1_21[129]}
   );
   gpc1_1 gpc1007 (
      {stage0_21[247]},
      {stage1_21[130]}
   );
   gpc1_1 gpc1008 (
      {stage0_21[248]},
      {stage1_21[131]}
   );
   gpc1_1 gpc1009 (
      {stage0_21[249]},
      {stage1_21[132]}
   );
   gpc1_1 gpc1010 (
      {stage0_21[250]},
      {stage1_21[133]}
   );
   gpc1_1 gpc1011 (
      {stage0_21[251]},
      {stage1_21[134]}
   );
   gpc1_1 gpc1012 (
      {stage0_21[252]},
      {stage1_21[135]}
   );
   gpc1_1 gpc1013 (
      {stage0_21[253]},
      {stage1_21[136]}
   );
   gpc1_1 gpc1014 (
      {stage0_21[254]},
      {stage1_21[137]}
   );
   gpc1_1 gpc1015 (
      {stage0_21[255]},
      {stage1_21[138]}
   );
   gpc1_1 gpc1016 (
      {stage0_22[246]},
      {stage1_22[84]}
   );
   gpc1_1 gpc1017 (
      {stage0_22[247]},
      {stage1_22[85]}
   );
   gpc1_1 gpc1018 (
      {stage0_22[248]},
      {stage1_22[86]}
   );
   gpc1_1 gpc1019 (
      {stage0_22[249]},
      {stage1_22[87]}
   );
   gpc1_1 gpc1020 (
      {stage0_22[250]},
      {stage1_22[88]}
   );
   gpc1_1 gpc1021 (
      {stage0_22[251]},
      {stage1_22[89]}
   );
   gpc1_1 gpc1022 (
      {stage0_22[252]},
      {stage1_22[90]}
   );
   gpc1_1 gpc1023 (
      {stage0_22[253]},
      {stage1_22[91]}
   );
   gpc1_1 gpc1024 (
      {stage0_22[254]},
      {stage1_22[92]}
   );
   gpc1_1 gpc1025 (
      {stage0_22[255]},
      {stage1_22[93]}
   );
   gpc1_1 gpc1026 (
      {stage0_23[246]},
      {stage1_23[84]}
   );
   gpc1_1 gpc1027 (
      {stage0_23[247]},
      {stage1_23[85]}
   );
   gpc1_1 gpc1028 (
      {stage0_23[248]},
      {stage1_23[86]}
   );
   gpc1_1 gpc1029 (
      {stage0_23[249]},
      {stage1_23[87]}
   );
   gpc1_1 gpc1030 (
      {stage0_23[250]},
      {stage1_23[88]}
   );
   gpc1_1 gpc1031 (
      {stage0_23[251]},
      {stage1_23[89]}
   );
   gpc1_1 gpc1032 (
      {stage0_23[252]},
      {stage1_23[90]}
   );
   gpc1_1 gpc1033 (
      {stage0_23[253]},
      {stage1_23[91]}
   );
   gpc1_1 gpc1034 (
      {stage0_23[254]},
      {stage1_23[92]}
   );
   gpc1_1 gpc1035 (
      {stage0_23[255]},
      {stage1_23[93]}
   );
   gpc1_1 gpc1036 (
      {stage0_24[96]},
      {stage1_24[94]}
   );
   gpc1_1 gpc1037 (
      {stage0_24[97]},
      {stage1_24[95]}
   );
   gpc1_1 gpc1038 (
      {stage0_24[98]},
      {stage1_24[96]}
   );
   gpc1_1 gpc1039 (
      {stage0_24[99]},
      {stage1_24[97]}
   );
   gpc1_1 gpc1040 (
      {stage0_24[100]},
      {stage1_24[98]}
   );
   gpc1_1 gpc1041 (
      {stage0_24[101]},
      {stage1_24[99]}
   );
   gpc1_1 gpc1042 (
      {stage0_24[102]},
      {stage1_24[100]}
   );
   gpc1_1 gpc1043 (
      {stage0_24[103]},
      {stage1_24[101]}
   );
   gpc1_1 gpc1044 (
      {stage0_24[104]},
      {stage1_24[102]}
   );
   gpc1_1 gpc1045 (
      {stage0_24[105]},
      {stage1_24[103]}
   );
   gpc1_1 gpc1046 (
      {stage0_24[106]},
      {stage1_24[104]}
   );
   gpc1_1 gpc1047 (
      {stage0_24[107]},
      {stage1_24[105]}
   );
   gpc1_1 gpc1048 (
      {stage0_24[108]},
      {stage1_24[106]}
   );
   gpc1_1 gpc1049 (
      {stage0_24[109]},
      {stage1_24[107]}
   );
   gpc1_1 gpc1050 (
      {stage0_24[110]},
      {stage1_24[108]}
   );
   gpc1_1 gpc1051 (
      {stage0_24[111]},
      {stage1_24[109]}
   );
   gpc1_1 gpc1052 (
      {stage0_24[112]},
      {stage1_24[110]}
   );
   gpc1_1 gpc1053 (
      {stage0_24[113]},
      {stage1_24[111]}
   );
   gpc1_1 gpc1054 (
      {stage0_24[114]},
      {stage1_24[112]}
   );
   gpc1_1 gpc1055 (
      {stage0_24[115]},
      {stage1_24[113]}
   );
   gpc1_1 gpc1056 (
      {stage0_24[116]},
      {stage1_24[114]}
   );
   gpc1_1 gpc1057 (
      {stage0_24[117]},
      {stage1_24[115]}
   );
   gpc1_1 gpc1058 (
      {stage0_24[118]},
      {stage1_24[116]}
   );
   gpc1_1 gpc1059 (
      {stage0_24[119]},
      {stage1_24[117]}
   );
   gpc1_1 gpc1060 (
      {stage0_24[120]},
      {stage1_24[118]}
   );
   gpc1_1 gpc1061 (
      {stage0_24[121]},
      {stage1_24[119]}
   );
   gpc1_1 gpc1062 (
      {stage0_24[122]},
      {stage1_24[120]}
   );
   gpc1_1 gpc1063 (
      {stage0_24[123]},
      {stage1_24[121]}
   );
   gpc1_1 gpc1064 (
      {stage0_24[124]},
      {stage1_24[122]}
   );
   gpc1_1 gpc1065 (
      {stage0_24[125]},
      {stage1_24[123]}
   );
   gpc1_1 gpc1066 (
      {stage0_24[126]},
      {stage1_24[124]}
   );
   gpc1_1 gpc1067 (
      {stage0_24[127]},
      {stage1_24[125]}
   );
   gpc1_1 gpc1068 (
      {stage0_24[128]},
      {stage1_24[126]}
   );
   gpc1_1 gpc1069 (
      {stage0_24[129]},
      {stage1_24[127]}
   );
   gpc1_1 gpc1070 (
      {stage0_24[130]},
      {stage1_24[128]}
   );
   gpc1_1 gpc1071 (
      {stage0_24[131]},
      {stage1_24[129]}
   );
   gpc1_1 gpc1072 (
      {stage0_24[132]},
      {stage1_24[130]}
   );
   gpc1_1 gpc1073 (
      {stage0_24[133]},
      {stage1_24[131]}
   );
   gpc1_1 gpc1074 (
      {stage0_24[134]},
      {stage1_24[132]}
   );
   gpc1_1 gpc1075 (
      {stage0_24[135]},
      {stage1_24[133]}
   );
   gpc1_1 gpc1076 (
      {stage0_24[136]},
      {stage1_24[134]}
   );
   gpc1_1 gpc1077 (
      {stage0_24[137]},
      {stage1_24[135]}
   );
   gpc1_1 gpc1078 (
      {stage0_24[138]},
      {stage1_24[136]}
   );
   gpc1_1 gpc1079 (
      {stage0_24[139]},
      {stage1_24[137]}
   );
   gpc1_1 gpc1080 (
      {stage0_24[140]},
      {stage1_24[138]}
   );
   gpc1_1 gpc1081 (
      {stage0_24[141]},
      {stage1_24[139]}
   );
   gpc1_1 gpc1082 (
      {stage0_24[142]},
      {stage1_24[140]}
   );
   gpc1_1 gpc1083 (
      {stage0_24[143]},
      {stage1_24[141]}
   );
   gpc1_1 gpc1084 (
      {stage0_24[144]},
      {stage1_24[142]}
   );
   gpc1_1 gpc1085 (
      {stage0_24[145]},
      {stage1_24[143]}
   );
   gpc1_1 gpc1086 (
      {stage0_24[146]},
      {stage1_24[144]}
   );
   gpc1_1 gpc1087 (
      {stage0_24[147]},
      {stage1_24[145]}
   );
   gpc1_1 gpc1088 (
      {stage0_24[148]},
      {stage1_24[146]}
   );
   gpc1_1 gpc1089 (
      {stage0_24[149]},
      {stage1_24[147]}
   );
   gpc1_1 gpc1090 (
      {stage0_24[150]},
      {stage1_24[148]}
   );
   gpc1_1 gpc1091 (
      {stage0_24[151]},
      {stage1_24[149]}
   );
   gpc1_1 gpc1092 (
      {stage0_24[152]},
      {stage1_24[150]}
   );
   gpc1_1 gpc1093 (
      {stage0_24[153]},
      {stage1_24[151]}
   );
   gpc1_1 gpc1094 (
      {stage0_24[154]},
      {stage1_24[152]}
   );
   gpc1_1 gpc1095 (
      {stage0_24[155]},
      {stage1_24[153]}
   );
   gpc1_1 gpc1096 (
      {stage0_24[156]},
      {stage1_24[154]}
   );
   gpc1_1 gpc1097 (
      {stage0_24[157]},
      {stage1_24[155]}
   );
   gpc1_1 gpc1098 (
      {stage0_24[158]},
      {stage1_24[156]}
   );
   gpc1_1 gpc1099 (
      {stage0_24[159]},
      {stage1_24[157]}
   );
   gpc1_1 gpc1100 (
      {stage0_24[160]},
      {stage1_24[158]}
   );
   gpc1_1 gpc1101 (
      {stage0_24[161]},
      {stage1_24[159]}
   );
   gpc1_1 gpc1102 (
      {stage0_24[162]},
      {stage1_24[160]}
   );
   gpc1_1 gpc1103 (
      {stage0_24[163]},
      {stage1_24[161]}
   );
   gpc1_1 gpc1104 (
      {stage0_24[164]},
      {stage1_24[162]}
   );
   gpc1_1 gpc1105 (
      {stage0_24[165]},
      {stage1_24[163]}
   );
   gpc1_1 gpc1106 (
      {stage0_24[166]},
      {stage1_24[164]}
   );
   gpc1_1 gpc1107 (
      {stage0_24[167]},
      {stage1_24[165]}
   );
   gpc1_1 gpc1108 (
      {stage0_24[168]},
      {stage1_24[166]}
   );
   gpc1_1 gpc1109 (
      {stage0_24[169]},
      {stage1_24[167]}
   );
   gpc1_1 gpc1110 (
      {stage0_24[170]},
      {stage1_24[168]}
   );
   gpc1_1 gpc1111 (
      {stage0_24[171]},
      {stage1_24[169]}
   );
   gpc1_1 gpc1112 (
      {stage0_24[172]},
      {stage1_24[170]}
   );
   gpc1_1 gpc1113 (
      {stage0_24[173]},
      {stage1_24[171]}
   );
   gpc1_1 gpc1114 (
      {stage0_24[174]},
      {stage1_24[172]}
   );
   gpc1_1 gpc1115 (
      {stage0_24[175]},
      {stage1_24[173]}
   );
   gpc1_1 gpc1116 (
      {stage0_24[176]},
      {stage1_24[174]}
   );
   gpc1_1 gpc1117 (
      {stage0_24[177]},
      {stage1_24[175]}
   );
   gpc1_1 gpc1118 (
      {stage0_24[178]},
      {stage1_24[176]}
   );
   gpc1_1 gpc1119 (
      {stage0_24[179]},
      {stage1_24[177]}
   );
   gpc1_1 gpc1120 (
      {stage0_24[180]},
      {stage1_24[178]}
   );
   gpc1_1 gpc1121 (
      {stage0_24[181]},
      {stage1_24[179]}
   );
   gpc1_1 gpc1122 (
      {stage0_24[182]},
      {stage1_24[180]}
   );
   gpc1_1 gpc1123 (
      {stage0_24[183]},
      {stage1_24[181]}
   );
   gpc1_1 gpc1124 (
      {stage0_24[184]},
      {stage1_24[182]}
   );
   gpc1_1 gpc1125 (
      {stage0_24[185]},
      {stage1_24[183]}
   );
   gpc1_1 gpc1126 (
      {stage0_24[186]},
      {stage1_24[184]}
   );
   gpc1_1 gpc1127 (
      {stage0_24[187]},
      {stage1_24[185]}
   );
   gpc1_1 gpc1128 (
      {stage0_24[188]},
      {stage1_24[186]}
   );
   gpc1_1 gpc1129 (
      {stage0_24[189]},
      {stage1_24[187]}
   );
   gpc1_1 gpc1130 (
      {stage0_24[190]},
      {stage1_24[188]}
   );
   gpc1_1 gpc1131 (
      {stage0_24[191]},
      {stage1_24[189]}
   );
   gpc1_1 gpc1132 (
      {stage0_24[192]},
      {stage1_24[190]}
   );
   gpc1_1 gpc1133 (
      {stage0_24[193]},
      {stage1_24[191]}
   );
   gpc1_1 gpc1134 (
      {stage0_24[194]},
      {stage1_24[192]}
   );
   gpc1_1 gpc1135 (
      {stage0_24[195]},
      {stage1_24[193]}
   );
   gpc1_1 gpc1136 (
      {stage0_24[196]},
      {stage1_24[194]}
   );
   gpc1_1 gpc1137 (
      {stage0_24[197]},
      {stage1_24[195]}
   );
   gpc1_1 gpc1138 (
      {stage0_24[198]},
      {stage1_24[196]}
   );
   gpc1_1 gpc1139 (
      {stage0_24[199]},
      {stage1_24[197]}
   );
   gpc1_1 gpc1140 (
      {stage0_24[200]},
      {stage1_24[198]}
   );
   gpc1_1 gpc1141 (
      {stage0_24[201]},
      {stage1_24[199]}
   );
   gpc1_1 gpc1142 (
      {stage0_24[202]},
      {stage1_24[200]}
   );
   gpc1_1 gpc1143 (
      {stage0_24[203]},
      {stage1_24[201]}
   );
   gpc1_1 gpc1144 (
      {stage0_24[204]},
      {stage1_24[202]}
   );
   gpc1_1 gpc1145 (
      {stage0_24[205]},
      {stage1_24[203]}
   );
   gpc1_1 gpc1146 (
      {stage0_24[206]},
      {stage1_24[204]}
   );
   gpc1_1 gpc1147 (
      {stage0_24[207]},
      {stage1_24[205]}
   );
   gpc1_1 gpc1148 (
      {stage0_24[208]},
      {stage1_24[206]}
   );
   gpc1_1 gpc1149 (
      {stage0_24[209]},
      {stage1_24[207]}
   );
   gpc1_1 gpc1150 (
      {stage0_24[210]},
      {stage1_24[208]}
   );
   gpc1_1 gpc1151 (
      {stage0_24[211]},
      {stage1_24[209]}
   );
   gpc1_1 gpc1152 (
      {stage0_24[212]},
      {stage1_24[210]}
   );
   gpc1_1 gpc1153 (
      {stage0_24[213]},
      {stage1_24[211]}
   );
   gpc1_1 gpc1154 (
      {stage0_24[214]},
      {stage1_24[212]}
   );
   gpc1_1 gpc1155 (
      {stage0_24[215]},
      {stage1_24[213]}
   );
   gpc1_1 gpc1156 (
      {stage0_24[216]},
      {stage1_24[214]}
   );
   gpc1_1 gpc1157 (
      {stage0_24[217]},
      {stage1_24[215]}
   );
   gpc1_1 gpc1158 (
      {stage0_24[218]},
      {stage1_24[216]}
   );
   gpc1_1 gpc1159 (
      {stage0_24[219]},
      {stage1_24[217]}
   );
   gpc1_1 gpc1160 (
      {stage0_24[220]},
      {stage1_24[218]}
   );
   gpc1_1 gpc1161 (
      {stage0_24[221]},
      {stage1_24[219]}
   );
   gpc1_1 gpc1162 (
      {stage0_24[222]},
      {stage1_24[220]}
   );
   gpc1_1 gpc1163 (
      {stage0_24[223]},
      {stage1_24[221]}
   );
   gpc1_1 gpc1164 (
      {stage0_24[224]},
      {stage1_24[222]}
   );
   gpc1_1 gpc1165 (
      {stage0_24[225]},
      {stage1_24[223]}
   );
   gpc1_1 gpc1166 (
      {stage0_24[226]},
      {stage1_24[224]}
   );
   gpc1_1 gpc1167 (
      {stage0_24[227]},
      {stage1_24[225]}
   );
   gpc1_1 gpc1168 (
      {stage0_24[228]},
      {stage1_24[226]}
   );
   gpc1_1 gpc1169 (
      {stage0_24[229]},
      {stage1_24[227]}
   );
   gpc1_1 gpc1170 (
      {stage0_24[230]},
      {stage1_24[228]}
   );
   gpc1_1 gpc1171 (
      {stage0_24[231]},
      {stage1_24[229]}
   );
   gpc1_1 gpc1172 (
      {stage0_24[232]},
      {stage1_24[230]}
   );
   gpc1_1 gpc1173 (
      {stage0_24[233]},
      {stage1_24[231]}
   );
   gpc1_1 gpc1174 (
      {stage0_24[234]},
      {stage1_24[232]}
   );
   gpc1_1 gpc1175 (
      {stage0_24[235]},
      {stage1_24[233]}
   );
   gpc1_1 gpc1176 (
      {stage0_24[236]},
      {stage1_24[234]}
   );
   gpc1_1 gpc1177 (
      {stage0_24[237]},
      {stage1_24[235]}
   );
   gpc1_1 gpc1178 (
      {stage0_24[238]},
      {stage1_24[236]}
   );
   gpc1_1 gpc1179 (
      {stage0_24[239]},
      {stage1_24[237]}
   );
   gpc1_1 gpc1180 (
      {stage0_24[240]},
      {stage1_24[238]}
   );
   gpc1_1 gpc1181 (
      {stage0_24[241]},
      {stage1_24[239]}
   );
   gpc1_1 gpc1182 (
      {stage0_24[242]},
      {stage1_24[240]}
   );
   gpc1_1 gpc1183 (
      {stage0_24[243]},
      {stage1_24[241]}
   );
   gpc1_1 gpc1184 (
      {stage0_24[244]},
      {stage1_24[242]}
   );
   gpc1_1 gpc1185 (
      {stage0_24[245]},
      {stage1_24[243]}
   );
   gpc1_1 gpc1186 (
      {stage0_24[246]},
      {stage1_24[244]}
   );
   gpc1_1 gpc1187 (
      {stage0_24[247]},
      {stage1_24[245]}
   );
   gpc1_1 gpc1188 (
      {stage0_24[248]},
      {stage1_24[246]}
   );
   gpc1_1 gpc1189 (
      {stage0_24[249]},
      {stage1_24[247]}
   );
   gpc1_1 gpc1190 (
      {stage0_24[250]},
      {stage1_24[248]}
   );
   gpc1_1 gpc1191 (
      {stage0_24[251]},
      {stage1_24[249]}
   );
   gpc1_1 gpc1192 (
      {stage0_24[252]},
      {stage1_24[250]}
   );
   gpc1_1 gpc1193 (
      {stage0_24[253]},
      {stage1_24[251]}
   );
   gpc1_1 gpc1194 (
      {stage0_24[254]},
      {stage1_24[252]}
   );
   gpc1_1 gpc1195 (
      {stage0_24[255]},
      {stage1_24[253]}
   );
   gpc1_1 gpc1196 (
      {stage0_25[222]},
      {stage1_25[84]}
   );
   gpc1_1 gpc1197 (
      {stage0_25[223]},
      {stage1_25[85]}
   );
   gpc1_1 gpc1198 (
      {stage0_25[224]},
      {stage1_25[86]}
   );
   gpc1_1 gpc1199 (
      {stage0_25[225]},
      {stage1_25[87]}
   );
   gpc1_1 gpc1200 (
      {stage0_25[226]},
      {stage1_25[88]}
   );
   gpc1_1 gpc1201 (
      {stage0_25[227]},
      {stage1_25[89]}
   );
   gpc1_1 gpc1202 (
      {stage0_25[228]},
      {stage1_25[90]}
   );
   gpc1_1 gpc1203 (
      {stage0_25[229]},
      {stage1_25[91]}
   );
   gpc1_1 gpc1204 (
      {stage0_25[230]},
      {stage1_25[92]}
   );
   gpc1_1 gpc1205 (
      {stage0_25[231]},
      {stage1_25[93]}
   );
   gpc1_1 gpc1206 (
      {stage0_25[232]},
      {stage1_25[94]}
   );
   gpc1_1 gpc1207 (
      {stage0_25[233]},
      {stage1_25[95]}
   );
   gpc1_1 gpc1208 (
      {stage0_25[234]},
      {stage1_25[96]}
   );
   gpc1_1 gpc1209 (
      {stage0_25[235]},
      {stage1_25[97]}
   );
   gpc1_1 gpc1210 (
      {stage0_25[236]},
      {stage1_25[98]}
   );
   gpc1_1 gpc1211 (
      {stage0_25[237]},
      {stage1_25[99]}
   );
   gpc1_1 gpc1212 (
      {stage0_25[238]},
      {stage1_25[100]}
   );
   gpc1_1 gpc1213 (
      {stage0_25[239]},
      {stage1_25[101]}
   );
   gpc1_1 gpc1214 (
      {stage0_25[240]},
      {stage1_25[102]}
   );
   gpc1_1 gpc1215 (
      {stage0_25[241]},
      {stage1_25[103]}
   );
   gpc1_1 gpc1216 (
      {stage0_25[242]},
      {stage1_25[104]}
   );
   gpc1_1 gpc1217 (
      {stage0_25[243]},
      {stage1_25[105]}
   );
   gpc1_1 gpc1218 (
      {stage0_25[244]},
      {stage1_25[106]}
   );
   gpc1_1 gpc1219 (
      {stage0_25[245]},
      {stage1_25[107]}
   );
   gpc1_1 gpc1220 (
      {stage0_25[246]},
      {stage1_25[108]}
   );
   gpc1_1 gpc1221 (
      {stage0_25[247]},
      {stage1_25[109]}
   );
   gpc1_1 gpc1222 (
      {stage0_25[248]},
      {stage1_25[110]}
   );
   gpc1_1 gpc1223 (
      {stage0_25[249]},
      {stage1_25[111]}
   );
   gpc1_1 gpc1224 (
      {stage0_25[250]},
      {stage1_25[112]}
   );
   gpc1_1 gpc1225 (
      {stage0_25[251]},
      {stage1_25[113]}
   );
   gpc1_1 gpc1226 (
      {stage0_25[252]},
      {stage1_25[114]}
   );
   gpc1_1 gpc1227 (
      {stage0_25[253]},
      {stage1_25[115]}
   );
   gpc1_1 gpc1228 (
      {stage0_25[254]},
      {stage1_25[116]}
   );
   gpc1_1 gpc1229 (
      {stage0_25[255]},
      {stage1_25[117]}
   );
   gpc1_1 gpc1230 (
      {stage0_26[72]},
      {stage1_26[53]}
   );
   gpc1_1 gpc1231 (
      {stage0_26[73]},
      {stage1_26[54]}
   );
   gpc1_1 gpc1232 (
      {stage0_26[74]},
      {stage1_26[55]}
   );
   gpc1_1 gpc1233 (
      {stage0_26[75]},
      {stage1_26[56]}
   );
   gpc1_1 gpc1234 (
      {stage0_26[76]},
      {stage1_26[57]}
   );
   gpc1_1 gpc1235 (
      {stage0_26[77]},
      {stage1_26[58]}
   );
   gpc1_1 gpc1236 (
      {stage0_26[78]},
      {stage1_26[59]}
   );
   gpc1_1 gpc1237 (
      {stage0_26[79]},
      {stage1_26[60]}
   );
   gpc1_1 gpc1238 (
      {stage0_26[80]},
      {stage1_26[61]}
   );
   gpc1_1 gpc1239 (
      {stage0_26[81]},
      {stage1_26[62]}
   );
   gpc1_1 gpc1240 (
      {stage0_26[82]},
      {stage1_26[63]}
   );
   gpc1_1 gpc1241 (
      {stage0_26[83]},
      {stage1_26[64]}
   );
   gpc1_1 gpc1242 (
      {stage0_26[84]},
      {stage1_26[65]}
   );
   gpc1_1 gpc1243 (
      {stage0_26[85]},
      {stage1_26[66]}
   );
   gpc1_1 gpc1244 (
      {stage0_26[86]},
      {stage1_26[67]}
   );
   gpc1_1 gpc1245 (
      {stage0_26[87]},
      {stage1_26[68]}
   );
   gpc1_1 gpc1246 (
      {stage0_26[88]},
      {stage1_26[69]}
   );
   gpc1_1 gpc1247 (
      {stage0_26[89]},
      {stage1_26[70]}
   );
   gpc1_1 gpc1248 (
      {stage0_26[90]},
      {stage1_26[71]}
   );
   gpc1_1 gpc1249 (
      {stage0_26[91]},
      {stage1_26[72]}
   );
   gpc1_1 gpc1250 (
      {stage0_26[92]},
      {stage1_26[73]}
   );
   gpc1_1 gpc1251 (
      {stage0_26[93]},
      {stage1_26[74]}
   );
   gpc1_1 gpc1252 (
      {stage0_26[94]},
      {stage1_26[75]}
   );
   gpc1_1 gpc1253 (
      {stage0_26[95]},
      {stage1_26[76]}
   );
   gpc1_1 gpc1254 (
      {stage0_26[96]},
      {stage1_26[77]}
   );
   gpc1_1 gpc1255 (
      {stage0_26[97]},
      {stage1_26[78]}
   );
   gpc1_1 gpc1256 (
      {stage0_26[98]},
      {stage1_26[79]}
   );
   gpc1_1 gpc1257 (
      {stage0_26[99]},
      {stage1_26[80]}
   );
   gpc1_1 gpc1258 (
      {stage0_26[100]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1259 (
      {stage0_26[101]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1260 (
      {stage0_26[102]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1261 (
      {stage0_26[103]},
      {stage1_26[84]}
   );
   gpc1_1 gpc1262 (
      {stage0_26[104]},
      {stage1_26[85]}
   );
   gpc1_1 gpc1263 (
      {stage0_26[105]},
      {stage1_26[86]}
   );
   gpc1_1 gpc1264 (
      {stage0_26[106]},
      {stage1_26[87]}
   );
   gpc1_1 gpc1265 (
      {stage0_26[107]},
      {stage1_26[88]}
   );
   gpc1_1 gpc1266 (
      {stage0_26[108]},
      {stage1_26[89]}
   );
   gpc1_1 gpc1267 (
      {stage0_26[109]},
      {stage1_26[90]}
   );
   gpc1_1 gpc1268 (
      {stage0_26[110]},
      {stage1_26[91]}
   );
   gpc1_1 gpc1269 (
      {stage0_26[111]},
      {stage1_26[92]}
   );
   gpc1_1 gpc1270 (
      {stage0_26[112]},
      {stage1_26[93]}
   );
   gpc1_1 gpc1271 (
      {stage0_26[113]},
      {stage1_26[94]}
   );
   gpc1_1 gpc1272 (
      {stage0_26[114]},
      {stage1_26[95]}
   );
   gpc1_1 gpc1273 (
      {stage0_26[115]},
      {stage1_26[96]}
   );
   gpc1_1 gpc1274 (
      {stage0_26[116]},
      {stage1_26[97]}
   );
   gpc1_1 gpc1275 (
      {stage0_26[117]},
      {stage1_26[98]}
   );
   gpc1_1 gpc1276 (
      {stage0_26[118]},
      {stage1_26[99]}
   );
   gpc1_1 gpc1277 (
      {stage0_26[119]},
      {stage1_26[100]}
   );
   gpc1_1 gpc1278 (
      {stage0_26[120]},
      {stage1_26[101]}
   );
   gpc1_1 gpc1279 (
      {stage0_26[121]},
      {stage1_26[102]}
   );
   gpc1_1 gpc1280 (
      {stage0_26[122]},
      {stage1_26[103]}
   );
   gpc1_1 gpc1281 (
      {stage0_26[123]},
      {stage1_26[104]}
   );
   gpc1_1 gpc1282 (
      {stage0_26[124]},
      {stage1_26[105]}
   );
   gpc1_1 gpc1283 (
      {stage0_26[125]},
      {stage1_26[106]}
   );
   gpc1_1 gpc1284 (
      {stage0_26[126]},
      {stage1_26[107]}
   );
   gpc1_1 gpc1285 (
      {stage0_26[127]},
      {stage1_26[108]}
   );
   gpc1_1 gpc1286 (
      {stage0_26[128]},
      {stage1_26[109]}
   );
   gpc1_1 gpc1287 (
      {stage0_26[129]},
      {stage1_26[110]}
   );
   gpc1_1 gpc1288 (
      {stage0_26[130]},
      {stage1_26[111]}
   );
   gpc1_1 gpc1289 (
      {stage0_26[131]},
      {stage1_26[112]}
   );
   gpc1_1 gpc1290 (
      {stage0_26[132]},
      {stage1_26[113]}
   );
   gpc1_1 gpc1291 (
      {stage0_26[133]},
      {stage1_26[114]}
   );
   gpc1_1 gpc1292 (
      {stage0_26[134]},
      {stage1_26[115]}
   );
   gpc1_1 gpc1293 (
      {stage0_26[135]},
      {stage1_26[116]}
   );
   gpc1_1 gpc1294 (
      {stage0_26[136]},
      {stage1_26[117]}
   );
   gpc1_1 gpc1295 (
      {stage0_26[137]},
      {stage1_26[118]}
   );
   gpc1_1 gpc1296 (
      {stage0_26[138]},
      {stage1_26[119]}
   );
   gpc1_1 gpc1297 (
      {stage0_26[139]},
      {stage1_26[120]}
   );
   gpc1_1 gpc1298 (
      {stage0_26[140]},
      {stage1_26[121]}
   );
   gpc1_1 gpc1299 (
      {stage0_26[141]},
      {stage1_26[122]}
   );
   gpc1_1 gpc1300 (
      {stage0_26[142]},
      {stage1_26[123]}
   );
   gpc1_1 gpc1301 (
      {stage0_26[143]},
      {stage1_26[124]}
   );
   gpc1_1 gpc1302 (
      {stage0_26[144]},
      {stage1_26[125]}
   );
   gpc1_1 gpc1303 (
      {stage0_26[145]},
      {stage1_26[126]}
   );
   gpc1_1 gpc1304 (
      {stage0_26[146]},
      {stage1_26[127]}
   );
   gpc1_1 gpc1305 (
      {stage0_26[147]},
      {stage1_26[128]}
   );
   gpc1_1 gpc1306 (
      {stage0_26[148]},
      {stage1_26[129]}
   );
   gpc1_1 gpc1307 (
      {stage0_26[149]},
      {stage1_26[130]}
   );
   gpc1_1 gpc1308 (
      {stage0_26[150]},
      {stage1_26[131]}
   );
   gpc1_1 gpc1309 (
      {stage0_26[151]},
      {stage1_26[132]}
   );
   gpc1_1 gpc1310 (
      {stage0_26[152]},
      {stage1_26[133]}
   );
   gpc1_1 gpc1311 (
      {stage0_26[153]},
      {stage1_26[134]}
   );
   gpc1_1 gpc1312 (
      {stage0_26[154]},
      {stage1_26[135]}
   );
   gpc1_1 gpc1313 (
      {stage0_26[155]},
      {stage1_26[136]}
   );
   gpc1_1 gpc1314 (
      {stage0_26[156]},
      {stage1_26[137]}
   );
   gpc1_1 gpc1315 (
      {stage0_26[157]},
      {stage1_26[138]}
   );
   gpc1_1 gpc1316 (
      {stage0_26[158]},
      {stage1_26[139]}
   );
   gpc1_1 gpc1317 (
      {stage0_26[159]},
      {stage1_26[140]}
   );
   gpc1_1 gpc1318 (
      {stage0_26[160]},
      {stage1_26[141]}
   );
   gpc1_1 gpc1319 (
      {stage0_26[161]},
      {stage1_26[142]}
   );
   gpc1_1 gpc1320 (
      {stage0_26[162]},
      {stage1_26[143]}
   );
   gpc1_1 gpc1321 (
      {stage0_26[163]},
      {stage1_26[144]}
   );
   gpc1_1 gpc1322 (
      {stage0_26[164]},
      {stage1_26[145]}
   );
   gpc1_1 gpc1323 (
      {stage0_26[165]},
      {stage1_26[146]}
   );
   gpc1_1 gpc1324 (
      {stage0_26[166]},
      {stage1_26[147]}
   );
   gpc1_1 gpc1325 (
      {stage0_26[167]},
      {stage1_26[148]}
   );
   gpc1_1 gpc1326 (
      {stage0_26[168]},
      {stage1_26[149]}
   );
   gpc1_1 gpc1327 (
      {stage0_26[169]},
      {stage1_26[150]}
   );
   gpc1_1 gpc1328 (
      {stage0_26[170]},
      {stage1_26[151]}
   );
   gpc1_1 gpc1329 (
      {stage0_26[171]},
      {stage1_26[152]}
   );
   gpc1_1 gpc1330 (
      {stage0_26[172]},
      {stage1_26[153]}
   );
   gpc1_1 gpc1331 (
      {stage0_26[173]},
      {stage1_26[154]}
   );
   gpc1_1 gpc1332 (
      {stage0_26[174]},
      {stage1_26[155]}
   );
   gpc1_1 gpc1333 (
      {stage0_26[175]},
      {stage1_26[156]}
   );
   gpc1_1 gpc1334 (
      {stage0_26[176]},
      {stage1_26[157]}
   );
   gpc1_1 gpc1335 (
      {stage0_26[177]},
      {stage1_26[158]}
   );
   gpc1_1 gpc1336 (
      {stage0_26[178]},
      {stage1_26[159]}
   );
   gpc1_1 gpc1337 (
      {stage0_26[179]},
      {stage1_26[160]}
   );
   gpc1_1 gpc1338 (
      {stage0_26[180]},
      {stage1_26[161]}
   );
   gpc1_1 gpc1339 (
      {stage0_26[181]},
      {stage1_26[162]}
   );
   gpc1_1 gpc1340 (
      {stage0_26[182]},
      {stage1_26[163]}
   );
   gpc1_1 gpc1341 (
      {stage0_26[183]},
      {stage1_26[164]}
   );
   gpc1_1 gpc1342 (
      {stage0_26[184]},
      {stage1_26[165]}
   );
   gpc1_1 gpc1343 (
      {stage0_26[185]},
      {stage1_26[166]}
   );
   gpc1_1 gpc1344 (
      {stage0_26[186]},
      {stage1_26[167]}
   );
   gpc1_1 gpc1345 (
      {stage0_26[187]},
      {stage1_26[168]}
   );
   gpc1_1 gpc1346 (
      {stage0_26[188]},
      {stage1_26[169]}
   );
   gpc1_1 gpc1347 (
      {stage0_26[189]},
      {stage1_26[170]}
   );
   gpc1_1 gpc1348 (
      {stage0_26[190]},
      {stage1_26[171]}
   );
   gpc1_1 gpc1349 (
      {stage0_26[191]},
      {stage1_26[172]}
   );
   gpc1_1 gpc1350 (
      {stage0_26[192]},
      {stage1_26[173]}
   );
   gpc1_1 gpc1351 (
      {stage0_26[193]},
      {stage1_26[174]}
   );
   gpc1_1 gpc1352 (
      {stage0_26[194]},
      {stage1_26[175]}
   );
   gpc1_1 gpc1353 (
      {stage0_26[195]},
      {stage1_26[176]}
   );
   gpc1_1 gpc1354 (
      {stage0_26[196]},
      {stage1_26[177]}
   );
   gpc1_1 gpc1355 (
      {stage0_26[197]},
      {stage1_26[178]}
   );
   gpc1_1 gpc1356 (
      {stage0_26[198]},
      {stage1_26[179]}
   );
   gpc1_1 gpc1357 (
      {stage0_26[199]},
      {stage1_26[180]}
   );
   gpc1_1 gpc1358 (
      {stage0_26[200]},
      {stage1_26[181]}
   );
   gpc1_1 gpc1359 (
      {stage0_26[201]},
      {stage1_26[182]}
   );
   gpc1_1 gpc1360 (
      {stage0_26[202]},
      {stage1_26[183]}
   );
   gpc1_1 gpc1361 (
      {stage0_26[203]},
      {stage1_26[184]}
   );
   gpc1_1 gpc1362 (
      {stage0_26[204]},
      {stage1_26[185]}
   );
   gpc1_1 gpc1363 (
      {stage0_26[205]},
      {stage1_26[186]}
   );
   gpc1_1 gpc1364 (
      {stage0_26[206]},
      {stage1_26[187]}
   );
   gpc1_1 gpc1365 (
      {stage0_26[207]},
      {stage1_26[188]}
   );
   gpc1_1 gpc1366 (
      {stage0_26[208]},
      {stage1_26[189]}
   );
   gpc1_1 gpc1367 (
      {stage0_26[209]},
      {stage1_26[190]}
   );
   gpc1_1 gpc1368 (
      {stage0_26[210]},
      {stage1_26[191]}
   );
   gpc1_1 gpc1369 (
      {stage0_26[211]},
      {stage1_26[192]}
   );
   gpc1_1 gpc1370 (
      {stage0_26[212]},
      {stage1_26[193]}
   );
   gpc1_1 gpc1371 (
      {stage0_26[213]},
      {stage1_26[194]}
   );
   gpc1_1 gpc1372 (
      {stage0_26[214]},
      {stage1_26[195]}
   );
   gpc1_1 gpc1373 (
      {stage0_26[215]},
      {stage1_26[196]}
   );
   gpc1_1 gpc1374 (
      {stage0_26[216]},
      {stage1_26[197]}
   );
   gpc1_1 gpc1375 (
      {stage0_26[217]},
      {stage1_26[198]}
   );
   gpc1_1 gpc1376 (
      {stage0_26[218]},
      {stage1_26[199]}
   );
   gpc1_1 gpc1377 (
      {stage0_26[219]},
      {stage1_26[200]}
   );
   gpc1_1 gpc1378 (
      {stage0_26[220]},
      {stage1_26[201]}
   );
   gpc1_1 gpc1379 (
      {stage0_26[221]},
      {stage1_26[202]}
   );
   gpc1_1 gpc1380 (
      {stage0_26[222]},
      {stage1_26[203]}
   );
   gpc1_1 gpc1381 (
      {stage0_26[223]},
      {stage1_26[204]}
   );
   gpc1_1 gpc1382 (
      {stage0_26[224]},
      {stage1_26[205]}
   );
   gpc1_1 gpc1383 (
      {stage0_26[225]},
      {stage1_26[206]}
   );
   gpc1_1 gpc1384 (
      {stage0_26[226]},
      {stage1_26[207]}
   );
   gpc1_1 gpc1385 (
      {stage0_26[227]},
      {stage1_26[208]}
   );
   gpc1_1 gpc1386 (
      {stage0_26[228]},
      {stage1_26[209]}
   );
   gpc1_1 gpc1387 (
      {stage0_26[229]},
      {stage1_26[210]}
   );
   gpc1_1 gpc1388 (
      {stage0_26[230]},
      {stage1_26[211]}
   );
   gpc1_1 gpc1389 (
      {stage0_26[231]},
      {stage1_26[212]}
   );
   gpc1_1 gpc1390 (
      {stage0_26[232]},
      {stage1_26[213]}
   );
   gpc1_1 gpc1391 (
      {stage0_26[233]},
      {stage1_26[214]}
   );
   gpc1_1 gpc1392 (
      {stage0_26[234]},
      {stage1_26[215]}
   );
   gpc1_1 gpc1393 (
      {stage0_26[235]},
      {stage1_26[216]}
   );
   gpc1_1 gpc1394 (
      {stage0_26[236]},
      {stage1_26[217]}
   );
   gpc1_1 gpc1395 (
      {stage0_26[237]},
      {stage1_26[218]}
   );
   gpc1_1 gpc1396 (
      {stage0_26[238]},
      {stage1_26[219]}
   );
   gpc1_1 gpc1397 (
      {stage0_26[239]},
      {stage1_26[220]}
   );
   gpc1_1 gpc1398 (
      {stage0_26[240]},
      {stage1_26[221]}
   );
   gpc1_1 gpc1399 (
      {stage0_26[241]},
      {stage1_26[222]}
   );
   gpc1_1 gpc1400 (
      {stage0_26[242]},
      {stage1_26[223]}
   );
   gpc1_1 gpc1401 (
      {stage0_26[243]},
      {stage1_26[224]}
   );
   gpc1_1 gpc1402 (
      {stage0_26[244]},
      {stage1_26[225]}
   );
   gpc1_1 gpc1403 (
      {stage0_26[245]},
      {stage1_26[226]}
   );
   gpc1_1 gpc1404 (
      {stage0_26[246]},
      {stage1_26[227]}
   );
   gpc1_1 gpc1405 (
      {stage0_26[247]},
      {stage1_26[228]}
   );
   gpc1_1 gpc1406 (
      {stage0_26[248]},
      {stage1_26[229]}
   );
   gpc1_1 gpc1407 (
      {stage0_26[249]},
      {stage1_26[230]}
   );
   gpc1_1 gpc1408 (
      {stage0_26[250]},
      {stage1_26[231]}
   );
   gpc1_1 gpc1409 (
      {stage0_26[251]},
      {stage1_26[232]}
   );
   gpc1_1 gpc1410 (
      {stage0_26[252]},
      {stage1_26[233]}
   );
   gpc1_1 gpc1411 (
      {stage0_26[253]},
      {stage1_26[234]}
   );
   gpc1_1 gpc1412 (
      {stage0_26[254]},
      {stage1_26[235]}
   );
   gpc1_1 gpc1413 (
      {stage0_26[255]},
      {stage1_26[236]}
   );
   gpc1_1 gpc1414 (
      {stage0_27[204]},
      {stage1_27[56]}
   );
   gpc1_1 gpc1415 (
      {stage0_27[205]},
      {stage1_27[57]}
   );
   gpc1_1 gpc1416 (
      {stage0_27[206]},
      {stage1_27[58]}
   );
   gpc1_1 gpc1417 (
      {stage0_27[207]},
      {stage1_27[59]}
   );
   gpc1_1 gpc1418 (
      {stage0_27[208]},
      {stage1_27[60]}
   );
   gpc1_1 gpc1419 (
      {stage0_27[209]},
      {stage1_27[61]}
   );
   gpc1_1 gpc1420 (
      {stage0_27[210]},
      {stage1_27[62]}
   );
   gpc1_1 gpc1421 (
      {stage0_27[211]},
      {stage1_27[63]}
   );
   gpc1_1 gpc1422 (
      {stage0_27[212]},
      {stage1_27[64]}
   );
   gpc1_1 gpc1423 (
      {stage0_27[213]},
      {stage1_27[65]}
   );
   gpc1_1 gpc1424 (
      {stage0_27[214]},
      {stage1_27[66]}
   );
   gpc1_1 gpc1425 (
      {stage0_27[215]},
      {stage1_27[67]}
   );
   gpc1_1 gpc1426 (
      {stage0_27[216]},
      {stage1_27[68]}
   );
   gpc1_1 gpc1427 (
      {stage0_27[217]},
      {stage1_27[69]}
   );
   gpc1_1 gpc1428 (
      {stage0_27[218]},
      {stage1_27[70]}
   );
   gpc1_1 gpc1429 (
      {stage0_27[219]},
      {stage1_27[71]}
   );
   gpc1_1 gpc1430 (
      {stage0_27[220]},
      {stage1_27[72]}
   );
   gpc1_1 gpc1431 (
      {stage0_27[221]},
      {stage1_27[73]}
   );
   gpc1_1 gpc1432 (
      {stage0_27[222]},
      {stage1_27[74]}
   );
   gpc1_1 gpc1433 (
      {stage0_27[223]},
      {stage1_27[75]}
   );
   gpc1_1 gpc1434 (
      {stage0_27[224]},
      {stage1_27[76]}
   );
   gpc1_1 gpc1435 (
      {stage0_27[225]},
      {stage1_27[77]}
   );
   gpc1_1 gpc1436 (
      {stage0_27[226]},
      {stage1_27[78]}
   );
   gpc1_1 gpc1437 (
      {stage0_27[227]},
      {stage1_27[79]}
   );
   gpc1_1 gpc1438 (
      {stage0_27[228]},
      {stage1_27[80]}
   );
   gpc1_1 gpc1439 (
      {stage0_27[229]},
      {stage1_27[81]}
   );
   gpc1_1 gpc1440 (
      {stage0_27[230]},
      {stage1_27[82]}
   );
   gpc1_1 gpc1441 (
      {stage0_27[231]},
      {stage1_27[83]}
   );
   gpc1_1 gpc1442 (
      {stage0_27[232]},
      {stage1_27[84]}
   );
   gpc1_1 gpc1443 (
      {stage0_27[233]},
      {stage1_27[85]}
   );
   gpc1_1 gpc1444 (
      {stage0_27[234]},
      {stage1_27[86]}
   );
   gpc1_1 gpc1445 (
      {stage0_27[235]},
      {stage1_27[87]}
   );
   gpc1_1 gpc1446 (
      {stage0_27[236]},
      {stage1_27[88]}
   );
   gpc1_1 gpc1447 (
      {stage0_27[237]},
      {stage1_27[89]}
   );
   gpc1_1 gpc1448 (
      {stage0_27[238]},
      {stage1_27[90]}
   );
   gpc1_1 gpc1449 (
      {stage0_27[239]},
      {stage1_27[91]}
   );
   gpc1_1 gpc1450 (
      {stage0_27[240]},
      {stage1_27[92]}
   );
   gpc1_1 gpc1451 (
      {stage0_27[241]},
      {stage1_27[93]}
   );
   gpc1_1 gpc1452 (
      {stage0_27[242]},
      {stage1_27[94]}
   );
   gpc1_1 gpc1453 (
      {stage0_27[243]},
      {stage1_27[95]}
   );
   gpc1_1 gpc1454 (
      {stage0_27[244]},
      {stage1_27[96]}
   );
   gpc1_1 gpc1455 (
      {stage0_27[245]},
      {stage1_27[97]}
   );
   gpc1_1 gpc1456 (
      {stage0_27[246]},
      {stage1_27[98]}
   );
   gpc1_1 gpc1457 (
      {stage0_27[247]},
      {stage1_27[99]}
   );
   gpc1_1 gpc1458 (
      {stage0_27[248]},
      {stage1_27[100]}
   );
   gpc1_1 gpc1459 (
      {stage0_27[249]},
      {stage1_27[101]}
   );
   gpc1_1 gpc1460 (
      {stage0_27[250]},
      {stage1_27[102]}
   );
   gpc1_1 gpc1461 (
      {stage0_27[251]},
      {stage1_27[103]}
   );
   gpc1_1 gpc1462 (
      {stage0_27[252]},
      {stage1_27[104]}
   );
   gpc1_1 gpc1463 (
      {stage0_27[253]},
      {stage1_27[105]}
   );
   gpc1_1 gpc1464 (
      {stage0_27[254]},
      {stage1_27[106]}
   );
   gpc1_1 gpc1465 (
      {stage0_27[255]},
      {stage1_27[107]}
   );
   gpc1_1 gpc1466 (
      {stage0_28[240]},
      {stage1_28[86]}
   );
   gpc1_1 gpc1467 (
      {stage0_28[241]},
      {stage1_28[87]}
   );
   gpc1_1 gpc1468 (
      {stage0_28[242]},
      {stage1_28[88]}
   );
   gpc1_1 gpc1469 (
      {stage0_28[243]},
      {stage1_28[89]}
   );
   gpc1_1 gpc1470 (
      {stage0_28[244]},
      {stage1_28[90]}
   );
   gpc1_1 gpc1471 (
      {stage0_28[245]},
      {stage1_28[91]}
   );
   gpc1_1 gpc1472 (
      {stage0_28[246]},
      {stage1_28[92]}
   );
   gpc1_1 gpc1473 (
      {stage0_28[247]},
      {stage1_28[93]}
   );
   gpc1_1 gpc1474 (
      {stage0_28[248]},
      {stage1_28[94]}
   );
   gpc1_1 gpc1475 (
      {stage0_28[249]},
      {stage1_28[95]}
   );
   gpc1_1 gpc1476 (
      {stage0_28[250]},
      {stage1_28[96]}
   );
   gpc1_1 gpc1477 (
      {stage0_28[251]},
      {stage1_28[97]}
   );
   gpc1_1 gpc1478 (
      {stage0_28[252]},
      {stage1_28[98]}
   );
   gpc1_1 gpc1479 (
      {stage0_28[253]},
      {stage1_28[99]}
   );
   gpc1_1 gpc1480 (
      {stage0_28[254]},
      {stage1_28[100]}
   );
   gpc1_1 gpc1481 (
      {stage0_28[255]},
      {stage1_28[101]}
   );
   gpc1_1 gpc1482 (
      {stage0_29[246]},
      {stage1_29[108]}
   );
   gpc1_1 gpc1483 (
      {stage0_29[247]},
      {stage1_29[109]}
   );
   gpc1_1 gpc1484 (
      {stage0_29[248]},
      {stage1_29[110]}
   );
   gpc1_1 gpc1485 (
      {stage0_29[249]},
      {stage1_29[111]}
   );
   gpc1_1 gpc1486 (
      {stage0_29[250]},
      {stage1_29[112]}
   );
   gpc1_1 gpc1487 (
      {stage0_29[251]},
      {stage1_29[113]}
   );
   gpc1_1 gpc1488 (
      {stage0_29[252]},
      {stage1_29[114]}
   );
   gpc1_1 gpc1489 (
      {stage0_29[253]},
      {stage1_29[115]}
   );
   gpc1_1 gpc1490 (
      {stage0_29[254]},
      {stage1_29[116]}
   );
   gpc1_1 gpc1491 (
      {stage0_29[255]},
      {stage1_29[117]}
   );
   gpc1_1 gpc1492 (
      {stage0_30[240]},
      {stage1_30[81]}
   );
   gpc1_1 gpc1493 (
      {stage0_30[241]},
      {stage1_30[82]}
   );
   gpc1_1 gpc1494 (
      {stage0_30[242]},
      {stage1_30[83]}
   );
   gpc1_1 gpc1495 (
      {stage0_30[243]},
      {stage1_30[84]}
   );
   gpc1_1 gpc1496 (
      {stage0_30[244]},
      {stage1_30[85]}
   );
   gpc1_1 gpc1497 (
      {stage0_30[245]},
      {stage1_30[86]}
   );
   gpc1_1 gpc1498 (
      {stage0_30[246]},
      {stage1_30[87]}
   );
   gpc1_1 gpc1499 (
      {stage0_30[247]},
      {stage1_30[88]}
   );
   gpc1_1 gpc1500 (
      {stage0_30[248]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1501 (
      {stage0_30[249]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1502 (
      {stage0_30[250]},
      {stage1_30[91]}
   );
   gpc1_1 gpc1503 (
      {stage0_30[251]},
      {stage1_30[92]}
   );
   gpc1_1 gpc1504 (
      {stage0_30[252]},
      {stage1_30[93]}
   );
   gpc1_1 gpc1505 (
      {stage0_30[253]},
      {stage1_30[94]}
   );
   gpc1_1 gpc1506 (
      {stage0_30[254]},
      {stage1_30[95]}
   );
   gpc1_1 gpc1507 (
      {stage0_30[255]},
      {stage1_30[96]}
   );
   gpc1_1 gpc1508 (
      {stage0_31[204]},
      {stage1_31[81]}
   );
   gpc1_1 gpc1509 (
      {stage0_31[205]},
      {stage1_31[82]}
   );
   gpc1_1 gpc1510 (
      {stage0_31[206]},
      {stage1_31[83]}
   );
   gpc1_1 gpc1511 (
      {stage0_31[207]},
      {stage1_31[84]}
   );
   gpc1_1 gpc1512 (
      {stage0_31[208]},
      {stage1_31[85]}
   );
   gpc1_1 gpc1513 (
      {stage0_31[209]},
      {stage1_31[86]}
   );
   gpc1_1 gpc1514 (
      {stage0_31[210]},
      {stage1_31[87]}
   );
   gpc1_1 gpc1515 (
      {stage0_31[211]},
      {stage1_31[88]}
   );
   gpc1_1 gpc1516 (
      {stage0_31[212]},
      {stage1_31[89]}
   );
   gpc1_1 gpc1517 (
      {stage0_31[213]},
      {stage1_31[90]}
   );
   gpc1_1 gpc1518 (
      {stage0_31[214]},
      {stage1_31[91]}
   );
   gpc1_1 gpc1519 (
      {stage0_31[215]},
      {stage1_31[92]}
   );
   gpc1_1 gpc1520 (
      {stage0_31[216]},
      {stage1_31[93]}
   );
   gpc1_1 gpc1521 (
      {stage0_31[217]},
      {stage1_31[94]}
   );
   gpc1_1 gpc1522 (
      {stage0_31[218]},
      {stage1_31[95]}
   );
   gpc1_1 gpc1523 (
      {stage0_31[219]},
      {stage1_31[96]}
   );
   gpc1_1 gpc1524 (
      {stage0_31[220]},
      {stage1_31[97]}
   );
   gpc1_1 gpc1525 (
      {stage0_31[221]},
      {stage1_31[98]}
   );
   gpc1_1 gpc1526 (
      {stage0_31[222]},
      {stage1_31[99]}
   );
   gpc1_1 gpc1527 (
      {stage0_31[223]},
      {stage1_31[100]}
   );
   gpc1_1 gpc1528 (
      {stage0_31[224]},
      {stage1_31[101]}
   );
   gpc1_1 gpc1529 (
      {stage0_31[225]},
      {stage1_31[102]}
   );
   gpc1_1 gpc1530 (
      {stage0_31[226]},
      {stage1_31[103]}
   );
   gpc1_1 gpc1531 (
      {stage0_31[227]},
      {stage1_31[104]}
   );
   gpc1_1 gpc1532 (
      {stage0_31[228]},
      {stage1_31[105]}
   );
   gpc1_1 gpc1533 (
      {stage0_31[229]},
      {stage1_31[106]}
   );
   gpc1_1 gpc1534 (
      {stage0_31[230]},
      {stage1_31[107]}
   );
   gpc1_1 gpc1535 (
      {stage0_31[231]},
      {stage1_31[108]}
   );
   gpc1_1 gpc1536 (
      {stage0_31[232]},
      {stage1_31[109]}
   );
   gpc1_1 gpc1537 (
      {stage0_31[233]},
      {stage1_31[110]}
   );
   gpc1_1 gpc1538 (
      {stage0_31[234]},
      {stage1_31[111]}
   );
   gpc1_1 gpc1539 (
      {stage0_31[235]},
      {stage1_31[112]}
   );
   gpc1_1 gpc1540 (
      {stage0_31[236]},
      {stage1_31[113]}
   );
   gpc1_1 gpc1541 (
      {stage0_31[237]},
      {stage1_31[114]}
   );
   gpc1_1 gpc1542 (
      {stage0_31[238]},
      {stage1_31[115]}
   );
   gpc1_1 gpc1543 (
      {stage0_31[239]},
      {stage1_31[116]}
   );
   gpc1_1 gpc1544 (
      {stage0_31[240]},
      {stage1_31[117]}
   );
   gpc1_1 gpc1545 (
      {stage0_31[241]},
      {stage1_31[118]}
   );
   gpc1_1 gpc1546 (
      {stage0_31[242]},
      {stage1_31[119]}
   );
   gpc1_1 gpc1547 (
      {stage0_31[243]},
      {stage1_31[120]}
   );
   gpc1_1 gpc1548 (
      {stage0_31[244]},
      {stage1_31[121]}
   );
   gpc1_1 gpc1549 (
      {stage0_31[245]},
      {stage1_31[122]}
   );
   gpc1_1 gpc1550 (
      {stage0_31[246]},
      {stage1_31[123]}
   );
   gpc1_1 gpc1551 (
      {stage0_31[247]},
      {stage1_31[124]}
   );
   gpc1_1 gpc1552 (
      {stage0_31[248]},
      {stage1_31[125]}
   );
   gpc1_1 gpc1553 (
      {stage0_31[249]},
      {stage1_31[126]}
   );
   gpc1_1 gpc1554 (
      {stage0_31[250]},
      {stage1_31[127]}
   );
   gpc1_1 gpc1555 (
      {stage0_31[251]},
      {stage1_31[128]}
   );
   gpc1_1 gpc1556 (
      {stage0_31[252]},
      {stage1_31[129]}
   );
   gpc1_1 gpc1557 (
      {stage0_31[253]},
      {stage1_31[130]}
   );
   gpc1_1 gpc1558 (
      {stage0_31[254]},
      {stage1_31[131]}
   );
   gpc1_1 gpc1559 (
      {stage0_31[255]},
      {stage1_31[132]}
   );
   gpc1163_5 gpc1560 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1561 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1562 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1563 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1564 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1565 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1566 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1567 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1568 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1569 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc1570 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc1571 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc1163_5 gpc1572 (
      {stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_2[12]},
      {stage1_3[12]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1573 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc1574 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[13]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc1575 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28]},
      {stage1_3[14]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc1576 (
      {stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage1_3[15]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[16],stage2_3[16],stage2_2[16]}
   );
   gpc615_5 gpc1577 (
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38]},
      {stage1_3[16]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[17],stage2_3[17],stage2_2[17]}
   );
   gpc615_5 gpc1578 (
      {stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43]},
      {stage1_3[17]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[18],stage2_3[18],stage2_2[18]}
   );
   gpc615_5 gpc1579 (
      {stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage1_3[18]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[19],stage2_3[19],stage2_2[19]}
   );
   gpc615_5 gpc1580 (
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_3[19]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[20],stage2_3[20],stage2_2[20]}
   );
   gpc615_5 gpc1581 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58]},
      {stage1_3[20]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[21],stage2_3[21],stage2_2[21]}
   );
   gpc615_5 gpc1582 (
      {stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage1_3[21]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[22],stage2_3[22],stage2_2[22]}
   );
   gpc615_5 gpc1583 (
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68]},
      {stage1_3[22]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc615_5 gpc1584 (
      {stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73]},
      {stage1_3[23]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[11],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc1585 (
      {stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77], stage1_2[78]},
      {stage1_3[24]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[12],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc615_5 gpc1586 (
      {stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage1_3[25]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[13],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc1587 (
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[14],stage2_5[14],stage2_4[27],stage2_3[27]}
   );
   gpc615_5 gpc1588 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[84]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[15],stage2_5[15],stage2_4[28],stage2_3[28]}
   );
   gpc615_5 gpc1589 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[85]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[16],stage2_5[16],stage2_4[29],stage2_3[29]}
   );
   gpc615_5 gpc1590 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[86]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[17],stage2_5[17],stage2_4[30],stage2_3[30]}
   );
   gpc615_5 gpc1591 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[87]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[18],stage2_5[18],stage2_4[31],stage2_3[31]}
   );
   gpc615_5 gpc1592 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[88]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[19],stage2_5[19],stage2_4[32],stage2_3[32]}
   );
   gpc615_5 gpc1593 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[89]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[20],stage2_5[20],stage2_4[33],stage2_3[33]}
   );
   gpc615_5 gpc1594 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[90]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[21],stage2_5[21],stage2_4[34],stage2_3[34]}
   );
   gpc615_5 gpc1595 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[91]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[22],stage2_5[22],stage2_4[35],stage2_3[35]}
   );
   gpc615_5 gpc1596 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[92]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[23],stage2_5[23],stage2_4[36],stage2_3[36]}
   );
   gpc615_5 gpc1597 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[93]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[24],stage2_5[24],stage2_4[37],stage2_3[37]}
   );
   gpc615_5 gpc1598 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[94]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[25],stage2_5[25],stage2_4[38],stage2_3[38]}
   );
   gpc207_4 gpc1599 (
      {stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[12],stage2_6[26],stage2_5[26],stage2_4[39]}
   );
   gpc606_5 gpc1600 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[13],stage2_6[27],stage2_5[27],stage2_4[40]}
   );
   gpc615_5 gpc1601 (
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112]},
      {stage1_5[72]},
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage2_8[1],stage2_7[14],stage2_6[28],stage2_5[28],stage2_4[41]}
   );
   gpc615_5 gpc1602 (
      {stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117]},
      {stage1_5[73]},
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19]},
      {stage2_8[2],stage2_7[15],stage2_6[29],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc1603 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[3],stage2_7[16],stage2_6[30],stage2_5[30]}
   );
   gpc606_5 gpc1604 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[4],stage2_7[17],stage2_6[31],stage2_5[31]}
   );
   gpc606_5 gpc1605 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[5],stage2_7[18],stage2_6[32],stage2_5[32]}
   );
   gpc606_5 gpc1606 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[6],stage2_7[19],stage2_6[33],stage2_5[33]}
   );
   gpc606_5 gpc1607 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[7],stage2_7[20],stage2_6[34],stage2_5[34]}
   );
   gpc606_5 gpc1608 (
      {stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108], stage1_5[109]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[8],stage2_7[21],stage2_6[35],stage2_5[35]}
   );
   gpc606_5 gpc1609 (
      {stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113], stage1_5[114], stage1_5[115]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[9],stage2_7[22],stage2_6[36],stage2_5[36]}
   );
   gpc606_5 gpc1610 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[10],stage2_7[23],stage2_6[37],stage2_5[37]}
   );
   gpc606_5 gpc1611 (
      {stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[8],stage2_8[11],stage2_7[24],stage2_6[38]}
   );
   gpc615_5 gpc1612 (
      {stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage1_7[48]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[9],stage2_8[12],stage2_7[25],stage2_6[39]}
   );
   gpc615_5 gpc1613 (
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_7[49]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[10],stage2_8[13],stage2_7[26],stage2_6[40]}
   );
   gpc615_5 gpc1614 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40]},
      {stage1_7[50]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[11],stage2_8[14],stage2_7[27],stage2_6[41]}
   );
   gpc615_5 gpc1615 (
      {stage1_6[41], stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45]},
      {stage1_7[51]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[12],stage2_8[15],stage2_7[28],stage2_6[42]}
   );
   gpc615_5 gpc1616 (
      {stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50]},
      {stage1_7[52]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[13],stage2_8[16],stage2_7[29],stage2_6[43]}
   );
   gpc615_5 gpc1617 (
      {stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage1_7[53]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[14],stage2_8[17],stage2_7[30],stage2_6[44]}
   );
   gpc615_5 gpc1618 (
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage1_7[54]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[15],stage2_8[18],stage2_7[31],stage2_6[45]}
   );
   gpc615_5 gpc1619 (
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_7[55]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[16],stage2_8[19],stage2_7[32],stage2_6[46]}
   );
   gpc615_5 gpc1620 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70]},
      {stage1_7[56]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[17],stage2_8[20],stage2_7[33],stage2_6[47]}
   );
   gpc615_5 gpc1621 (
      {stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75]},
      {stage1_7[57]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[18],stage2_8[21],stage2_7[34],stage2_6[48]}
   );
   gpc615_5 gpc1622 (
      {stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80]},
      {stage1_7[58]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[19],stage2_8[22],stage2_7[35],stage2_6[49]}
   );
   gpc615_5 gpc1623 (
      {stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage1_7[59]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[20],stage2_8[23],stage2_7[36],stage2_6[50]}
   );
   gpc615_5 gpc1624 (
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_7[60]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[21],stage2_8[24],stage2_7[37],stage2_6[51]}
   );
   gpc615_5 gpc1625 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_7[61]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[22],stage2_8[25],stage2_7[38],stage2_6[52]}
   );
   gpc615_5 gpc1626 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[90]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[15],stage2_9[23],stage2_8[26],stage2_7[39]}
   );
   gpc615_5 gpc1627 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[91]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[16],stage2_9[24],stage2_8[27],stage2_7[40]}
   );
   gpc615_5 gpc1628 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[92]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[17],stage2_9[25],stage2_8[28],stage2_7[41]}
   );
   gpc615_5 gpc1629 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[93]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[18],stage2_9[26],stage2_8[29],stage2_7[42]}
   );
   gpc615_5 gpc1630 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[94]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[19],stage2_9[27],stage2_8[30],stage2_7[43]}
   );
   gpc615_5 gpc1631 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[95]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[20],stage2_9[28],stage2_8[31],stage2_7[44]}
   );
   gpc606_5 gpc1632 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[6],stage2_10[21],stage2_9[29]}
   );
   gpc606_5 gpc1633 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[1],stage2_11[7],stage2_10[22],stage2_9[30]}
   );
   gpc606_5 gpc1634 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[2],stage2_11[8],stage2_10[23],stage2_9[31]}
   );
   gpc606_5 gpc1635 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[3],stage2_11[9],stage2_10[24],stage2_9[32]}
   );
   gpc606_5 gpc1636 (
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[4],stage2_11[10],stage2_10[25],stage2_9[33]}
   );
   gpc606_5 gpc1637 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[5],stage2_11[11],stage2_10[26],stage2_9[34]}
   );
   gpc606_5 gpc1638 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[6],stage2_11[12],stage2_10[27],stage2_9[35]}
   );
   gpc606_5 gpc1639 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[7],stage2_11[13],stage2_10[28],stage2_9[36]}
   );
   gpc606_5 gpc1640 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[8],stage2_11[14],stage2_10[29],stage2_9[37]}
   );
   gpc606_5 gpc1641 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[9],stage2_11[15],stage2_10[30],stage2_9[38]}
   );
   gpc606_5 gpc1642 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[10],stage2_11[16],stage2_10[31],stage2_9[39]}
   );
   gpc615_5 gpc1643 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106]},
      {stage1_10[0]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[11],stage2_11[17],stage2_10[32],stage2_9[40]}
   );
   gpc606_5 gpc1644 (
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[12],stage2_12[12],stage2_11[18],stage2_10[33]}
   );
   gpc606_5 gpc1645 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[13],stage2_12[13],stage2_11[19],stage2_10[34]}
   );
   gpc606_5 gpc1646 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[14],stage2_12[14],stage2_11[20],stage2_10[35]}
   );
   gpc606_5 gpc1647 (
      {stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[15],stage2_12[15],stage2_11[21],stage2_10[36]}
   );
   gpc606_5 gpc1648 (
      {stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[16],stage2_12[16],stage2_11[22],stage2_10[37]}
   );
   gpc606_5 gpc1649 (
      {stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[17],stage2_12[17],stage2_11[23],stage2_10[38]}
   );
   gpc606_5 gpc1650 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[18],stage2_12[18],stage2_11[24],stage2_10[39]}
   );
   gpc606_5 gpc1651 (
      {stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[19],stage2_12[19],stage2_11[25],stage2_10[40]}
   );
   gpc606_5 gpc1652 (
      {stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[20],stage2_12[20],stage2_11[26],stage2_10[41]}
   );
   gpc606_5 gpc1653 (
      {stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[21],stage2_12[21],stage2_11[27],stage2_10[42]}
   );
   gpc606_5 gpc1654 (
      {stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65], stage1_10[66]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[22],stage2_12[22],stage2_11[28],stage2_10[43]}
   );
   gpc606_5 gpc1655 (
      {stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[23],stage2_12[23],stage2_11[29],stage2_10[44]}
   );
   gpc606_5 gpc1656 (
      {stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[24],stage2_12[24],stage2_11[30],stage2_10[45]}
   );
   gpc606_5 gpc1657 (
      {stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[25],stage2_12[25],stage2_11[31],stage2_10[46]}
   );
   gpc606_5 gpc1658 (
      {stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[26],stage2_12[26],stage2_11[32],stage2_10[47]}
   );
   gpc606_5 gpc1659 (
      {stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[27],stage2_12[27],stage2_11[33],stage2_10[48]}
   );
   gpc615_5 gpc1660 (
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76]},
      {stage1_12[96]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[16],stage2_13[28],stage2_12[28],stage2_11[34]}
   );
   gpc615_5 gpc1661 (
      {stage1_11[77], stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81]},
      {stage1_12[97]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[17],stage2_13[29],stage2_12[29],stage2_11[35]}
   );
   gpc615_5 gpc1662 (
      {stage1_11[82], stage1_11[83], stage1_11[84], stage1_11[85], stage1_11[86]},
      {stage1_12[98]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[18],stage2_13[30],stage2_12[30],stage2_11[36]}
   );
   gpc615_5 gpc1663 (
      {stage1_11[87], stage1_11[88], stage1_11[89], stage1_11[90], stage1_11[91]},
      {stage1_12[99]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[19],stage2_13[31],stage2_12[31],stage2_11[37]}
   );
   gpc615_5 gpc1664 (
      {stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95], stage1_11[96]},
      {stage1_12[100]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[20],stage2_13[32],stage2_12[32],stage2_11[38]}
   );
   gpc615_5 gpc1665 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage1_12[101]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[21],stage2_13[33],stage2_12[33],stage2_11[39]}
   );
   gpc615_5 gpc1666 (
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106]},
      {stage1_12[102]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[22],stage2_13[34],stage2_12[34],stage2_11[40]}
   );
   gpc615_5 gpc1667 (
      {stage1_11[107], stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111]},
      {stage1_12[103]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[23],stage2_13[35],stage2_12[35],stage2_11[41]}
   );
   gpc615_5 gpc1668 (
      {stage1_11[112], stage1_11[113], stage1_11[114], stage1_11[115], stage1_11[116]},
      {stage1_12[104]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[24],stage2_13[36],stage2_12[36],stage2_11[42]}
   );
   gpc615_5 gpc1669 (
      {stage1_11[117], stage1_11[118], stage1_11[119], stage1_11[120], stage1_11[121]},
      {stage1_12[105]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[25],stage2_13[37],stage2_12[37],stage2_11[43]}
   );
   gpc615_5 gpc1670 (
      {stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125], stage1_11[126]},
      {stage1_12[106]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[26],stage2_13[38],stage2_12[38],stage2_11[44]}
   );
   gpc606_5 gpc1671 (
      {stage1_12[107], stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[11],stage2_14[27],stage2_13[39],stage2_12[39]}
   );
   gpc606_5 gpc1672 (
      {stage1_12[113], stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[12],stage2_14[28],stage2_13[40],stage2_12[40]}
   );
   gpc606_5 gpc1673 (
      {stage1_12[119], stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[13],stage2_14[29],stage2_13[41],stage2_12[41]}
   );
   gpc606_5 gpc1674 (
      {stage1_12[125], stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[14],stage2_14[30],stage2_13[42],stage2_12[42]}
   );
   gpc606_5 gpc1675 (
      {stage1_12[131], stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[15],stage2_14[31],stage2_13[43],stage2_12[43]}
   );
   gpc606_5 gpc1676 (
      {stage1_12[137], stage1_12[138], stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[16],stage2_14[32],stage2_13[44],stage2_12[44]}
   );
   gpc606_5 gpc1677 (
      {stage1_12[143], stage1_12[144], stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[17],stage2_14[33],stage2_13[45],stage2_12[45]}
   );
   gpc606_5 gpc1678 (
      {stage1_12[149], stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[18],stage2_14[34],stage2_13[46],stage2_12[46]}
   );
   gpc606_5 gpc1679 (
      {stage1_12[155], stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[19],stage2_14[35],stage2_13[47],stage2_12[47]}
   );
   gpc606_5 gpc1680 (
      {stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[20],stage2_14[36],stage2_13[48],stage2_12[48]}
   );
   gpc606_5 gpc1681 (
      {stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[21],stage2_14[37],stage2_13[49],stage2_12[49]}
   );
   gpc606_5 gpc1682 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[11],stage2_15[22],stage2_14[38],stage2_13[50]}
   );
   gpc606_5 gpc1683 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[12],stage2_15[23],stage2_14[39],stage2_13[51]}
   );
   gpc606_5 gpc1684 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[13],stage2_15[24],stage2_14[40],stage2_13[52]}
   );
   gpc606_5 gpc1685 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[14],stage2_15[25],stage2_14[41],stage2_13[53]}
   );
   gpc615_5 gpc1686 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[15],stage2_15[26]}
   );
   gpc615_5 gpc1687 (
      {stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[16],stage2_15[27]}
   );
   gpc615_5 gpc1688 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38]},
      {stage1_16[2]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[17],stage2_15[28]}
   );
   gpc615_5 gpc1689 (
      {stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_16[3]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[3],stage2_17[7],stage2_16[18],stage2_15[29]}
   );
   gpc615_5 gpc1690 (
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48]},
      {stage1_16[4]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[4],stage2_17[8],stage2_16[19],stage2_15[30]}
   );
   gpc615_5 gpc1691 (
      {stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage1_16[5]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[5],stage2_17[9],stage2_16[20],stage2_15[31]}
   );
   gpc615_5 gpc1692 (
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58]},
      {stage1_16[6]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[6],stage2_17[10],stage2_16[21],stage2_15[32]}
   );
   gpc615_5 gpc1693 (
      {stage1_15[59], stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63]},
      {stage1_16[7]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[7],stage2_17[11],stage2_16[22],stage2_15[33]}
   );
   gpc615_5 gpc1694 (
      {stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67], stage1_15[68]},
      {stage1_16[8]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[8],stage2_17[12],stage2_16[23],stage2_15[34]}
   );
   gpc615_5 gpc1695 (
      {stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage1_16[9]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[9],stage2_17[13],stage2_16[24],stage2_15[35]}
   );
   gpc615_5 gpc1696 (
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78]},
      {stage1_16[10]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[10],stage2_17[14],stage2_16[25],stage2_15[36]}
   );
   gpc615_5 gpc1697 (
      {stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage1_16[11]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[11],stage2_17[15],stage2_16[26],stage2_15[37]}
   );
   gpc606_5 gpc1698 (
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[12],stage2_18[12],stage2_17[16],stage2_16[27]}
   );
   gpc606_5 gpc1699 (
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[13],stage2_18[13],stage2_17[17],stage2_16[28]}
   );
   gpc606_5 gpc1700 (
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[14],stage2_18[14],stage2_17[18],stage2_16[29]}
   );
   gpc606_5 gpc1701 (
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[15],stage2_18[15],stage2_17[19],stage2_16[30]}
   );
   gpc606_5 gpc1702 (
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[16],stage2_18[16],stage2_17[20],stage2_16[31]}
   );
   gpc606_5 gpc1703 (
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[17],stage2_18[17],stage2_17[21],stage2_16[32]}
   );
   gpc606_5 gpc1704 (
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[18],stage2_18[18],stage2_17[22],stage2_16[33]}
   );
   gpc606_5 gpc1705 (
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[19],stage2_18[19],stage2_17[23],stage2_16[34]}
   );
   gpc606_5 gpc1706 (
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[20],stage2_18[20],stage2_17[24],stage2_16[35]}
   );
   gpc606_5 gpc1707 (
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[21],stage2_18[21],stage2_17[25],stage2_16[36]}
   );
   gpc606_5 gpc1708 (
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[22],stage2_18[22],stage2_17[26],stage2_16[37]}
   );
   gpc606_5 gpc1709 (
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[23],stage2_18[23],stage2_17[27],stage2_16[38]}
   );
   gpc606_5 gpc1710 (
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[24],stage2_18[24],stage2_17[28],stage2_16[39]}
   );
   gpc606_5 gpc1711 (
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[25],stage2_18[25],stage2_17[29],stage2_16[40]}
   );
   gpc606_5 gpc1712 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[14],stage2_19[26],stage2_18[26],stage2_17[30]}
   );
   gpc606_5 gpc1713 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[15],stage2_19[27],stage2_18[27],stage2_17[31]}
   );
   gpc606_5 gpc1714 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[16],stage2_19[28],stage2_18[28],stage2_17[32]}
   );
   gpc606_5 gpc1715 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[17],stage2_19[29],stage2_18[29],stage2_17[33]}
   );
   gpc606_5 gpc1716 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[18],stage2_19[30],stage2_18[30],stage2_17[34]}
   );
   gpc606_5 gpc1717 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[19],stage2_19[31],stage2_18[31],stage2_17[35]}
   );
   gpc615_5 gpc1718 (
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88]},
      {stage1_19[36]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[6],stage2_20[20],stage2_19[32],stage2_18[32]}
   );
   gpc615_5 gpc1719 (
      {stage1_18[89], stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93]},
      {stage1_19[37]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[7],stage2_20[21],stage2_19[33],stage2_18[33]}
   );
   gpc615_5 gpc1720 (
      {stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42]},
      {stage1_20[12]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[2],stage2_21[8],stage2_20[22],stage2_19[34]}
   );
   gpc615_5 gpc1721 (
      {stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_20[13]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[3],stage2_21[9],stage2_20[23],stage2_19[35]}
   );
   gpc615_5 gpc1722 (
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52]},
      {stage1_20[14]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[4],stage2_21[10],stage2_20[24],stage2_19[36]}
   );
   gpc615_5 gpc1723 (
      {stage1_19[53], stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57]},
      {stage1_20[15]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[5],stage2_21[11],stage2_20[25],stage2_19[37]}
   );
   gpc615_5 gpc1724 (
      {stage1_19[58], stage1_19[59], stage1_19[60], stage1_19[61], stage1_19[62]},
      {stage1_20[16]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[6],stage2_21[12],stage2_20[26],stage2_19[38]}
   );
   gpc615_5 gpc1725 (
      {stage1_19[63], stage1_19[64], stage1_19[65], stage1_19[66], stage1_19[67]},
      {stage1_20[17]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[7],stage2_21[13],stage2_20[27],stage2_19[39]}
   );
   gpc615_5 gpc1726 (
      {stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71], stage1_19[72]},
      {stage1_20[18]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[8],stage2_21[14],stage2_20[28],stage2_19[40]}
   );
   gpc615_5 gpc1727 (
      {stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage1_20[19]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[9],stage2_21[15],stage2_20[29],stage2_19[41]}
   );
   gpc615_5 gpc1728 (
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82]},
      {stage1_20[20]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[10],stage2_21[16],stage2_20[30],stage2_19[42]}
   );
   gpc615_5 gpc1729 (
      {stage1_19[83], stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87]},
      {stage1_20[21]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[11],stage2_21[17],stage2_20[31],stage2_19[43]}
   );
   gpc615_5 gpc1730 (
      {stage1_19[88], stage1_19[89], stage1_19[90], stage1_19[91], stage1_19[92]},
      {stage1_20[22]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[12],stage2_21[18],stage2_20[32],stage2_19[44]}
   );
   gpc606_5 gpc1731 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[11],stage2_22[13],stage2_21[19]}
   );
   gpc606_5 gpc1732 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[1],stage2_23[12],stage2_22[14],stage2_21[20]}
   );
   gpc606_5 gpc1733 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[2],stage2_23[13],stage2_22[15],stage2_21[21]}
   );
   gpc606_5 gpc1734 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[3],stage2_23[14],stage2_22[16],stage2_21[22]}
   );
   gpc606_5 gpc1735 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[4],stage2_23[15],stage2_22[17]}
   );
   gpc606_5 gpc1736 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[5],stage2_23[16],stage2_22[18]}
   );
   gpc606_5 gpc1737 (
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[6],stage2_23[17],stage2_22[19]}
   );
   gpc606_5 gpc1738 (
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[7],stage2_23[18],stage2_22[20]}
   );
   gpc606_5 gpc1739 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[8],stage2_23[19],stage2_22[21]}
   );
   gpc606_5 gpc1740 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[9],stage2_24[9],stage2_23[20],stage2_22[22]}
   );
   gpc606_5 gpc1741 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[10],stage2_24[10],stage2_23[21],stage2_22[23]}
   );
   gpc606_5 gpc1742 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[11],stage2_24[11],stage2_23[22],stage2_22[24]}
   );
   gpc606_5 gpc1743 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[12],stage2_24[12],stage2_23[23],stage2_22[25]}
   );
   gpc606_5 gpc1744 (
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[13],stage2_24[13],stage2_23[24],stage2_22[26]}
   );
   gpc606_5 gpc1745 (
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[14],stage2_24[14],stage2_23[25],stage2_22[27]}
   );
   gpc606_5 gpc1746 (
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[15],stage2_24[15],stage2_23[26],stage2_22[28]}
   );
   gpc615_5 gpc1747 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76]},
      {stage1_23[24]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[16],stage2_24[16],stage2_23[27],stage2_22[29]}
   );
   gpc606_5 gpc1748 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29], stage1_23[30]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[13],stage2_25[17],stage2_24[17],stage2_23[28]}
   );
   gpc606_5 gpc1749 (
      {stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[14],stage2_25[18],stage2_24[18],stage2_23[29]}
   );
   gpc606_5 gpc1750 (
      {stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[15],stage2_25[19],stage2_24[19],stage2_23[30]}
   );
   gpc606_5 gpc1751 (
      {stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47], stage1_23[48]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[16],stage2_25[20],stage2_24[20],stage2_23[31]}
   );
   gpc606_5 gpc1752 (
      {stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53], stage1_23[54]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[17],stage2_25[21],stage2_24[21],stage2_23[32]}
   );
   gpc606_5 gpc1753 (
      {stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59], stage1_23[60]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[18],stage2_25[22],stage2_24[22],stage2_23[33]}
   );
   gpc606_5 gpc1754 (
      {stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[19],stage2_25[23],stage2_24[23],stage2_23[34]}
   );
   gpc606_5 gpc1755 (
      {stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[20],stage2_25[24],stage2_24[24],stage2_23[35]}
   );
   gpc606_5 gpc1756 (
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[21],stage2_25[25],stage2_24[25]}
   );
   gpc615_5 gpc1757 (
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88]},
      {stage1_25[48]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[22],stage2_25[26],stage2_24[26]}
   );
   gpc615_5 gpc1758 (
      {stage1_24[89], stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93]},
      {stage1_25[49]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[23],stage2_25[27],stage2_24[27]}
   );
   gpc615_5 gpc1759 (
      {stage1_24[94], stage1_24[95], stage1_24[96], stage1_24[97], stage1_24[98]},
      {stage1_25[50]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[24],stage2_25[28],stage2_24[28]}
   );
   gpc615_5 gpc1760 (
      {stage1_24[99], stage1_24[100], stage1_24[101], stage1_24[102], stage1_24[103]},
      {stage1_25[51]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[12],stage2_26[25],stage2_25[29],stage2_24[29]}
   );
   gpc615_5 gpc1761 (
      {stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107], stage1_24[108]},
      {stage1_25[52]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[13],stage2_26[26],stage2_25[30],stage2_24[30]}
   );
   gpc615_5 gpc1762 (
      {stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage1_25[53]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[14],stage2_26[27],stage2_25[31],stage2_24[31]}
   );
   gpc615_5 gpc1763 (
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118]},
      {stage1_25[54]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[15],stage2_26[28],stage2_25[32],stage2_24[32]}
   );
   gpc615_5 gpc1764 (
      {stage1_24[119], stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123]},
      {stage1_25[55]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[16],stage2_26[29],stage2_25[33],stage2_24[33]}
   );
   gpc615_5 gpc1765 (
      {stage1_24[124], stage1_24[125], stage1_24[126], stage1_24[127], stage1_24[128]},
      {stage1_25[56]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[17],stage2_26[30],stage2_25[34],stage2_24[34]}
   );
   gpc615_5 gpc1766 (
      {stage1_24[129], stage1_24[130], stage1_24[131], stage1_24[132], stage1_24[133]},
      {stage1_25[57]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[18],stage2_26[31],stage2_25[35],stage2_24[35]}
   );
   gpc615_5 gpc1767 (
      {stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137], stage1_24[138]},
      {stage1_25[58]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[19],stage2_26[32],stage2_25[36],stage2_24[36]}
   );
   gpc615_5 gpc1768 (
      {stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143]},
      {stage1_25[59]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[20],stage2_26[33],stage2_25[37],stage2_24[37]}
   );
   gpc615_5 gpc1769 (
      {stage1_24[144], stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148]},
      {stage1_25[60]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[21],stage2_26[34],stage2_25[38],stage2_24[38]}
   );
   gpc615_5 gpc1770 (
      {stage1_24[149], stage1_24[150], stage1_24[151], stage1_24[152], stage1_24[153]},
      {stage1_25[61]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[22],stage2_26[35],stage2_25[39],stage2_24[39]}
   );
   gpc615_5 gpc1771 (
      {stage1_24[154], stage1_24[155], stage1_24[156], stage1_24[157], stage1_24[158]},
      {stage1_25[62]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[23],stage2_26[36],stage2_25[40],stage2_24[40]}
   );
   gpc615_5 gpc1772 (
      {stage1_24[159], stage1_24[160], stage1_24[161], stage1_24[162], stage1_24[163]},
      {stage1_25[63]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[24],stage2_26[37],stage2_25[41],stage2_24[41]}
   );
   gpc615_5 gpc1773 (
      {stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167], stage1_24[168]},
      {stage1_25[64]},
      {stage1_26[102], stage1_26[103], stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107]},
      {stage2_28[17],stage2_27[25],stage2_26[38],stage2_25[42],stage2_24[42]}
   );
   gpc615_5 gpc1774 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_25[65]},
      {stage1_26[108], stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage2_28[18],stage2_27[26],stage2_26[39],stage2_25[43],stage2_24[43]}
   );
   gpc615_5 gpc1775 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178]},
      {stage1_25[66]},
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage2_28[19],stage2_27[27],stage2_26[40],stage2_25[44],stage2_24[44]}
   );
   gpc615_5 gpc1776 (
      {stage1_24[179], stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183]},
      {stage1_25[67]},
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage2_28[20],stage2_27[28],stage2_26[41],stage2_25[45],stage2_24[45]}
   );
   gpc615_5 gpc1777 (
      {stage1_24[184], stage1_24[185], stage1_24[186], stage1_24[187], stage1_24[188]},
      {stage1_25[68]},
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130], stage1_26[131]},
      {stage2_28[21],stage2_27[29],stage2_26[42],stage2_25[46],stage2_24[46]}
   );
   gpc615_5 gpc1778 (
      {stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192], stage1_24[193]},
      {stage1_25[69]},
      {stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135], stage1_26[136], stage1_26[137]},
      {stage2_28[22],stage2_27[30],stage2_26[43],stage2_25[47],stage2_24[47]}
   );
   gpc615_5 gpc1779 (
      {stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197], stage1_24[198]},
      {stage1_25[70]},
      {stage1_26[138], stage1_26[139], stage1_26[140], stage1_26[141], stage1_26[142], stage1_26[143]},
      {stage2_28[23],stage2_27[31],stage2_26[44],stage2_25[48],stage2_24[48]}
   );
   gpc615_5 gpc1780 (
      {stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203]},
      {stage1_25[71]},
      {stage1_26[144], stage1_26[145], stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149]},
      {stage2_28[24],stage2_27[32],stage2_26[45],stage2_25[49],stage2_24[49]}
   );
   gpc615_5 gpc1781 (
      {stage1_24[204], stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208]},
      {stage1_25[72]},
      {stage1_26[150], stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154], stage1_26[155]},
      {stage2_28[25],stage2_27[33],stage2_26[46],stage2_25[50],stage2_24[50]}
   );
   gpc615_5 gpc1782 (
      {stage1_24[209], stage1_24[210], stage1_24[211], stage1_24[212], stage1_24[213]},
      {stage1_25[73]},
      {stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159], stage1_26[160], stage1_26[161]},
      {stage2_28[26],stage2_27[34],stage2_26[47],stage2_25[51],stage2_24[51]}
   );
   gpc615_5 gpc1783 (
      {stage1_24[214], stage1_24[215], stage1_24[216], stage1_24[217], stage1_24[218]},
      {stage1_25[74]},
      {stage1_26[162], stage1_26[163], stage1_26[164], stage1_26[165], stage1_26[166], stage1_26[167]},
      {stage2_28[27],stage2_27[35],stage2_26[48],stage2_25[52],stage2_24[52]}
   );
   gpc615_5 gpc1784 (
      {stage1_24[219], stage1_24[220], stage1_24[221], stage1_24[222], stage1_24[223]},
      {stage1_25[75]},
      {stage1_26[168], stage1_26[169], stage1_26[170], stage1_26[171], stage1_26[172], stage1_26[173]},
      {stage2_28[28],stage2_27[36],stage2_26[49],stage2_25[53],stage2_24[53]}
   );
   gpc615_5 gpc1785 (
      {stage1_24[224], stage1_24[225], stage1_24[226], stage1_24[227], stage1_24[228]},
      {stage1_25[76]},
      {stage1_26[174], stage1_26[175], stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179]},
      {stage2_28[29],stage2_27[37],stage2_26[50],stage2_25[54],stage2_24[54]}
   );
   gpc615_5 gpc1786 (
      {stage1_24[229], stage1_24[230], stage1_24[231], stage1_24[232], stage1_24[233]},
      {stage1_25[77]},
      {stage1_26[180], stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184], stage1_26[185]},
      {stage2_28[30],stage2_27[38],stage2_26[51],stage2_25[55],stage2_24[55]}
   );
   gpc615_5 gpc1787 (
      {stage1_24[234], stage1_24[235], stage1_24[236], stage1_24[237], stage1_24[238]},
      {stage1_25[78]},
      {stage1_26[186], stage1_26[187], stage1_26[188], stage1_26[189], stage1_26[190], stage1_26[191]},
      {stage2_28[31],stage2_27[39],stage2_26[52],stage2_25[56],stage2_24[56]}
   );
   gpc615_5 gpc1788 (
      {stage1_24[239], stage1_24[240], stage1_24[241], stage1_24[242], stage1_24[243]},
      {stage1_25[79]},
      {stage1_26[192], stage1_26[193], stage1_26[194], stage1_26[195], stage1_26[196], stage1_26[197]},
      {stage2_28[32],stage2_27[40],stage2_26[53],stage2_25[57],stage2_24[57]}
   );
   gpc615_5 gpc1789 (
      {stage1_24[244], stage1_24[245], stage1_24[246], stage1_24[247], stage1_24[248]},
      {stage1_25[80]},
      {stage1_26[198], stage1_26[199], stage1_26[200], stage1_26[201], stage1_26[202], stage1_26[203]},
      {stage2_28[33],stage2_27[41],stage2_26[54],stage2_25[58],stage2_24[58]}
   );
   gpc606_5 gpc1790 (
      {stage1_25[81], stage1_25[82], stage1_25[83], stage1_25[84], stage1_25[85], stage1_25[86]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[34],stage2_27[42],stage2_26[55],stage2_25[59]}
   );
   gpc606_5 gpc1791 (
      {stage1_25[87], stage1_25[88], stage1_25[89], stage1_25[90], stage1_25[91], stage1_25[92]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[35],stage2_27[43],stage2_26[56],stage2_25[60]}
   );
   gpc606_5 gpc1792 (
      {stage1_25[93], stage1_25[94], stage1_25[95], stage1_25[96], stage1_25[97], stage1_25[98]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[36],stage2_27[44],stage2_26[57],stage2_25[61]}
   );
   gpc606_5 gpc1793 (
      {stage1_25[99], stage1_25[100], stage1_25[101], stage1_25[102], stage1_25[103], stage1_25[104]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[37],stage2_27[45],stage2_26[58],stage2_25[62]}
   );
   gpc606_5 gpc1794 (
      {stage1_25[105], stage1_25[106], stage1_25[107], stage1_25[108], stage1_25[109], stage1_25[110]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[38],stage2_27[46],stage2_26[59],stage2_25[63]}
   );
   gpc606_5 gpc1795 (
      {stage1_25[111], stage1_25[112], stage1_25[113], stage1_25[114], stage1_25[115], stage1_25[116]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[39],stage2_27[47],stage2_26[60],stage2_25[64]}
   );
   gpc615_5 gpc1796 (
      {stage1_26[204], stage1_26[205], stage1_26[206], stage1_26[207], stage1_26[208]},
      {stage1_27[36]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[6],stage2_28[40],stage2_27[48],stage2_26[61]}
   );
   gpc615_5 gpc1797 (
      {stage1_26[209], stage1_26[210], stage1_26[211], stage1_26[212], stage1_26[213]},
      {stage1_27[37]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[7],stage2_28[41],stage2_27[49],stage2_26[62]}
   );
   gpc615_5 gpc1798 (
      {stage1_26[214], stage1_26[215], stage1_26[216], stage1_26[217], stage1_26[218]},
      {stage1_27[38]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[8],stage2_28[42],stage2_27[50],stage2_26[63]}
   );
   gpc615_5 gpc1799 (
      {stage1_26[219], stage1_26[220], stage1_26[221], stage1_26[222], stage1_26[223]},
      {stage1_27[39]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[9],stage2_28[43],stage2_27[51],stage2_26[64]}
   );
   gpc615_5 gpc1800 (
      {stage1_26[224], stage1_26[225], stage1_26[226], stage1_26[227], stage1_26[228]},
      {stage1_27[40]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[10],stage2_28[44],stage2_27[52],stage2_26[65]}
   );
   gpc615_5 gpc1801 (
      {stage1_26[229], stage1_26[230], stage1_26[231], stage1_26[232], stage1_26[233]},
      {stage1_27[41]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[11],stage2_28[45],stage2_27[53],stage2_26[66]}
   );
   gpc615_5 gpc1802 (
      {stage1_26[234], stage1_26[235], stage1_26[236], 1'b0, 1'b0},
      {stage1_27[42]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[12],stage2_28[46],stage2_27[54],stage2_26[67]}
   );
   gpc615_5 gpc1803 (
      {stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage1_28[42]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[13],stage2_28[47],stage2_27[55]}
   );
   gpc615_5 gpc1804 (
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_28[43]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[14],stage2_28[48],stage2_27[56]}
   );
   gpc615_5 gpc1805 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[44]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[9],stage2_29[15],stage2_28[49],stage2_27[57]}
   );
   gpc615_5 gpc1806 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[45]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[10],stage2_29[16],stage2_28[50],stage2_27[58]}
   );
   gpc615_5 gpc1807 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[46]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[11],stage2_29[17],stage2_28[51],stage2_27[59]}
   );
   gpc615_5 gpc1808 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[47]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[12],stage2_29[18],stage2_28[52],stage2_27[60]}
   );
   gpc606_5 gpc1809 (
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[6],stage2_30[13],stage2_29[19],stage2_28[53]}
   );
   gpc606_5 gpc1810 (
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[7],stage2_30[14],stage2_29[20],stage2_28[54]}
   );
   gpc606_5 gpc1811 (
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[8],stage2_30[15],stage2_29[21],stage2_28[55]}
   );
   gpc606_5 gpc1812 (
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[9],stage2_30[16],stage2_29[22],stage2_28[56]}
   );
   gpc606_5 gpc1813 (
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[10],stage2_30[17],stage2_29[23],stage2_28[57]}
   );
   gpc606_5 gpc1814 (
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[11],stage2_30[18],stage2_29[24],stage2_28[58]}
   );
   gpc606_5 gpc1815 (
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[12],stage2_30[19],stage2_29[25],stage2_28[59]}
   );
   gpc606_5 gpc1816 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[7],stage2_31[13],stage2_30[20],stage2_29[26]}
   );
   gpc606_5 gpc1817 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[8],stage2_31[14],stage2_30[21],stage2_29[27]}
   );
   gpc606_5 gpc1818 (
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[9],stage2_31[15],stage2_30[22],stage2_29[28]}
   );
   gpc606_5 gpc1819 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[10],stage2_31[16],stage2_30[23],stage2_29[29]}
   );
   gpc606_5 gpc1820 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[11],stage2_31[17],stage2_30[24],stage2_29[30]}
   );
   gpc606_5 gpc1821 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[12],stage2_31[18],stage2_30[25],stage2_29[31]}
   );
   gpc606_5 gpc1822 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[13],stage2_31[19],stage2_30[26],stage2_29[32]}
   );
   gpc606_5 gpc1823 (
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[14],stage2_31[20],stage2_30[27],stage2_29[33]}
   );
   gpc606_5 gpc1824 (
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[15],stage2_31[21],stage2_30[28],stage2_29[34]}
   );
   gpc606_5 gpc1825 (
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[16],stage2_31[22],stage2_30[29],stage2_29[35]}
   );
   gpc606_5 gpc1826 (
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[17],stage2_31[23],stage2_30[30],stage2_29[36]}
   );
   gpc606_5 gpc1827 (
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage2_33[11],stage2_32[18],stage2_31[24],stage2_30[31],stage2_29[37]}
   );
   gpc606_5 gpc1828 (
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage2_33[12],stage2_32[19],stage2_31[25],stage2_30[32],stage2_29[38]}
   );
   gpc606_5 gpc1829 (
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], 1'b0, 1'b0},
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage2_33[13],stage2_32[20],stage2_31[26],stage2_30[33],stage2_29[39]}
   );
   gpc615_5 gpc1830 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46]},
      {stage1_31[84]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[14],stage2_32[21],stage2_31[27],stage2_30[34]}
   );
   gpc615_5 gpc1831 (
      {stage1_30[47], stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51]},
      {stage1_31[85]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[15],stage2_32[22],stage2_31[28],stage2_30[35]}
   );
   gpc615_5 gpc1832 (
      {stage1_30[52], stage1_30[53], stage1_30[54], stage1_30[55], stage1_30[56]},
      {stage1_31[86]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[16],stage2_32[23],stage2_31[29],stage2_30[36]}
   );
   gpc615_5 gpc1833 (
      {stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61]},
      {stage1_31[87]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[17],stage2_32[24],stage2_31[30],stage2_30[37]}
   );
   gpc615_5 gpc1834 (
      {stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66]},
      {stage1_31[88]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[18],stage2_32[25],stage2_31[31],stage2_30[38]}
   );
   gpc615_5 gpc1835 (
      {stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_31[89]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[19],stage2_32[26],stage2_31[32],stage2_30[39]}
   );
   gpc615_5 gpc1836 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76]},
      {stage1_31[90]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[20],stage2_32[27],stage2_31[33],stage2_30[40]}
   );
   gpc615_5 gpc1837 (
      {stage1_30[77], stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81]},
      {stage1_31[91]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[21],stage2_32[28],stage2_31[34],stage2_30[41]}
   );
   gpc615_5 gpc1838 (
      {stage1_30[82], stage1_30[83], stage1_30[84], stage1_30[85], stage1_30[86]},
      {stage1_31[92]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[22],stage2_32[29],stage2_31[35],stage2_30[42]}
   );
   gpc615_5 gpc1839 (
      {stage1_30[87], stage1_30[88], stage1_30[89], stage1_30[90], stage1_30[91]},
      {stage1_31[93]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[23],stage2_32[30],stage2_31[36],stage2_30[43]}
   );
   gpc615_5 gpc1840 (
      {stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95], stage1_30[96]},
      {stage1_31[94]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[24],stage2_32[31],stage2_31[37],stage2_30[44]}
   );
   gpc606_5 gpc1841 (
      {stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[11],stage2_33[25],stage2_32[32],stage2_31[38]}
   );
   gpc606_5 gpc1842 (
      {stage1_31[101], stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[12],stage2_33[26],stage2_32[33],stage2_31[39]}
   );
   gpc606_5 gpc1843 (
      {stage1_31[107], stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[13],stage2_33[27],stage2_32[34],stage2_31[40]}
   );
   gpc606_5 gpc1844 (
      {stage1_31[113], stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[14],stage2_33[28],stage2_32[35],stage2_31[41]}
   );
   gpc615_5 gpc1845 (
      {stage1_31[119], stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123]},
      {stage1_32[66]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[15],stage2_33[29],stage2_32[36],stage2_31[42]}
   );
   gpc615_5 gpc1846 (
      {stage1_31[124], stage1_31[125], stage1_31[126], stage1_31[127], stage1_31[128]},
      {stage1_32[67]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], 1'b0, 1'b0},
      {stage2_35[5],stage2_34[16],stage2_33[30],stage2_32[37],stage2_31[43]}
   );
   gpc1_1 gpc1847 (
      {stage1_0[39]},
      {stage2_0[13]}
   );
   gpc1_1 gpc1848 (
      {stage1_0[40]},
      {stage2_0[14]}
   );
   gpc1_1 gpc1849 (
      {stage1_0[41]},
      {stage2_0[15]}
   );
   gpc1_1 gpc1850 (
      {stage1_0[42]},
      {stage2_0[16]}
   );
   gpc1_1 gpc1851 (
      {stage1_0[43]},
      {stage2_0[17]}
   );
   gpc1_1 gpc1852 (
      {stage1_0[44]},
      {stage2_0[18]}
   );
   gpc1_1 gpc1853 (
      {stage1_0[45]},
      {stage2_0[19]}
   );
   gpc1_1 gpc1854 (
      {stage1_0[46]},
      {stage2_0[20]}
   );
   gpc1_1 gpc1855 (
      {stage1_0[47]},
      {stage2_0[21]}
   );
   gpc1_1 gpc1856 (
      {stage1_0[48]},
      {stage2_0[22]}
   );
   gpc1_1 gpc1857 (
      {stage1_0[49]},
      {stage2_0[23]}
   );
   gpc1_1 gpc1858 (
      {stage1_1[78]},
      {stage2_1[13]}
   );
   gpc1_1 gpc1859 (
      {stage1_1[79]},
      {stage2_1[14]}
   );
   gpc1_1 gpc1860 (
      {stage1_1[80]},
      {stage2_1[15]}
   );
   gpc1_1 gpc1861 (
      {stage1_1[81]},
      {stage2_1[16]}
   );
   gpc1_1 gpc1862 (
      {stage1_1[82]},
      {stage2_1[17]}
   );
   gpc1_1 gpc1863 (
      {stage1_1[83]},
      {stage2_1[18]}
   );
   gpc1_1 gpc1864 (
      {stage1_1[84]},
      {stage2_1[19]}
   );
   gpc1_1 gpc1865 (
      {stage1_1[85]},
      {stage2_1[20]}
   );
   gpc1_1 gpc1866 (
      {stage1_1[86]},
      {stage2_1[21]}
   );
   gpc1_1 gpc1867 (
      {stage1_1[87]},
      {stage2_1[22]}
   );
   gpc1_1 gpc1868 (
      {stage1_1[88]},
      {stage2_1[23]}
   );
   gpc1_1 gpc1869 (
      {stage1_1[89]},
      {stage2_1[24]}
   );
   gpc1_1 gpc1870 (
      {stage1_1[90]},
      {stage2_1[25]}
   );
   gpc1_1 gpc1871 (
      {stage1_1[91]},
      {stage2_1[26]}
   );
   gpc1_1 gpc1872 (
      {stage1_1[92]},
      {stage2_1[27]}
   );
   gpc1_1 gpc1873 (
      {stage1_1[93]},
      {stage2_1[28]}
   );
   gpc1_1 gpc1874 (
      {stage1_1[94]},
      {stage2_1[29]}
   );
   gpc1_1 gpc1875 (
      {stage1_1[95]},
      {stage2_1[30]}
   );
   gpc1_1 gpc1876 (
      {stage1_1[96]},
      {stage2_1[31]}
   );
   gpc1_1 gpc1877 (
      {stage1_1[97]},
      {stage2_1[32]}
   );
   gpc1_1 gpc1878 (
      {stage1_2[84]},
      {stage2_2[27]}
   );
   gpc1_1 gpc1879 (
      {stage1_2[85]},
      {stage2_2[28]}
   );
   gpc1_1 gpc1880 (
      {stage1_2[86]},
      {stage2_2[29]}
   );
   gpc1_1 gpc1881 (
      {stage1_2[87]},
      {stage2_2[30]}
   );
   gpc1_1 gpc1882 (
      {stage1_2[88]},
      {stage2_2[31]}
   );
   gpc1_1 gpc1883 (
      {stage1_2[89]},
      {stage2_2[32]}
   );
   gpc1_1 gpc1884 (
      {stage1_2[90]},
      {stage2_2[33]}
   );
   gpc1_1 gpc1885 (
      {stage1_2[91]},
      {stage2_2[34]}
   );
   gpc1_1 gpc1886 (
      {stage1_3[87]},
      {stage2_3[39]}
   );
   gpc1_1 gpc1887 (
      {stage1_3[88]},
      {stage2_3[40]}
   );
   gpc1_1 gpc1888 (
      {stage1_3[89]},
      {stage2_3[41]}
   );
   gpc1_1 gpc1889 (
      {stage1_3[90]},
      {stage2_3[42]}
   );
   gpc1_1 gpc1890 (
      {stage1_4[118]},
      {stage2_4[43]}
   );
   gpc1_1 gpc1891 (
      {stage1_4[119]},
      {stage2_4[44]}
   );
   gpc1_1 gpc1892 (
      {stage1_4[120]},
      {stage2_4[45]}
   );
   gpc1_1 gpc1893 (
      {stage1_4[121]},
      {stage2_4[46]}
   );
   gpc1_1 gpc1894 (
      {stage1_4[122]},
      {stage2_4[47]}
   );
   gpc1_1 gpc1895 (
      {stage1_4[123]},
      {stage2_4[48]}
   );
   gpc1_1 gpc1896 (
      {stage1_4[124]},
      {stage2_4[49]}
   );
   gpc1_1 gpc1897 (
      {stage1_4[125]},
      {stage2_4[50]}
   );
   gpc1_1 gpc1898 (
      {stage1_4[126]},
      {stage2_4[51]}
   );
   gpc1_1 gpc1899 (
      {stage1_4[127]},
      {stage2_4[52]}
   );
   gpc1_1 gpc1900 (
      {stage1_4[128]},
      {stage2_4[53]}
   );
   gpc1_1 gpc1901 (
      {stage1_4[129]},
      {stage2_4[54]}
   );
   gpc1_1 gpc1902 (
      {stage1_4[130]},
      {stage2_4[55]}
   );
   gpc1_1 gpc1903 (
      {stage1_4[131]},
      {stage2_4[56]}
   );
   gpc1_1 gpc1904 (
      {stage1_4[132]},
      {stage2_4[57]}
   );
   gpc1_1 gpc1905 (
      {stage1_4[133]},
      {stage2_4[58]}
   );
   gpc1_1 gpc1906 (
      {stage1_4[134]},
      {stage2_4[59]}
   );
   gpc1_1 gpc1907 (
      {stage1_4[135]},
      {stage2_4[60]}
   );
   gpc1_1 gpc1908 (
      {stage1_4[136]},
      {stage2_4[61]}
   );
   gpc1_1 gpc1909 (
      {stage1_4[137]},
      {stage2_4[62]}
   );
   gpc1_1 gpc1910 (
      {stage1_4[138]},
      {stage2_4[63]}
   );
   gpc1_1 gpc1911 (
      {stage1_4[139]},
      {stage2_4[64]}
   );
   gpc1_1 gpc1912 (
      {stage1_4[140]},
      {stage2_4[65]}
   );
   gpc1_1 gpc1913 (
      {stage1_4[141]},
      {stage2_4[66]}
   );
   gpc1_1 gpc1914 (
      {stage1_4[142]},
      {stage2_4[67]}
   );
   gpc1_1 gpc1915 (
      {stage1_4[143]},
      {stage2_4[68]}
   );
   gpc1_1 gpc1916 (
      {stage1_4[144]},
      {stage2_4[69]}
   );
   gpc1_1 gpc1917 (
      {stage1_4[145]},
      {stage2_4[70]}
   );
   gpc1_1 gpc1918 (
      {stage1_4[146]},
      {stage2_4[71]}
   );
   gpc1_1 gpc1919 (
      {stage1_4[147]},
      {stage2_4[72]}
   );
   gpc1_1 gpc1920 (
      {stage1_4[148]},
      {stage2_4[73]}
   );
   gpc1_1 gpc1921 (
      {stage1_5[122]},
      {stage2_5[38]}
   );
   gpc1_1 gpc1922 (
      {stage1_5[123]},
      {stage2_5[39]}
   );
   gpc1_1 gpc1923 (
      {stage1_5[124]},
      {stage2_5[40]}
   );
   gpc1_1 gpc1924 (
      {stage1_5[125]},
      {stage2_5[41]}
   );
   gpc1_1 gpc1925 (
      {stage1_7[92]},
      {stage2_7[45]}
   );
   gpc1_1 gpc1926 (
      {stage1_7[93]},
      {stage2_7[46]}
   );
   gpc1_1 gpc1927 (
      {stage1_7[94]},
      {stage2_7[47]}
   );
   gpc1_1 gpc1928 (
      {stage1_7[95]},
      {stage2_7[48]}
   );
   gpc1_1 gpc1929 (
      {stage1_7[96]},
      {stage2_7[49]}
   );
   gpc1_1 gpc1930 (
      {stage1_7[97]},
      {stage2_7[50]}
   );
   gpc1_1 gpc1931 (
      {stage1_7[98]},
      {stage2_7[51]}
   );
   gpc1_1 gpc1932 (
      {stage1_7[99]},
      {stage2_7[52]}
   );
   gpc1_1 gpc1933 (
      {stage1_7[100]},
      {stage2_7[53]}
   );
   gpc1_1 gpc1934 (
      {stage1_8[96]},
      {stage2_8[32]}
   );
   gpc1_1 gpc1935 (
      {stage1_8[97]},
      {stage2_8[33]}
   );
   gpc1_1 gpc1936 (
      {stage1_8[98]},
      {stage2_8[34]}
   );
   gpc1_1 gpc1937 (
      {stage1_8[99]},
      {stage2_8[35]}
   );
   gpc1_1 gpc1938 (
      {stage1_8[100]},
      {stage2_8[36]}
   );
   gpc1_1 gpc1939 (
      {stage1_8[101]},
      {stage2_8[37]}
   );
   gpc1_1 gpc1940 (
      {stage1_8[102]},
      {stage2_8[38]}
   );
   gpc1_1 gpc1941 (
      {stage1_8[103]},
      {stage2_8[39]}
   );
   gpc1_1 gpc1942 (
      {stage1_8[104]},
      {stage2_8[40]}
   );
   gpc1_1 gpc1943 (
      {stage1_8[105]},
      {stage2_8[41]}
   );
   gpc1_1 gpc1944 (
      {stage1_8[106]},
      {stage2_8[42]}
   );
   gpc1_1 gpc1945 (
      {stage1_8[107]},
      {stage2_8[43]}
   );
   gpc1_1 gpc1946 (
      {stage1_8[108]},
      {stage2_8[44]}
   );
   gpc1_1 gpc1947 (
      {stage1_8[109]},
      {stage2_8[45]}
   );
   gpc1_1 gpc1948 (
      {stage1_8[110]},
      {stage2_8[46]}
   );
   gpc1_1 gpc1949 (
      {stage1_8[111]},
      {stage2_8[47]}
   );
   gpc1_1 gpc1950 (
      {stage1_8[112]},
      {stage2_8[48]}
   );
   gpc1_1 gpc1951 (
      {stage1_8[113]},
      {stage2_8[49]}
   );
   gpc1_1 gpc1952 (
      {stage1_8[114]},
      {stage2_8[50]}
   );
   gpc1_1 gpc1953 (
      {stage1_8[115]},
      {stage2_8[51]}
   );
   gpc1_1 gpc1954 (
      {stage1_8[116]},
      {stage2_8[52]}
   );
   gpc1_1 gpc1955 (
      {stage1_8[117]},
      {stage2_8[53]}
   );
   gpc1_1 gpc1956 (
      {stage1_8[118]},
      {stage2_8[54]}
   );
   gpc1_1 gpc1957 (
      {stage1_8[119]},
      {stage2_8[55]}
   );
   gpc1_1 gpc1958 (
      {stage1_9[107]},
      {stage2_9[41]}
   );
   gpc1_1 gpc1959 (
      {stage1_9[108]},
      {stage2_9[42]}
   );
   gpc1_1 gpc1960 (
      {stage1_9[109]},
      {stage2_9[43]}
   );
   gpc1_1 gpc1961 (
      {stage1_9[110]},
      {stage2_9[44]}
   );
   gpc1_1 gpc1962 (
      {stage1_9[111]},
      {stage2_9[45]}
   );
   gpc1_1 gpc1963 (
      {stage1_9[112]},
      {stage2_9[46]}
   );
   gpc1_1 gpc1964 (
      {stage1_9[113]},
      {stage2_9[47]}
   );
   gpc1_1 gpc1965 (
      {stage1_9[114]},
      {stage2_9[48]}
   );
   gpc1_1 gpc1966 (
      {stage1_9[115]},
      {stage2_9[49]}
   );
   gpc1_1 gpc1967 (
      {stage1_9[116]},
      {stage2_9[50]}
   );
   gpc1_1 gpc1968 (
      {stage1_9[117]},
      {stage2_9[51]}
   );
   gpc1_1 gpc1969 (
      {stage1_9[118]},
      {stage2_9[52]}
   );
   gpc1_1 gpc1970 (
      {stage1_9[119]},
      {stage2_9[53]}
   );
   gpc1_1 gpc1971 (
      {stage1_9[120]},
      {stage2_9[54]}
   );
   gpc1_1 gpc1972 (
      {stage1_9[121]},
      {stage2_9[55]}
   );
   gpc1_1 gpc1973 (
      {stage1_9[122]},
      {stage2_9[56]}
   );
   gpc1_1 gpc1974 (
      {stage1_9[123]},
      {stage2_9[57]}
   );
   gpc1_1 gpc1975 (
      {stage1_9[124]},
      {stage2_9[58]}
   );
   gpc1_1 gpc1976 (
      {stage1_9[125]},
      {stage2_9[59]}
   );
   gpc1_1 gpc1977 (
      {stage1_9[126]},
      {stage2_9[60]}
   );
   gpc1_1 gpc1978 (
      {stage1_9[127]},
      {stage2_9[61]}
   );
   gpc1_1 gpc1979 (
      {stage1_9[128]},
      {stage2_9[62]}
   );
   gpc1_1 gpc1980 (
      {stage1_9[129]},
      {stage2_9[63]}
   );
   gpc1_1 gpc1981 (
      {stage1_9[130]},
      {stage2_9[64]}
   );
   gpc1_1 gpc1982 (
      {stage1_9[131]},
      {stage2_9[65]}
   );
   gpc1_1 gpc1983 (
      {stage1_11[127]},
      {stage2_11[45]}
   );
   gpc1_1 gpc1984 (
      {stage1_11[128]},
      {stage2_11[46]}
   );
   gpc1_1 gpc1985 (
      {stage1_11[129]},
      {stage2_11[47]}
   );
   gpc1_1 gpc1986 (
      {stage1_11[130]},
      {stage2_11[48]}
   );
   gpc1_1 gpc1987 (
      {stage1_11[131]},
      {stage2_11[49]}
   );
   gpc1_1 gpc1988 (
      {stage1_11[132]},
      {stage2_11[50]}
   );
   gpc1_1 gpc1989 (
      {stage1_11[133]},
      {stage2_11[51]}
   );
   gpc1_1 gpc1990 (
      {stage1_11[134]},
      {stage2_11[52]}
   );
   gpc1_1 gpc1991 (
      {stage1_11[135]},
      {stage2_11[53]}
   );
   gpc1_1 gpc1992 (
      {stage1_11[136]},
      {stage2_11[54]}
   );
   gpc1_1 gpc1993 (
      {stage1_11[137]},
      {stage2_11[55]}
   );
   gpc1_1 gpc1994 (
      {stage1_11[138]},
      {stage2_11[56]}
   );
   gpc1_1 gpc1995 (
      {stage1_11[139]},
      {stage2_11[57]}
   );
   gpc1_1 gpc1996 (
      {stage1_12[173]},
      {stage2_12[50]}
   );
   gpc1_1 gpc1997 (
      {stage1_12[174]},
      {stage2_12[51]}
   );
   gpc1_1 gpc1998 (
      {stage1_12[175]},
      {stage2_12[52]}
   );
   gpc1_1 gpc1999 (
      {stage1_12[176]},
      {stage2_12[53]}
   );
   gpc1_1 gpc2000 (
      {stage1_12[177]},
      {stage2_12[54]}
   );
   gpc1_1 gpc2001 (
      {stage1_12[178]},
      {stage2_12[55]}
   );
   gpc1_1 gpc2002 (
      {stage1_12[179]},
      {stage2_12[56]}
   );
   gpc1_1 gpc2003 (
      {stage1_12[180]},
      {stage2_12[57]}
   );
   gpc1_1 gpc2004 (
      {stage1_12[181]},
      {stage2_12[58]}
   );
   gpc1_1 gpc2005 (
      {stage1_12[182]},
      {stage2_12[59]}
   );
   gpc1_1 gpc2006 (
      {stage1_12[183]},
      {stage2_12[60]}
   );
   gpc1_1 gpc2007 (
      {stage1_12[184]},
      {stage2_12[61]}
   );
   gpc1_1 gpc2008 (
      {stage1_12[185]},
      {stage2_12[62]}
   );
   gpc1_1 gpc2009 (
      {stage1_12[186]},
      {stage2_12[63]}
   );
   gpc1_1 gpc2010 (
      {stage1_12[187]},
      {stage2_12[64]}
   );
   gpc1_1 gpc2011 (
      {stage1_12[188]},
      {stage2_12[65]}
   );
   gpc1_1 gpc2012 (
      {stage1_12[189]},
      {stage2_12[66]}
   );
   gpc1_1 gpc2013 (
      {stage1_12[190]},
      {stage2_12[67]}
   );
   gpc1_1 gpc2014 (
      {stage1_12[191]},
      {stage2_12[68]}
   );
   gpc1_1 gpc2015 (
      {stage1_12[192]},
      {stage2_12[69]}
   );
   gpc1_1 gpc2016 (
      {stage1_12[193]},
      {stage2_12[70]}
   );
   gpc1_1 gpc2017 (
      {stage1_12[194]},
      {stage2_12[71]}
   );
   gpc1_1 gpc2018 (
      {stage1_12[195]},
      {stage2_12[72]}
   );
   gpc1_1 gpc2019 (
      {stage1_12[196]},
      {stage2_12[73]}
   );
   gpc1_1 gpc2020 (
      {stage1_12[197]},
      {stage2_12[74]}
   );
   gpc1_1 gpc2021 (
      {stage1_13[90]},
      {stage2_13[54]}
   );
   gpc1_1 gpc2022 (
      {stage1_13[91]},
      {stage2_13[55]}
   );
   gpc1_1 gpc2023 (
      {stage1_13[92]},
      {stage2_13[56]}
   );
   gpc1_1 gpc2024 (
      {stage1_14[66]},
      {stage2_14[42]}
   );
   gpc1_1 gpc2025 (
      {stage1_14[67]},
      {stage2_14[43]}
   );
   gpc1_1 gpc2026 (
      {stage1_14[68]},
      {stage2_14[44]}
   );
   gpc1_1 gpc2027 (
      {stage1_14[69]},
      {stage2_14[45]}
   );
   gpc1_1 gpc2028 (
      {stage1_14[70]},
      {stage2_14[46]}
   );
   gpc1_1 gpc2029 (
      {stage1_14[71]},
      {stage2_14[47]}
   );
   gpc1_1 gpc2030 (
      {stage1_14[72]},
      {stage2_14[48]}
   );
   gpc1_1 gpc2031 (
      {stage1_14[73]},
      {stage2_14[49]}
   );
   gpc1_1 gpc2032 (
      {stage1_14[74]},
      {stage2_14[50]}
   );
   gpc1_1 gpc2033 (
      {stage1_14[75]},
      {stage2_14[51]}
   );
   gpc1_1 gpc2034 (
      {stage1_14[76]},
      {stage2_14[52]}
   );
   gpc1_1 gpc2035 (
      {stage1_14[77]},
      {stage2_14[53]}
   );
   gpc1_1 gpc2036 (
      {stage1_14[78]},
      {stage2_14[54]}
   );
   gpc1_1 gpc2037 (
      {stage1_14[79]},
      {stage2_14[55]}
   );
   gpc1_1 gpc2038 (
      {stage1_14[80]},
      {stage2_14[56]}
   );
   gpc1_1 gpc2039 (
      {stage1_14[81]},
      {stage2_14[57]}
   );
   gpc1_1 gpc2040 (
      {stage1_14[82]},
      {stage2_14[58]}
   );
   gpc1_1 gpc2041 (
      {stage1_14[83]},
      {stage2_14[59]}
   );
   gpc1_1 gpc2042 (
      {stage1_14[84]},
      {stage2_14[60]}
   );
   gpc1_1 gpc2043 (
      {stage1_14[85]},
      {stage2_14[61]}
   );
   gpc1_1 gpc2044 (
      {stage1_14[86]},
      {stage2_14[62]}
   );
   gpc1_1 gpc2045 (
      {stage1_14[87]},
      {stage2_14[63]}
   );
   gpc1_1 gpc2046 (
      {stage1_14[88]},
      {stage2_14[64]}
   );
   gpc1_1 gpc2047 (
      {stage1_14[89]},
      {stage2_14[65]}
   );
   gpc1_1 gpc2048 (
      {stage1_14[90]},
      {stage2_14[66]}
   );
   gpc1_1 gpc2049 (
      {stage1_14[91]},
      {stage2_14[67]}
   );
   gpc1_1 gpc2050 (
      {stage1_14[92]},
      {stage2_14[68]}
   );
   gpc1_1 gpc2051 (
      {stage1_14[93]},
      {stage2_14[69]}
   );
   gpc1_1 gpc2052 (
      {stage1_14[94]},
      {stage2_14[70]}
   );
   gpc1_1 gpc2053 (
      {stage1_14[95]},
      {stage2_14[71]}
   );
   gpc1_1 gpc2054 (
      {stage1_14[96]},
      {stage2_14[72]}
   );
   gpc1_1 gpc2055 (
      {stage1_14[97]},
      {stage2_14[73]}
   );
   gpc1_1 gpc2056 (
      {stage1_14[98]},
      {stage2_14[74]}
   );
   gpc1_1 gpc2057 (
      {stage1_14[99]},
      {stage2_14[75]}
   );
   gpc1_1 gpc2058 (
      {stage1_14[100]},
      {stage2_14[76]}
   );
   gpc1_1 gpc2059 (
      {stage1_14[101]},
      {stage2_14[77]}
   );
   gpc1_1 gpc2060 (
      {stage1_14[102]},
      {stage2_14[78]}
   );
   gpc1_1 gpc2061 (
      {stage1_14[103]},
      {stage2_14[79]}
   );
   gpc1_1 gpc2062 (
      {stage1_14[104]},
      {stage2_14[80]}
   );
   gpc1_1 gpc2063 (
      {stage1_14[105]},
      {stage2_14[81]}
   );
   gpc1_1 gpc2064 (
      {stage1_14[106]},
      {stage2_14[82]}
   );
   gpc1_1 gpc2065 (
      {stage1_14[107]},
      {stage2_14[83]}
   );
   gpc1_1 gpc2066 (
      {stage1_14[108]},
      {stage2_14[84]}
   );
   gpc1_1 gpc2067 (
      {stage1_14[109]},
      {stage2_14[85]}
   );
   gpc1_1 gpc2068 (
      {stage1_14[110]},
      {stage2_14[86]}
   );
   gpc1_1 gpc2069 (
      {stage1_14[111]},
      {stage2_14[87]}
   );
   gpc1_1 gpc2070 (
      {stage1_14[112]},
      {stage2_14[88]}
   );
   gpc1_1 gpc2071 (
      {stage1_14[113]},
      {stage2_14[89]}
   );
   gpc1_1 gpc2072 (
      {stage1_15[84]},
      {stage2_15[38]}
   );
   gpc1_1 gpc2073 (
      {stage1_15[85]},
      {stage2_15[39]}
   );
   gpc1_1 gpc2074 (
      {stage1_15[86]},
      {stage2_15[40]}
   );
   gpc1_1 gpc2075 (
      {stage1_15[87]},
      {stage2_15[41]}
   );
   gpc1_1 gpc2076 (
      {stage1_15[88]},
      {stage2_15[42]}
   );
   gpc1_1 gpc2077 (
      {stage1_15[89]},
      {stage2_15[43]}
   );
   gpc1_1 gpc2078 (
      {stage1_15[90]},
      {stage2_15[44]}
   );
   gpc1_1 gpc2079 (
      {stage1_15[91]},
      {stage2_15[45]}
   );
   gpc1_1 gpc2080 (
      {stage1_15[92]},
      {stage2_15[46]}
   );
   gpc1_1 gpc2081 (
      {stage1_17[108]},
      {stage2_17[36]}
   );
   gpc1_1 gpc2082 (
      {stage1_17[109]},
      {stage2_17[37]}
   );
   gpc1_1 gpc2083 (
      {stage1_17[110]},
      {stage2_17[38]}
   );
   gpc1_1 gpc2084 (
      {stage1_17[111]},
      {stage2_17[39]}
   );
   gpc1_1 gpc2085 (
      {stage1_17[112]},
      {stage2_17[40]}
   );
   gpc1_1 gpc2086 (
      {stage1_17[113]},
      {stage2_17[41]}
   );
   gpc1_1 gpc2087 (
      {stage1_17[114]},
      {stage2_17[42]}
   );
   gpc1_1 gpc2088 (
      {stage1_17[115]},
      {stage2_17[43]}
   );
   gpc1_1 gpc2089 (
      {stage1_17[116]},
      {stage2_17[44]}
   );
   gpc1_1 gpc2090 (
      {stage1_17[117]},
      {stage2_17[45]}
   );
   gpc1_1 gpc2091 (
      {stage1_17[118]},
      {stage2_17[46]}
   );
   gpc1_1 gpc2092 (
      {stage1_17[119]},
      {stage2_17[47]}
   );
   gpc1_1 gpc2093 (
      {stage1_17[120]},
      {stage2_17[48]}
   );
   gpc1_1 gpc2094 (
      {stage1_17[121]},
      {stage2_17[49]}
   );
   gpc1_1 gpc2095 (
      {stage1_17[122]},
      {stage2_17[50]}
   );
   gpc1_1 gpc2096 (
      {stage1_17[123]},
      {stage2_17[51]}
   );
   gpc1_1 gpc2097 (
      {stage1_17[124]},
      {stage2_17[52]}
   );
   gpc1_1 gpc2098 (
      {stage1_17[125]},
      {stage2_17[53]}
   );
   gpc1_1 gpc2099 (
      {stage1_17[126]},
      {stage2_17[54]}
   );
   gpc1_1 gpc2100 (
      {stage1_18[94]},
      {stage2_18[34]}
   );
   gpc1_1 gpc2101 (
      {stage1_18[95]},
      {stage2_18[35]}
   );
   gpc1_1 gpc2102 (
      {stage1_18[96]},
      {stage2_18[36]}
   );
   gpc1_1 gpc2103 (
      {stage1_18[97]},
      {stage2_18[37]}
   );
   gpc1_1 gpc2104 (
      {stage1_18[98]},
      {stage2_18[38]}
   );
   gpc1_1 gpc2105 (
      {stage1_18[99]},
      {stage2_18[39]}
   );
   gpc1_1 gpc2106 (
      {stage1_18[100]},
      {stage2_18[40]}
   );
   gpc1_1 gpc2107 (
      {stage1_18[101]},
      {stage2_18[41]}
   );
   gpc1_1 gpc2108 (
      {stage1_18[102]},
      {stage2_18[42]}
   );
   gpc1_1 gpc2109 (
      {stage1_18[103]},
      {stage2_18[43]}
   );
   gpc1_1 gpc2110 (
      {stage1_18[104]},
      {stage2_18[44]}
   );
   gpc1_1 gpc2111 (
      {stage1_18[105]},
      {stage2_18[45]}
   );
   gpc1_1 gpc2112 (
      {stage1_18[106]},
      {stage2_18[46]}
   );
   gpc1_1 gpc2113 (
      {stage1_18[107]},
      {stage2_18[47]}
   );
   gpc1_1 gpc2114 (
      {stage1_18[108]},
      {stage2_18[48]}
   );
   gpc1_1 gpc2115 (
      {stage1_18[109]},
      {stage2_18[49]}
   );
   gpc1_1 gpc2116 (
      {stage1_18[110]},
      {stage2_18[50]}
   );
   gpc1_1 gpc2117 (
      {stage1_18[111]},
      {stage2_18[51]}
   );
   gpc1_1 gpc2118 (
      {stage1_18[112]},
      {stage2_18[52]}
   );
   gpc1_1 gpc2119 (
      {stage1_18[113]},
      {stage2_18[53]}
   );
   gpc1_1 gpc2120 (
      {stage1_18[114]},
      {stage2_18[54]}
   );
   gpc1_1 gpc2121 (
      {stage1_18[115]},
      {stage2_18[55]}
   );
   gpc1_1 gpc2122 (
      {stage1_18[116]},
      {stage2_18[56]}
   );
   gpc1_1 gpc2123 (
      {stage1_18[117]},
      {stage2_18[57]}
   );
   gpc1_1 gpc2124 (
      {stage1_18[118]},
      {stage2_18[58]}
   );
   gpc1_1 gpc2125 (
      {stage1_18[119]},
      {stage2_18[59]}
   );
   gpc1_1 gpc2126 (
      {stage1_18[120]},
      {stage2_18[60]}
   );
   gpc1_1 gpc2127 (
      {stage1_18[121]},
      {stage2_18[61]}
   );
   gpc1_1 gpc2128 (
      {stage1_18[122]},
      {stage2_18[62]}
   );
   gpc1_1 gpc2129 (
      {stage1_18[123]},
      {stage2_18[63]}
   );
   gpc1_1 gpc2130 (
      {stage1_18[124]},
      {stage2_18[64]}
   );
   gpc1_1 gpc2131 (
      {stage1_18[125]},
      {stage2_18[65]}
   );
   gpc1_1 gpc2132 (
      {stage1_18[126]},
      {stage2_18[66]}
   );
   gpc1_1 gpc2133 (
      {stage1_18[127]},
      {stage2_18[67]}
   );
   gpc1_1 gpc2134 (
      {stage1_18[128]},
      {stage2_18[68]}
   );
   gpc1_1 gpc2135 (
      {stage1_18[129]},
      {stage2_18[69]}
   );
   gpc1_1 gpc2136 (
      {stage1_18[130]},
      {stage2_18[70]}
   );
   gpc1_1 gpc2137 (
      {stage1_18[131]},
      {stage2_18[71]}
   );
   gpc1_1 gpc2138 (
      {stage1_18[132]},
      {stage2_18[72]}
   );
   gpc1_1 gpc2139 (
      {stage1_18[133]},
      {stage2_18[73]}
   );
   gpc1_1 gpc2140 (
      {stage1_18[134]},
      {stage2_18[74]}
   );
   gpc1_1 gpc2141 (
      {stage1_18[135]},
      {stage2_18[75]}
   );
   gpc1_1 gpc2142 (
      {stage1_18[136]},
      {stage2_18[76]}
   );
   gpc1_1 gpc2143 (
      {stage1_18[137]},
      {stage2_18[77]}
   );
   gpc1_1 gpc2144 (
      {stage1_18[138]},
      {stage2_18[78]}
   );
   gpc1_1 gpc2145 (
      {stage1_18[139]},
      {stage2_18[79]}
   );
   gpc1_1 gpc2146 (
      {stage1_18[140]},
      {stage2_18[80]}
   );
   gpc1_1 gpc2147 (
      {stage1_18[141]},
      {stage2_18[81]}
   );
   gpc1_1 gpc2148 (
      {stage1_18[142]},
      {stage2_18[82]}
   );
   gpc1_1 gpc2149 (
      {stage1_18[143]},
      {stage2_18[83]}
   );
   gpc1_1 gpc2150 (
      {stage1_18[144]},
      {stage2_18[84]}
   );
   gpc1_1 gpc2151 (
      {stage1_18[145]},
      {stage2_18[85]}
   );
   gpc1_1 gpc2152 (
      {stage1_18[146]},
      {stage2_18[86]}
   );
   gpc1_1 gpc2153 (
      {stage1_18[147]},
      {stage2_18[87]}
   );
   gpc1_1 gpc2154 (
      {stage1_18[148]},
      {stage2_18[88]}
   );
   gpc1_1 gpc2155 (
      {stage1_18[149]},
      {stage2_18[89]}
   );
   gpc1_1 gpc2156 (
      {stage1_18[150]},
      {stage2_18[90]}
   );
   gpc1_1 gpc2157 (
      {stage1_19[93]},
      {stage2_19[45]}
   );
   gpc1_1 gpc2158 (
      {stage1_20[23]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2159 (
      {stage1_20[24]},
      {stage2_20[34]}
   );
   gpc1_1 gpc2160 (
      {stage1_20[25]},
      {stage2_20[35]}
   );
   gpc1_1 gpc2161 (
      {stage1_20[26]},
      {stage2_20[36]}
   );
   gpc1_1 gpc2162 (
      {stage1_20[27]},
      {stage2_20[37]}
   );
   gpc1_1 gpc2163 (
      {stage1_20[28]},
      {stage2_20[38]}
   );
   gpc1_1 gpc2164 (
      {stage1_20[29]},
      {stage2_20[39]}
   );
   gpc1_1 gpc2165 (
      {stage1_20[30]},
      {stage2_20[40]}
   );
   gpc1_1 gpc2166 (
      {stage1_20[31]},
      {stage2_20[41]}
   );
   gpc1_1 gpc2167 (
      {stage1_20[32]},
      {stage2_20[42]}
   );
   gpc1_1 gpc2168 (
      {stage1_20[33]},
      {stage2_20[43]}
   );
   gpc1_1 gpc2169 (
      {stage1_20[34]},
      {stage2_20[44]}
   );
   gpc1_1 gpc2170 (
      {stage1_20[35]},
      {stage2_20[45]}
   );
   gpc1_1 gpc2171 (
      {stage1_20[36]},
      {stage2_20[46]}
   );
   gpc1_1 gpc2172 (
      {stage1_20[37]},
      {stage2_20[47]}
   );
   gpc1_1 gpc2173 (
      {stage1_20[38]},
      {stage2_20[48]}
   );
   gpc1_1 gpc2174 (
      {stage1_20[39]},
      {stage2_20[49]}
   );
   gpc1_1 gpc2175 (
      {stage1_20[40]},
      {stage2_20[50]}
   );
   gpc1_1 gpc2176 (
      {stage1_20[41]},
      {stage2_20[51]}
   );
   gpc1_1 gpc2177 (
      {stage1_20[42]},
      {stage2_20[52]}
   );
   gpc1_1 gpc2178 (
      {stage1_20[43]},
      {stage2_20[53]}
   );
   gpc1_1 gpc2179 (
      {stage1_20[44]},
      {stage2_20[54]}
   );
   gpc1_1 gpc2180 (
      {stage1_20[45]},
      {stage2_20[55]}
   );
   gpc1_1 gpc2181 (
      {stage1_20[46]},
      {stage2_20[56]}
   );
   gpc1_1 gpc2182 (
      {stage1_20[47]},
      {stage2_20[57]}
   );
   gpc1_1 gpc2183 (
      {stage1_20[48]},
      {stage2_20[58]}
   );
   gpc1_1 gpc2184 (
      {stage1_20[49]},
      {stage2_20[59]}
   );
   gpc1_1 gpc2185 (
      {stage1_20[50]},
      {stage2_20[60]}
   );
   gpc1_1 gpc2186 (
      {stage1_20[51]},
      {stage2_20[61]}
   );
   gpc1_1 gpc2187 (
      {stage1_20[52]},
      {stage2_20[62]}
   );
   gpc1_1 gpc2188 (
      {stage1_20[53]},
      {stage2_20[63]}
   );
   gpc1_1 gpc2189 (
      {stage1_20[54]},
      {stage2_20[64]}
   );
   gpc1_1 gpc2190 (
      {stage1_20[55]},
      {stage2_20[65]}
   );
   gpc1_1 gpc2191 (
      {stage1_20[56]},
      {stage2_20[66]}
   );
   gpc1_1 gpc2192 (
      {stage1_20[57]},
      {stage2_20[67]}
   );
   gpc1_1 gpc2193 (
      {stage1_20[58]},
      {stage2_20[68]}
   );
   gpc1_1 gpc2194 (
      {stage1_20[59]},
      {stage2_20[69]}
   );
   gpc1_1 gpc2195 (
      {stage1_20[60]},
      {stage2_20[70]}
   );
   gpc1_1 gpc2196 (
      {stage1_20[61]},
      {stage2_20[71]}
   );
   gpc1_1 gpc2197 (
      {stage1_20[62]},
      {stage2_20[72]}
   );
   gpc1_1 gpc2198 (
      {stage1_20[63]},
      {stage2_20[73]}
   );
   gpc1_1 gpc2199 (
      {stage1_20[64]},
      {stage2_20[74]}
   );
   gpc1_1 gpc2200 (
      {stage1_20[65]},
      {stage2_20[75]}
   );
   gpc1_1 gpc2201 (
      {stage1_20[66]},
      {stage2_20[76]}
   );
   gpc1_1 gpc2202 (
      {stage1_20[67]},
      {stage2_20[77]}
   );
   gpc1_1 gpc2203 (
      {stage1_20[68]},
      {stage2_20[78]}
   );
   gpc1_1 gpc2204 (
      {stage1_20[69]},
      {stage2_20[79]}
   );
   gpc1_1 gpc2205 (
      {stage1_20[70]},
      {stage2_20[80]}
   );
   gpc1_1 gpc2206 (
      {stage1_20[71]},
      {stage2_20[81]}
   );
   gpc1_1 gpc2207 (
      {stage1_20[72]},
      {stage2_20[82]}
   );
   gpc1_1 gpc2208 (
      {stage1_20[73]},
      {stage2_20[83]}
   );
   gpc1_1 gpc2209 (
      {stage1_20[74]},
      {stage2_20[84]}
   );
   gpc1_1 gpc2210 (
      {stage1_20[75]},
      {stage2_20[85]}
   );
   gpc1_1 gpc2211 (
      {stage1_20[76]},
      {stage2_20[86]}
   );
   gpc1_1 gpc2212 (
      {stage1_20[77]},
      {stage2_20[87]}
   );
   gpc1_1 gpc2213 (
      {stage1_20[78]},
      {stage2_20[88]}
   );
   gpc1_1 gpc2214 (
      {stage1_20[79]},
      {stage2_20[89]}
   );
   gpc1_1 gpc2215 (
      {stage1_20[80]},
      {stage2_20[90]}
   );
   gpc1_1 gpc2216 (
      {stage1_20[81]},
      {stage2_20[91]}
   );
   gpc1_1 gpc2217 (
      {stage1_20[82]},
      {stage2_20[92]}
   );
   gpc1_1 gpc2218 (
      {stage1_20[83]},
      {stage2_20[93]}
   );
   gpc1_1 gpc2219 (
      {stage1_20[84]},
      {stage2_20[94]}
   );
   gpc1_1 gpc2220 (
      {stage1_20[85]},
      {stage2_20[95]}
   );
   gpc1_1 gpc2221 (
      {stage1_20[86]},
      {stage2_20[96]}
   );
   gpc1_1 gpc2222 (
      {stage1_20[87]},
      {stage2_20[97]}
   );
   gpc1_1 gpc2223 (
      {stage1_20[88]},
      {stage2_20[98]}
   );
   gpc1_1 gpc2224 (
      {stage1_20[89]},
      {stage2_20[99]}
   );
   gpc1_1 gpc2225 (
      {stage1_20[90]},
      {stage2_20[100]}
   );
   gpc1_1 gpc2226 (
      {stage1_20[91]},
      {stage2_20[101]}
   );
   gpc1_1 gpc2227 (
      {stage1_20[92]},
      {stage2_20[102]}
   );
   gpc1_1 gpc2228 (
      {stage1_20[93]},
      {stage2_20[103]}
   );
   gpc1_1 gpc2229 (
      {stage1_20[94]},
      {stage2_20[104]}
   );
   gpc1_1 gpc2230 (
      {stage1_20[95]},
      {stage2_20[105]}
   );
   gpc1_1 gpc2231 (
      {stage1_20[96]},
      {stage2_20[106]}
   );
   gpc1_1 gpc2232 (
      {stage1_20[97]},
      {stage2_20[107]}
   );
   gpc1_1 gpc2233 (
      {stage1_20[98]},
      {stage2_20[108]}
   );
   gpc1_1 gpc2234 (
      {stage1_20[99]},
      {stage2_20[109]}
   );
   gpc1_1 gpc2235 (
      {stage1_20[100]},
      {stage2_20[110]}
   );
   gpc1_1 gpc2236 (
      {stage1_20[101]},
      {stage2_20[111]}
   );
   gpc1_1 gpc2237 (
      {stage1_20[102]},
      {stage2_20[112]}
   );
   gpc1_1 gpc2238 (
      {stage1_20[103]},
      {stage2_20[113]}
   );
   gpc1_1 gpc2239 (
      {stage1_20[104]},
      {stage2_20[114]}
   );
   gpc1_1 gpc2240 (
      {stage1_20[105]},
      {stage2_20[115]}
   );
   gpc1_1 gpc2241 (
      {stage1_20[106]},
      {stage2_20[116]}
   );
   gpc1_1 gpc2242 (
      {stage1_20[107]},
      {stage2_20[117]}
   );
   gpc1_1 gpc2243 (
      {stage1_20[108]},
      {stage2_20[118]}
   );
   gpc1_1 gpc2244 (
      {stage1_20[109]},
      {stage2_20[119]}
   );
   gpc1_1 gpc2245 (
      {stage1_20[110]},
      {stage2_20[120]}
   );
   gpc1_1 gpc2246 (
      {stage1_20[111]},
      {stage2_20[121]}
   );
   gpc1_1 gpc2247 (
      {stage1_20[112]},
      {stage2_20[122]}
   );
   gpc1_1 gpc2248 (
      {stage1_20[113]},
      {stage2_20[123]}
   );
   gpc1_1 gpc2249 (
      {stage1_20[114]},
      {stage2_20[124]}
   );
   gpc1_1 gpc2250 (
      {stage1_20[115]},
      {stage2_20[125]}
   );
   gpc1_1 gpc2251 (
      {stage1_21[90]},
      {stage2_21[23]}
   );
   gpc1_1 gpc2252 (
      {stage1_21[91]},
      {stage2_21[24]}
   );
   gpc1_1 gpc2253 (
      {stage1_21[92]},
      {stage2_21[25]}
   );
   gpc1_1 gpc2254 (
      {stage1_21[93]},
      {stage2_21[26]}
   );
   gpc1_1 gpc2255 (
      {stage1_21[94]},
      {stage2_21[27]}
   );
   gpc1_1 gpc2256 (
      {stage1_21[95]},
      {stage2_21[28]}
   );
   gpc1_1 gpc2257 (
      {stage1_21[96]},
      {stage2_21[29]}
   );
   gpc1_1 gpc2258 (
      {stage1_21[97]},
      {stage2_21[30]}
   );
   gpc1_1 gpc2259 (
      {stage1_21[98]},
      {stage2_21[31]}
   );
   gpc1_1 gpc2260 (
      {stage1_21[99]},
      {stage2_21[32]}
   );
   gpc1_1 gpc2261 (
      {stage1_21[100]},
      {stage2_21[33]}
   );
   gpc1_1 gpc2262 (
      {stage1_21[101]},
      {stage2_21[34]}
   );
   gpc1_1 gpc2263 (
      {stage1_21[102]},
      {stage2_21[35]}
   );
   gpc1_1 gpc2264 (
      {stage1_21[103]},
      {stage2_21[36]}
   );
   gpc1_1 gpc2265 (
      {stage1_21[104]},
      {stage2_21[37]}
   );
   gpc1_1 gpc2266 (
      {stage1_21[105]},
      {stage2_21[38]}
   );
   gpc1_1 gpc2267 (
      {stage1_21[106]},
      {stage2_21[39]}
   );
   gpc1_1 gpc2268 (
      {stage1_21[107]},
      {stage2_21[40]}
   );
   gpc1_1 gpc2269 (
      {stage1_21[108]},
      {stage2_21[41]}
   );
   gpc1_1 gpc2270 (
      {stage1_21[109]},
      {stage2_21[42]}
   );
   gpc1_1 gpc2271 (
      {stage1_21[110]},
      {stage2_21[43]}
   );
   gpc1_1 gpc2272 (
      {stage1_21[111]},
      {stage2_21[44]}
   );
   gpc1_1 gpc2273 (
      {stage1_21[112]},
      {stage2_21[45]}
   );
   gpc1_1 gpc2274 (
      {stage1_21[113]},
      {stage2_21[46]}
   );
   gpc1_1 gpc2275 (
      {stage1_21[114]},
      {stage2_21[47]}
   );
   gpc1_1 gpc2276 (
      {stage1_21[115]},
      {stage2_21[48]}
   );
   gpc1_1 gpc2277 (
      {stage1_21[116]},
      {stage2_21[49]}
   );
   gpc1_1 gpc2278 (
      {stage1_21[117]},
      {stage2_21[50]}
   );
   gpc1_1 gpc2279 (
      {stage1_21[118]},
      {stage2_21[51]}
   );
   gpc1_1 gpc2280 (
      {stage1_21[119]},
      {stage2_21[52]}
   );
   gpc1_1 gpc2281 (
      {stage1_21[120]},
      {stage2_21[53]}
   );
   gpc1_1 gpc2282 (
      {stage1_21[121]},
      {stage2_21[54]}
   );
   gpc1_1 gpc2283 (
      {stage1_21[122]},
      {stage2_21[55]}
   );
   gpc1_1 gpc2284 (
      {stage1_21[123]},
      {stage2_21[56]}
   );
   gpc1_1 gpc2285 (
      {stage1_21[124]},
      {stage2_21[57]}
   );
   gpc1_1 gpc2286 (
      {stage1_21[125]},
      {stage2_21[58]}
   );
   gpc1_1 gpc2287 (
      {stage1_21[126]},
      {stage2_21[59]}
   );
   gpc1_1 gpc2288 (
      {stage1_21[127]},
      {stage2_21[60]}
   );
   gpc1_1 gpc2289 (
      {stage1_21[128]},
      {stage2_21[61]}
   );
   gpc1_1 gpc2290 (
      {stage1_21[129]},
      {stage2_21[62]}
   );
   gpc1_1 gpc2291 (
      {stage1_21[130]},
      {stage2_21[63]}
   );
   gpc1_1 gpc2292 (
      {stage1_21[131]},
      {stage2_21[64]}
   );
   gpc1_1 gpc2293 (
      {stage1_21[132]},
      {stage2_21[65]}
   );
   gpc1_1 gpc2294 (
      {stage1_21[133]},
      {stage2_21[66]}
   );
   gpc1_1 gpc2295 (
      {stage1_21[134]},
      {stage2_21[67]}
   );
   gpc1_1 gpc2296 (
      {stage1_21[135]},
      {stage2_21[68]}
   );
   gpc1_1 gpc2297 (
      {stage1_21[136]},
      {stage2_21[69]}
   );
   gpc1_1 gpc2298 (
      {stage1_21[137]},
      {stage2_21[70]}
   );
   gpc1_1 gpc2299 (
      {stage1_21[138]},
      {stage2_21[71]}
   );
   gpc1_1 gpc2300 (
      {stage1_22[77]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2301 (
      {stage1_22[78]},
      {stage2_22[31]}
   );
   gpc1_1 gpc2302 (
      {stage1_22[79]},
      {stage2_22[32]}
   );
   gpc1_1 gpc2303 (
      {stage1_22[80]},
      {stage2_22[33]}
   );
   gpc1_1 gpc2304 (
      {stage1_22[81]},
      {stage2_22[34]}
   );
   gpc1_1 gpc2305 (
      {stage1_22[82]},
      {stage2_22[35]}
   );
   gpc1_1 gpc2306 (
      {stage1_22[83]},
      {stage2_22[36]}
   );
   gpc1_1 gpc2307 (
      {stage1_22[84]},
      {stage2_22[37]}
   );
   gpc1_1 gpc2308 (
      {stage1_22[85]},
      {stage2_22[38]}
   );
   gpc1_1 gpc2309 (
      {stage1_22[86]},
      {stage2_22[39]}
   );
   gpc1_1 gpc2310 (
      {stage1_22[87]},
      {stage2_22[40]}
   );
   gpc1_1 gpc2311 (
      {stage1_22[88]},
      {stage2_22[41]}
   );
   gpc1_1 gpc2312 (
      {stage1_22[89]},
      {stage2_22[42]}
   );
   gpc1_1 gpc2313 (
      {stage1_22[90]},
      {stage2_22[43]}
   );
   gpc1_1 gpc2314 (
      {stage1_22[91]},
      {stage2_22[44]}
   );
   gpc1_1 gpc2315 (
      {stage1_22[92]},
      {stage2_22[45]}
   );
   gpc1_1 gpc2316 (
      {stage1_22[93]},
      {stage2_22[46]}
   );
   gpc1_1 gpc2317 (
      {stage1_23[73]},
      {stage2_23[36]}
   );
   gpc1_1 gpc2318 (
      {stage1_23[74]},
      {stage2_23[37]}
   );
   gpc1_1 gpc2319 (
      {stage1_23[75]},
      {stage2_23[38]}
   );
   gpc1_1 gpc2320 (
      {stage1_23[76]},
      {stage2_23[39]}
   );
   gpc1_1 gpc2321 (
      {stage1_23[77]},
      {stage2_23[40]}
   );
   gpc1_1 gpc2322 (
      {stage1_23[78]},
      {stage2_23[41]}
   );
   gpc1_1 gpc2323 (
      {stage1_23[79]},
      {stage2_23[42]}
   );
   gpc1_1 gpc2324 (
      {stage1_23[80]},
      {stage2_23[43]}
   );
   gpc1_1 gpc2325 (
      {stage1_23[81]},
      {stage2_23[44]}
   );
   gpc1_1 gpc2326 (
      {stage1_23[82]},
      {stage2_23[45]}
   );
   gpc1_1 gpc2327 (
      {stage1_23[83]},
      {stage2_23[46]}
   );
   gpc1_1 gpc2328 (
      {stage1_23[84]},
      {stage2_23[47]}
   );
   gpc1_1 gpc2329 (
      {stage1_23[85]},
      {stage2_23[48]}
   );
   gpc1_1 gpc2330 (
      {stage1_23[86]},
      {stage2_23[49]}
   );
   gpc1_1 gpc2331 (
      {stage1_23[87]},
      {stage2_23[50]}
   );
   gpc1_1 gpc2332 (
      {stage1_23[88]},
      {stage2_23[51]}
   );
   gpc1_1 gpc2333 (
      {stage1_23[89]},
      {stage2_23[52]}
   );
   gpc1_1 gpc2334 (
      {stage1_23[90]},
      {stage2_23[53]}
   );
   gpc1_1 gpc2335 (
      {stage1_23[91]},
      {stage2_23[54]}
   );
   gpc1_1 gpc2336 (
      {stage1_23[92]},
      {stage2_23[55]}
   );
   gpc1_1 gpc2337 (
      {stage1_23[93]},
      {stage2_23[56]}
   );
   gpc1_1 gpc2338 (
      {stage1_24[249]},
      {stage2_24[59]}
   );
   gpc1_1 gpc2339 (
      {stage1_24[250]},
      {stage2_24[60]}
   );
   gpc1_1 gpc2340 (
      {stage1_24[251]},
      {stage2_24[61]}
   );
   gpc1_1 gpc2341 (
      {stage1_24[252]},
      {stage2_24[62]}
   );
   gpc1_1 gpc2342 (
      {stage1_24[253]},
      {stage2_24[63]}
   );
   gpc1_1 gpc2343 (
      {stage1_25[117]},
      {stage2_25[65]}
   );
   gpc1_1 gpc2344 (
      {stage1_27[73]},
      {stage2_27[61]}
   );
   gpc1_1 gpc2345 (
      {stage1_27[74]},
      {stage2_27[62]}
   );
   gpc1_1 gpc2346 (
      {stage1_27[75]},
      {stage2_27[63]}
   );
   gpc1_1 gpc2347 (
      {stage1_27[76]},
      {stage2_27[64]}
   );
   gpc1_1 gpc2348 (
      {stage1_27[77]},
      {stage2_27[65]}
   );
   gpc1_1 gpc2349 (
      {stage1_27[78]},
      {stage2_27[66]}
   );
   gpc1_1 gpc2350 (
      {stage1_27[79]},
      {stage2_27[67]}
   );
   gpc1_1 gpc2351 (
      {stage1_27[80]},
      {stage2_27[68]}
   );
   gpc1_1 gpc2352 (
      {stage1_27[81]},
      {stage2_27[69]}
   );
   gpc1_1 gpc2353 (
      {stage1_27[82]},
      {stage2_27[70]}
   );
   gpc1_1 gpc2354 (
      {stage1_27[83]},
      {stage2_27[71]}
   );
   gpc1_1 gpc2355 (
      {stage1_27[84]},
      {stage2_27[72]}
   );
   gpc1_1 gpc2356 (
      {stage1_27[85]},
      {stage2_27[73]}
   );
   gpc1_1 gpc2357 (
      {stage1_27[86]},
      {stage2_27[74]}
   );
   gpc1_1 gpc2358 (
      {stage1_27[87]},
      {stage2_27[75]}
   );
   gpc1_1 gpc2359 (
      {stage1_27[88]},
      {stage2_27[76]}
   );
   gpc1_1 gpc2360 (
      {stage1_27[89]},
      {stage2_27[77]}
   );
   gpc1_1 gpc2361 (
      {stage1_27[90]},
      {stage2_27[78]}
   );
   gpc1_1 gpc2362 (
      {stage1_27[91]},
      {stage2_27[79]}
   );
   gpc1_1 gpc2363 (
      {stage1_27[92]},
      {stage2_27[80]}
   );
   gpc1_1 gpc2364 (
      {stage1_27[93]},
      {stage2_27[81]}
   );
   gpc1_1 gpc2365 (
      {stage1_27[94]},
      {stage2_27[82]}
   );
   gpc1_1 gpc2366 (
      {stage1_27[95]},
      {stage2_27[83]}
   );
   gpc1_1 gpc2367 (
      {stage1_27[96]},
      {stage2_27[84]}
   );
   gpc1_1 gpc2368 (
      {stage1_27[97]},
      {stage2_27[85]}
   );
   gpc1_1 gpc2369 (
      {stage1_27[98]},
      {stage2_27[86]}
   );
   gpc1_1 gpc2370 (
      {stage1_27[99]},
      {stage2_27[87]}
   );
   gpc1_1 gpc2371 (
      {stage1_27[100]},
      {stage2_27[88]}
   );
   gpc1_1 gpc2372 (
      {stage1_27[101]},
      {stage2_27[89]}
   );
   gpc1_1 gpc2373 (
      {stage1_27[102]},
      {stage2_27[90]}
   );
   gpc1_1 gpc2374 (
      {stage1_27[103]},
      {stage2_27[91]}
   );
   gpc1_1 gpc2375 (
      {stage1_27[104]},
      {stage2_27[92]}
   );
   gpc1_1 gpc2376 (
      {stage1_27[105]},
      {stage2_27[93]}
   );
   gpc1_1 gpc2377 (
      {stage1_27[106]},
      {stage2_27[94]}
   );
   gpc1_1 gpc2378 (
      {stage1_27[107]},
      {stage2_27[95]}
   );
   gpc1_1 gpc2379 (
      {stage1_28[90]},
      {stage2_28[60]}
   );
   gpc1_1 gpc2380 (
      {stage1_28[91]},
      {stage2_28[61]}
   );
   gpc1_1 gpc2381 (
      {stage1_28[92]},
      {stage2_28[62]}
   );
   gpc1_1 gpc2382 (
      {stage1_28[93]},
      {stage2_28[63]}
   );
   gpc1_1 gpc2383 (
      {stage1_28[94]},
      {stage2_28[64]}
   );
   gpc1_1 gpc2384 (
      {stage1_28[95]},
      {stage2_28[65]}
   );
   gpc1_1 gpc2385 (
      {stage1_28[96]},
      {stage2_28[66]}
   );
   gpc1_1 gpc2386 (
      {stage1_28[97]},
      {stage2_28[67]}
   );
   gpc1_1 gpc2387 (
      {stage1_28[98]},
      {stage2_28[68]}
   );
   gpc1_1 gpc2388 (
      {stage1_28[99]},
      {stage2_28[69]}
   );
   gpc1_1 gpc2389 (
      {stage1_28[100]},
      {stage2_28[70]}
   );
   gpc1_1 gpc2390 (
      {stage1_28[101]},
      {stage2_28[71]}
   );
   gpc1_1 gpc2391 (
      {stage1_31[129]},
      {stage2_31[44]}
   );
   gpc1_1 gpc2392 (
      {stage1_31[130]},
      {stage2_31[45]}
   );
   gpc1_1 gpc2393 (
      {stage1_31[131]},
      {stage2_31[46]}
   );
   gpc1_1 gpc2394 (
      {stage1_31[132]},
      {stage2_31[47]}
   );
   gpc1_1 gpc2395 (
      {stage1_32[68]},
      {stage2_32[38]}
   );
   gpc1_1 gpc2396 (
      {stage1_32[69]},
      {stage2_32[39]}
   );
   gpc1_1 gpc2397 (
      {stage1_32[70]},
      {stage2_32[40]}
   );
   gpc1_1 gpc2398 (
      {stage1_32[71]},
      {stage2_32[41]}
   );
   gpc1_1 gpc2399 (
      {stage1_32[72]},
      {stage2_32[42]}
   );
   gpc1_1 gpc2400 (
      {stage1_32[73]},
      {stage2_32[43]}
   );
   gpc117_4 gpc2401 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_1[0]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc117_4 gpc2402 (
      {stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13]},
      {stage2_1[1]},
      {stage2_2[1]},
      {stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc2403 (
      {stage2_0[14], stage2_0[15], stage2_0[16]},
      {stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7]},
      {stage2_2[2]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc2404 (
      {stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21]},
      {stage2_1[8]},
      {stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8]},
      {stage3_4[1],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc2405 (
      {stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc2406 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[3],stage3_3[5]}
   );
   gpc615_5 gpc2407 (
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[2],stage3_4[4],stage3_3[6]}
   );
   gpc615_5 gpc2408 (
      {stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[3],stage3_4[5],stage3_3[7]}
   );
   gpc606_5 gpc2409 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[4],stage3_4[6]}
   );
   gpc606_5 gpc2410 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc2411 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25], stage2_4[26]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[6],stage3_4[8]}
   );
   gpc615_5 gpc2412 (
      {stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage2_5[18]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[6],stage3_6[7],stage3_5[7],stage3_4[9]}
   );
   gpc615_5 gpc2413 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36]},
      {stage2_5[19]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[7],stage3_6[8],stage3_5[8],stage3_4[10]}
   );
   gpc615_5 gpc2414 (
      {stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage2_5[20]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[8],stage3_6[9],stage3_5[9],stage3_4[11]}
   );
   gpc615_5 gpc2415 (
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46]},
      {stage2_5[21]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[9],stage3_6[10],stage3_5[10],stage3_4[12]}
   );
   gpc615_5 gpc2416 (
      {stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51]},
      {stage2_5[22]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[10],stage3_6[11],stage3_5[11],stage3_4[13]}
   );
   gpc606_5 gpc2417 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[11],stage3_6[12],stage3_5[12]}
   );
   gpc606_5 gpc2418 (
      {stage2_5[29], stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[9],stage3_7[12],stage3_6[13],stage3_5[13]}
   );
   gpc606_5 gpc2419 (
      {stage2_5[35], stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[10],stage3_7[13],stage3_6[14],stage3_5[14]}
   );
   gpc615_5 gpc2420 (
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[3],stage3_8[11],stage3_7[14]}
   );
   gpc615_5 gpc2421 (
      {stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[4],stage3_8[12],stage3_7[15]}
   );
   gpc615_5 gpc2422 (
      {stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32]},
      {stage2_8[2]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[2],stage3_9[5],stage3_8[13],stage3_7[16]}
   );
   gpc615_5 gpc2423 (
      {stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37]},
      {stage2_8[3]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[3],stage3_9[6],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc2424 (
      {stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41], stage2_7[42]},
      {stage2_8[4]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[4],stage3_9[7],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc2425 (
      {stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage2_8[5]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[5],stage3_9[8],stage3_8[16],stage3_7[19]}
   );
   gpc623_5 gpc2426 (
      {stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[6], stage2_8[7]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[6],stage3_9[9],stage3_8[17],stage3_7[20]}
   );
   gpc606_5 gpc2427 (
      {stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[7],stage3_10[7],stage3_9[10],stage3_8[18]}
   );
   gpc606_5 gpc2428 (
      {stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[8],stage3_10[8],stage3_9[11],stage3_8[19]}
   );
   gpc606_5 gpc2429 (
      {stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[9],stage3_10[9],stage3_9[12],stage3_8[20]}
   );
   gpc606_5 gpc2430 (
      {stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30], stage2_8[31]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[10],stage3_10[10],stage3_9[13],stage3_8[21]}
   );
   gpc606_5 gpc2431 (
      {stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36], stage2_8[37]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[11],stage3_10[11],stage3_9[14],stage3_8[22]}
   );
   gpc606_5 gpc2432 (
      {stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[12],stage3_10[12],stage3_9[15],stage3_8[23]}
   );
   gpc606_5 gpc2433 (
      {stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[13],stage3_10[13],stage3_9[16],stage3_8[24]}
   );
   gpc615_5 gpc2434 (
      {stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_9[42]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[14],stage3_10[14],stage3_9[17],stage3_8[25]}
   );
   gpc606_5 gpc2435 (
      {stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[8],stage3_11[15],stage3_10[15],stage3_9[18]}
   );
   gpc606_5 gpc2436 (
      {stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[9],stage3_11[16],stage3_10[16],stage3_9[19]}
   );
   gpc606_5 gpc2437 (
      {stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[10],stage3_11[17],stage3_10[17],stage3_9[20]}
   );
   gpc615_5 gpc2438 (
      {stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage2_10[48]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[11],stage3_11[18],stage3_10[18],stage3_9[21]}
   );
   gpc615_5 gpc2439 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[4],stage3_12[12],stage3_11[19]}
   );
   gpc615_5 gpc2440 (
      {stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage2_12[1]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[5],stage3_12[13],stage3_11[20]}
   );
   gpc615_5 gpc2441 (
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_12[2]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[6],stage3_12[14],stage3_11[21]}
   );
   gpc615_5 gpc2442 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43]},
      {stage2_12[3]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[7],stage3_12[15],stage3_11[22]}
   );
   gpc615_5 gpc2443 (
      {stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48]},
      {stage2_12[4]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[8],stage3_12[16],stage3_11[23]}
   );
   gpc615_5 gpc2444 (
      {stage2_11[49], stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53]},
      {stage2_12[5]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[5],stage3_13[9],stage3_12[17],stage3_11[24]}
   );
   gpc615_5 gpc2445 (
      {stage2_11[54], stage2_11[55], stage2_11[56], stage2_11[57], 1'b0},
      {stage2_12[6]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[6],stage3_13[10],stage3_12[18],stage3_11[25]}
   );
   gpc606_5 gpc2446 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[7],stage3_14[7],stage3_13[11],stage3_12[19]}
   );
   gpc606_5 gpc2447 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[8],stage3_14[8],stage3_13[12],stage3_12[20]}
   );
   gpc606_5 gpc2448 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[9],stage3_14[9],stage3_13[13],stage3_12[21]}
   );
   gpc606_5 gpc2449 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[10],stage3_14[10],stage3_13[14],stage3_12[22]}
   );
   gpc606_5 gpc2450 (
      {stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35], stage2_12[36]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[11],stage3_14[11],stage3_13[15],stage3_12[23]}
   );
   gpc606_5 gpc2451 (
      {stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41], stage2_12[42]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[12],stage3_14[12],stage3_13[16],stage3_12[24]}
   );
   gpc606_5 gpc2452 (
      {stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47], stage2_12[48]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[13],stage3_14[13],stage3_13[17],stage3_12[25]}
   );
   gpc606_5 gpc2453 (
      {stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53], stage2_12[54]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[14],stage3_14[14],stage3_13[18],stage3_12[26]}
   );
   gpc606_5 gpc2454 (
      {stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59], stage2_12[60]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[15],stage3_14[15],stage3_13[19],stage3_12[27]}
   );
   gpc606_5 gpc2455 (
      {stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65], stage2_12[66]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[16],stage3_14[16],stage3_13[20],stage3_12[28]}
   );
   gpc606_5 gpc2456 (
      {stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[17],stage3_14[17],stage3_13[21],stage3_12[29]}
   );
   gpc615_5 gpc2457 (
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[11],stage3_15[18],stage3_14[18]}
   );
   gpc615_5 gpc2458 (
      {stage2_14[71], stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[12],stage3_15[19],stage3_14[19]}
   );
   gpc615_5 gpc2459 (
      {stage2_14[76], stage2_14[77], stage2_14[78], stage2_14[79], stage2_14[80]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[13],stage3_15[20],stage3_14[20]}
   );
   gpc615_5 gpc2460 (
      {stage2_14[81], stage2_14[82], stage2_14[83], stage2_14[84], stage2_14[85]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[14],stage3_15[21],stage3_14[21]}
   );
   gpc615_5 gpc2461 (
      {stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8]},
      {stage2_16[24]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[4],stage3_17[4],stage3_16[15],stage3_15[22]}
   );
   gpc615_5 gpc2462 (
      {stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13]},
      {stage2_16[25]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[5],stage3_17[5],stage3_16[16],stage3_15[23]}
   );
   gpc615_5 gpc2463 (
      {stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18]},
      {stage2_16[26]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[6],stage3_17[6],stage3_16[17],stage3_15[24]}
   );
   gpc615_5 gpc2464 (
      {stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage2_16[27]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[7],stage3_17[7],stage3_16[18],stage3_15[25]}
   );
   gpc615_5 gpc2465 (
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28]},
      {stage2_16[28]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[8],stage3_17[8],stage3_16[19],stage3_15[26]}
   );
   gpc615_5 gpc2466 (
      {stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_16[29]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[9],stage3_17[9],stage3_16[20],stage3_15[27]}
   );
   gpc615_5 gpc2467 (
      {stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38]},
      {stage2_16[30]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[10],stage3_17[10],stage3_16[21],stage3_15[28]}
   );
   gpc615_5 gpc2468 (
      {stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43]},
      {stage2_16[31]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[11],stage3_17[11],stage3_16[22],stage3_15[29]}
   );
   gpc606_5 gpc2469 (
      {stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35], stage2_16[36], stage2_16[37]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[8],stage3_18[12],stage3_17[12],stage3_16[23]}
   );
   gpc615_5 gpc2470 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[0]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[9],stage3_18[13]}
   );
   gpc615_5 gpc2471 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[1]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[10],stage3_18[14]}
   );
   gpc615_5 gpc2472 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[2]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[3],stage3_19[11],stage3_18[15]}
   );
   gpc615_5 gpc2473 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[3]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[4],stage3_19[12],stage3_18[16]}
   );
   gpc615_5 gpc2474 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[4]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[5],stage3_19[13],stage3_18[17]}
   );
   gpc615_5 gpc2475 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage2_19[5]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[6],stage3_19[14],stage3_18[18]}
   );
   gpc615_5 gpc2476 (
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40]},
      {stage2_19[6]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[7],stage3_19[15],stage3_18[19]}
   );
   gpc615_5 gpc2477 (
      {stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45]},
      {stage2_19[7]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[7],stage3_20[8],stage3_19[16],stage3_18[20]}
   );
   gpc615_5 gpc2478 (
      {stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50]},
      {stage2_19[8]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[8],stage3_20[9],stage3_19[17],stage3_18[21]}
   );
   gpc615_5 gpc2479 (
      {stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55]},
      {stage2_19[9]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[9],stage3_20[10],stage3_19[18],stage3_18[22]}
   );
   gpc615_5 gpc2480 (
      {stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_19[10]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[10],stage3_20[11],stage3_19[19],stage3_18[23]}
   );
   gpc615_5 gpc2481 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65]},
      {stage2_19[11]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[11],stage3_21[11],stage3_20[12],stage3_19[20],stage3_18[24]}
   );
   gpc615_5 gpc2482 (
      {stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70]},
      {stage2_19[12]},
      {stage2_20[72], stage2_20[73], stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77]},
      {stage3_22[12],stage3_21[12],stage3_20[13],stage3_19[21],stage3_18[25]}
   );
   gpc615_5 gpc2483 (
      {stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74], stage2_18[75]},
      {stage2_19[13]},
      {stage2_20[78], stage2_20[79], stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83]},
      {stage3_22[13],stage3_21[13],stage3_20[14],stage3_19[22],stage3_18[26]}
   );
   gpc615_5 gpc2484 (
      {stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79], stage2_18[80]},
      {stage2_19[14]},
      {stage2_20[84], stage2_20[85], stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89]},
      {stage3_22[14],stage3_21[14],stage3_20[15],stage3_19[23],stage3_18[27]}
   );
   gpc615_5 gpc2485 (
      {stage2_19[15], stage2_19[16], stage2_19[17], stage2_19[18], stage2_19[19]},
      {stage2_20[90]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[15],stage3_21[15],stage3_20[16],stage3_19[24]}
   );
   gpc615_5 gpc2486 (
      {stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23], stage2_19[24]},
      {stage2_20[91]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[16],stage3_21[16],stage3_20[17],stage3_19[25]}
   );
   gpc615_5 gpc2487 (
      {stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_20[92]},
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage3_23[2],stage3_22[17],stage3_21[17],stage3_20[18],stage3_19[26]}
   );
   gpc615_5 gpc2488 (
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34]},
      {stage2_20[93]},
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage3_23[3],stage3_22[18],stage3_21[18],stage3_20[19],stage3_19[27]}
   );
   gpc615_5 gpc2489 (
      {stage2_19[35], stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39]},
      {stage2_20[94]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[4],stage3_22[19],stage3_21[19],stage3_20[20],stage3_19[28]}
   );
   gpc606_5 gpc2490 (
      {stage2_20[95], stage2_20[96], stage2_20[97], stage2_20[98], stage2_20[99], stage2_20[100]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[5],stage3_22[20],stage3_21[20],stage3_20[21]}
   );
   gpc606_5 gpc2491 (
      {stage2_20[101], stage2_20[102], stage2_20[103], stage2_20[104], stage2_20[105], stage2_20[106]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[6],stage3_22[21],stage3_21[21],stage3_20[22]}
   );
   gpc606_5 gpc2492 (
      {stage2_20[107], stage2_20[108], stage2_20[109], stage2_20[110], stage2_20[111], stage2_20[112]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[7],stage3_22[22],stage3_21[22],stage3_20[23]}
   );
   gpc1343_5 gpc2493 (
      {stage2_21[30], stage2_21[31], stage2_21[32]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21]},
      {stage2_23[0], stage2_23[1], stage2_23[2]},
      {stage2_24[0]},
      {stage3_25[0],stage3_24[3],stage3_23[8],stage3_22[23],stage3_21[23]}
   );
   gpc1343_5 gpc2494 (
      {stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage2_22[22], stage2_22[23], stage2_22[24], stage2_22[25]},
      {stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage2_24[1]},
      {stage3_25[1],stage3_24[4],stage3_23[9],stage3_22[24],stage3_21[24]}
   );
   gpc1343_5 gpc2495 (
      {stage2_21[36], stage2_21[37], stage2_21[38]},
      {stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_23[6], stage2_23[7], stage2_23[8]},
      {stage2_24[2]},
      {stage3_25[2],stage3_24[5],stage3_23[10],stage3_22[25],stage3_21[25]}
   );
   gpc615_5 gpc2496 (
      {stage2_21[39], stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43]},
      {stage2_22[30]},
      {stage2_23[9], stage2_23[10], stage2_23[11], stage2_23[12], stage2_23[13], stage2_23[14]},
      {stage3_25[3],stage3_24[6],stage3_23[11],stage3_22[26],stage3_21[26]}
   );
   gpc615_5 gpc2497 (
      {stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47], stage2_21[48]},
      {stage2_22[31]},
      {stage2_23[15], stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20]},
      {stage3_25[4],stage3_24[7],stage3_23[12],stage3_22[27],stage3_21[27]}
   );
   gpc615_5 gpc2498 (
      {stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage2_22[32]},
      {stage2_23[21], stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage3_25[5],stage3_24[8],stage3_23[13],stage3_22[28],stage3_21[28]}
   );
   gpc615_5 gpc2499 (
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58]},
      {stage2_22[33]},
      {stage2_23[27], stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32]},
      {stage3_25[6],stage3_24[9],stage3_23[14],stage3_22[29],stage3_21[29]}
   );
   gpc615_5 gpc2500 (
      {stage2_21[59], stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63]},
      {stage2_22[34]},
      {stage2_23[33], stage2_23[34], stage2_23[35], stage2_23[36], stage2_23[37], stage2_23[38]},
      {stage3_25[7],stage3_24[10],stage3_23[15],stage3_22[30],stage3_21[30]}
   );
   gpc615_5 gpc2501 (
      {stage2_21[64], stage2_21[65], stage2_21[66], stage2_21[67], stage2_21[68]},
      {stage2_22[35]},
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44]},
      {stage3_25[8],stage3_24[11],stage3_23[16],stage3_22[31],stage3_21[31]}
   );
   gpc615_5 gpc2502 (
      {stage2_21[69], stage2_21[70], stage2_21[71], 1'b0, 1'b0},
      {stage2_22[36]},
      {stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage3_25[9],stage3_24[12],stage3_23[17],stage3_22[32],stage3_21[32]}
   );
   gpc615_5 gpc2503 (
      {stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage2_23[51]},
      {stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6], stage2_24[7], stage2_24[8]},
      {stage3_26[0],stage3_25[10],stage3_24[13],stage3_23[18],stage3_22[33]}
   );
   gpc615_5 gpc2504 (
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46]},
      {stage2_23[52]},
      {stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13], stage2_24[14]},
      {stage3_26[1],stage3_25[11],stage3_24[14],stage3_23[19],stage3_22[34]}
   );
   gpc615_5 gpc2505 (
      {stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56], 1'b0},
      {stage2_24[15]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[2],stage3_25[12],stage3_24[15],stage3_23[20]}
   );
   gpc606_5 gpc2506 (
      {stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[3],stage3_25[13],stage3_24[16]}
   );
   gpc606_5 gpc2507 (
      {stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[2],stage3_26[4],stage3_25[14],stage3_24[17]}
   );
   gpc606_5 gpc2508 (
      {stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[3],stage3_26[5],stage3_25[15],stage3_24[18]}
   );
   gpc606_5 gpc2509 (
      {stage2_24[34], stage2_24[35], stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[4],stage3_26[6],stage3_25[16],stage3_24[19]}
   );
   gpc606_5 gpc2510 (
      {stage2_24[40], stage2_24[41], stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[5],stage3_26[7],stage3_25[17],stage3_24[20]}
   );
   gpc606_5 gpc2511 (
      {stage2_24[46], stage2_24[47], stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51]},
      {stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage3_28[5],stage3_27[6],stage3_26[8],stage3_25[18],stage3_24[21]}
   );
   gpc606_5 gpc2512 (
      {stage2_24[52], stage2_24[53], stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57]},
      {stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage3_28[6],stage3_27[7],stage3_26[9],stage3_25[19],stage3_24[22]}
   );
   gpc606_5 gpc2513 (
      {stage2_24[58], stage2_24[59], stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63]},
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage3_28[7],stage3_27[8],stage3_26[10],stage3_25[20],stage3_24[23]}
   );
   gpc606_5 gpc2514 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[8],stage3_27[9],stage3_26[11],stage3_25[21]}
   );
   gpc606_5 gpc2515 (
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[9],stage3_27[10],stage3_26[12],stage3_25[22]}
   );
   gpc606_5 gpc2516 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[10],stage3_27[11],stage3_26[13],stage3_25[23]}
   );
   gpc606_5 gpc2517 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[11],stage3_27[12],stage3_26[14],stage3_25[24]}
   );
   gpc606_5 gpc2518 (
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[12],stage3_27[13],stage3_26[15],stage3_25[25]}
   );
   gpc606_5 gpc2519 (
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage2_27[30], stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage3_29[5],stage3_28[13],stage3_27[14],stage3_26[16],stage3_25[26]}
   );
   gpc606_5 gpc2520 (
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage2_27[36], stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage3_29[6],stage3_28[14],stage3_27[15],stage3_26[17],stage3_25[27]}
   );
   gpc606_5 gpc2521 (
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46], stage2_27[47]},
      {stage3_29[7],stage3_28[15],stage3_27[16],stage3_26[18],stage3_25[28]}
   );
   gpc606_5 gpc2522 (
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53]},
      {stage3_29[8],stage3_28[16],stage3_27[17],stage3_26[19],stage3_25[29]}
   );
   gpc615_5 gpc2523 (
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_27[54]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[9],stage3_28[17],stage3_27[18],stage3_26[20]}
   );
   gpc615_5 gpc2524 (
      {stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57]},
      {stage2_27[55]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[10],stage3_28[18],stage3_27[19],stage3_26[21]}
   );
   gpc615_5 gpc2525 (
      {stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_27[56]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[11],stage3_28[19],stage3_27[20],stage3_26[22]}
   );
   gpc615_5 gpc2526 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67]},
      {stage2_27[57]},
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage3_30[3],stage3_29[12],stage3_28[20],stage3_27[21],stage3_26[23]}
   );
   gpc606_5 gpc2527 (
      {stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61], stage2_27[62], stage2_27[63]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[4],stage3_29[13],stage3_28[21],stage3_27[22]}
   );
   gpc615_5 gpc2528 (
      {stage2_27[64], stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68]},
      {stage2_28[24]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[5],stage3_29[14],stage3_28[22],stage3_27[23]}
   );
   gpc615_5 gpc2529 (
      {stage2_27[69], stage2_27[70], stage2_27[71], stage2_27[72], stage2_27[73]},
      {stage2_28[25]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[6],stage3_29[15],stage3_28[23],stage3_27[24]}
   );
   gpc615_5 gpc2530 (
      {stage2_27[74], stage2_27[75], stage2_27[76], stage2_27[77], stage2_27[78]},
      {stage2_28[26]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[7],stage3_29[16],stage3_28[24],stage3_27[25]}
   );
   gpc615_5 gpc2531 (
      {stage2_27[79], stage2_27[80], stage2_27[81], stage2_27[82], stage2_27[83]},
      {stage2_28[27]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[8],stage3_29[17],stage3_28[25],stage3_27[26]}
   );
   gpc606_5 gpc2532 (
      {stage2_28[28], stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[5],stage3_30[9],stage3_29[18],stage3_28[26]}
   );
   gpc606_5 gpc2533 (
      {stage2_28[34], stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38], stage2_28[39]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[6],stage3_30[10],stage3_29[19],stage3_28[27]}
   );
   gpc606_5 gpc2534 (
      {stage2_28[40], stage2_28[41], stage2_28[42], stage2_28[43], stage2_28[44], stage2_28[45]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[7],stage3_30[11],stage3_29[20],stage3_28[28]}
   );
   gpc606_5 gpc2535 (
      {stage2_28[46], stage2_28[47], stage2_28[48], stage2_28[49], stage2_28[50], stage2_28[51]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[8],stage3_30[12],stage3_29[21],stage3_28[29]}
   );
   gpc606_5 gpc2536 (
      {stage2_28[52], stage2_28[53], stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[9],stage3_30[13],stage3_29[22],stage3_28[30]}
   );
   gpc606_5 gpc2537 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[5],stage3_31[10],stage3_30[14],stage3_29[23]}
   );
   gpc615_5 gpc2538 (
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[6],stage3_31[11],stage3_30[15]}
   );
   gpc615_5 gpc2539 (
      {stage2_30[35], stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39]},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[7],stage3_31[12],stage3_30[16]}
   );
   gpc615_5 gpc2540 (
      {stage2_30[40], stage2_30[41], stage2_30[42], stage2_30[43], stage2_30[44]},
      {stage2_31[8]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[3],stage3_32[8],stage3_31[13],stage3_30[17]}
   );
   gpc615_5 gpc2541 (
      {stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12], stage2_31[13]},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[3],stage3_33[4],stage3_32[9],stage3_31[14]}
   );
   gpc615_5 gpc2542 (
      {stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17], stage2_31[18]},
      {stage2_32[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[4],stage3_33[5],stage3_32[10],stage3_31[15]}
   );
   gpc615_5 gpc2543 (
      {stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_32[20]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[5],stage3_33[6],stage3_32[11],stage3_31[16]}
   );
   gpc615_5 gpc2544 (
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage2_32[21]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[6],stage3_33[7],stage3_32[12],stage3_31[17]}
   );
   gpc606_5 gpc2545 (
      {stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[4],stage3_34[7],stage3_33[8],stage3_32[13]}
   );
   gpc606_5 gpc2546 (
      {stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[5],stage3_34[8],stage3_33[9],stage3_32[14]}
   );
   gpc606_5 gpc2547 (
      {stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], 1'b0},
      {stage3_36[2],stage3_35[6],stage3_34[9],stage3_33[10],stage3_32[15]}
   );
   gpc1_1 gpc2548 (
      {stage2_0[22]},
      {stage3_0[4]}
   );
   gpc1_1 gpc2549 (
      {stage2_0[23]},
      {stage3_0[5]}
   );
   gpc1_1 gpc2550 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc2551 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc2552 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc2553 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc2554 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc2555 (
      {stage2_1[14]},
      {stage3_1[9]}
   );
   gpc1_1 gpc2556 (
      {stage2_1[15]},
      {stage3_1[10]}
   );
   gpc1_1 gpc2557 (
      {stage2_1[16]},
      {stage3_1[11]}
   );
   gpc1_1 gpc2558 (
      {stage2_1[17]},
      {stage3_1[12]}
   );
   gpc1_1 gpc2559 (
      {stage2_1[18]},
      {stage3_1[13]}
   );
   gpc1_1 gpc2560 (
      {stage2_1[19]},
      {stage3_1[14]}
   );
   gpc1_1 gpc2561 (
      {stage2_1[20]},
      {stage3_1[15]}
   );
   gpc1_1 gpc2562 (
      {stage2_1[21]},
      {stage3_1[16]}
   );
   gpc1_1 gpc2563 (
      {stage2_1[22]},
      {stage3_1[17]}
   );
   gpc1_1 gpc2564 (
      {stage2_1[23]},
      {stage3_1[18]}
   );
   gpc1_1 gpc2565 (
      {stage2_1[24]},
      {stage3_1[19]}
   );
   gpc1_1 gpc2566 (
      {stage2_1[25]},
      {stage3_1[20]}
   );
   gpc1_1 gpc2567 (
      {stage2_1[26]},
      {stage3_1[21]}
   );
   gpc1_1 gpc2568 (
      {stage2_1[27]},
      {stage3_1[22]}
   );
   gpc1_1 gpc2569 (
      {stage2_1[28]},
      {stage3_1[23]}
   );
   gpc1_1 gpc2570 (
      {stage2_1[29]},
      {stage3_1[24]}
   );
   gpc1_1 gpc2571 (
      {stage2_1[30]},
      {stage3_1[25]}
   );
   gpc1_1 gpc2572 (
      {stage2_1[31]},
      {stage3_1[26]}
   );
   gpc1_1 gpc2573 (
      {stage2_1[32]},
      {stage3_1[27]}
   );
   gpc1_1 gpc2574 (
      {stage2_2[15]},
      {stage3_2[5]}
   );
   gpc1_1 gpc2575 (
      {stage2_2[16]},
      {stage3_2[6]}
   );
   gpc1_1 gpc2576 (
      {stage2_2[17]},
      {stage3_2[7]}
   );
   gpc1_1 gpc2577 (
      {stage2_2[18]},
      {stage3_2[8]}
   );
   gpc1_1 gpc2578 (
      {stage2_2[19]},
      {stage3_2[9]}
   );
   gpc1_1 gpc2579 (
      {stage2_2[20]},
      {stage3_2[10]}
   );
   gpc1_1 gpc2580 (
      {stage2_2[21]},
      {stage3_2[11]}
   );
   gpc1_1 gpc2581 (
      {stage2_2[22]},
      {stage3_2[12]}
   );
   gpc1_1 gpc2582 (
      {stage2_2[23]},
      {stage3_2[13]}
   );
   gpc1_1 gpc2583 (
      {stage2_2[24]},
      {stage3_2[14]}
   );
   gpc1_1 gpc2584 (
      {stage2_2[25]},
      {stage3_2[15]}
   );
   gpc1_1 gpc2585 (
      {stage2_2[26]},
      {stage3_2[16]}
   );
   gpc1_1 gpc2586 (
      {stage2_2[27]},
      {stage3_2[17]}
   );
   gpc1_1 gpc2587 (
      {stage2_2[28]},
      {stage3_2[18]}
   );
   gpc1_1 gpc2588 (
      {stage2_2[29]},
      {stage3_2[19]}
   );
   gpc1_1 gpc2589 (
      {stage2_2[30]},
      {stage3_2[20]}
   );
   gpc1_1 gpc2590 (
      {stage2_2[31]},
      {stage3_2[21]}
   );
   gpc1_1 gpc2591 (
      {stage2_2[32]},
      {stage3_2[22]}
   );
   gpc1_1 gpc2592 (
      {stage2_2[33]},
      {stage3_2[23]}
   );
   gpc1_1 gpc2593 (
      {stage2_2[34]},
      {stage3_2[24]}
   );
   gpc1_1 gpc2594 (
      {stage2_3[16]},
      {stage3_3[8]}
   );
   gpc1_1 gpc2595 (
      {stage2_3[17]},
      {stage3_3[9]}
   );
   gpc1_1 gpc2596 (
      {stage2_3[18]},
      {stage3_3[10]}
   );
   gpc1_1 gpc2597 (
      {stage2_3[19]},
      {stage3_3[11]}
   );
   gpc1_1 gpc2598 (
      {stage2_3[20]},
      {stage3_3[12]}
   );
   gpc1_1 gpc2599 (
      {stage2_3[21]},
      {stage3_3[13]}
   );
   gpc1_1 gpc2600 (
      {stage2_3[22]},
      {stage3_3[14]}
   );
   gpc1_1 gpc2601 (
      {stage2_3[23]},
      {stage3_3[15]}
   );
   gpc1_1 gpc2602 (
      {stage2_3[24]},
      {stage3_3[16]}
   );
   gpc1_1 gpc2603 (
      {stage2_3[25]},
      {stage3_3[17]}
   );
   gpc1_1 gpc2604 (
      {stage2_3[26]},
      {stage3_3[18]}
   );
   gpc1_1 gpc2605 (
      {stage2_3[27]},
      {stage3_3[19]}
   );
   gpc1_1 gpc2606 (
      {stage2_3[28]},
      {stage3_3[20]}
   );
   gpc1_1 gpc2607 (
      {stage2_3[29]},
      {stage3_3[21]}
   );
   gpc1_1 gpc2608 (
      {stage2_3[30]},
      {stage3_3[22]}
   );
   gpc1_1 gpc2609 (
      {stage2_3[31]},
      {stage3_3[23]}
   );
   gpc1_1 gpc2610 (
      {stage2_3[32]},
      {stage3_3[24]}
   );
   gpc1_1 gpc2611 (
      {stage2_3[33]},
      {stage3_3[25]}
   );
   gpc1_1 gpc2612 (
      {stage2_3[34]},
      {stage3_3[26]}
   );
   gpc1_1 gpc2613 (
      {stage2_3[35]},
      {stage3_3[27]}
   );
   gpc1_1 gpc2614 (
      {stage2_3[36]},
      {stage3_3[28]}
   );
   gpc1_1 gpc2615 (
      {stage2_3[37]},
      {stage3_3[29]}
   );
   gpc1_1 gpc2616 (
      {stage2_3[38]},
      {stage3_3[30]}
   );
   gpc1_1 gpc2617 (
      {stage2_3[39]},
      {stage3_3[31]}
   );
   gpc1_1 gpc2618 (
      {stage2_3[40]},
      {stage3_3[32]}
   );
   gpc1_1 gpc2619 (
      {stage2_3[41]},
      {stage3_3[33]}
   );
   gpc1_1 gpc2620 (
      {stage2_3[42]},
      {stage3_3[34]}
   );
   gpc1_1 gpc2621 (
      {stage2_4[52]},
      {stage3_4[14]}
   );
   gpc1_1 gpc2622 (
      {stage2_4[53]},
      {stage3_4[15]}
   );
   gpc1_1 gpc2623 (
      {stage2_4[54]},
      {stage3_4[16]}
   );
   gpc1_1 gpc2624 (
      {stage2_4[55]},
      {stage3_4[17]}
   );
   gpc1_1 gpc2625 (
      {stage2_4[56]},
      {stage3_4[18]}
   );
   gpc1_1 gpc2626 (
      {stage2_4[57]},
      {stage3_4[19]}
   );
   gpc1_1 gpc2627 (
      {stage2_4[58]},
      {stage3_4[20]}
   );
   gpc1_1 gpc2628 (
      {stage2_4[59]},
      {stage3_4[21]}
   );
   gpc1_1 gpc2629 (
      {stage2_4[60]},
      {stage3_4[22]}
   );
   gpc1_1 gpc2630 (
      {stage2_4[61]},
      {stage3_4[23]}
   );
   gpc1_1 gpc2631 (
      {stage2_4[62]},
      {stage3_4[24]}
   );
   gpc1_1 gpc2632 (
      {stage2_4[63]},
      {stage3_4[25]}
   );
   gpc1_1 gpc2633 (
      {stage2_4[64]},
      {stage3_4[26]}
   );
   gpc1_1 gpc2634 (
      {stage2_4[65]},
      {stage3_4[27]}
   );
   gpc1_1 gpc2635 (
      {stage2_4[66]},
      {stage3_4[28]}
   );
   gpc1_1 gpc2636 (
      {stage2_4[67]},
      {stage3_4[29]}
   );
   gpc1_1 gpc2637 (
      {stage2_4[68]},
      {stage3_4[30]}
   );
   gpc1_1 gpc2638 (
      {stage2_4[69]},
      {stage3_4[31]}
   );
   gpc1_1 gpc2639 (
      {stage2_4[70]},
      {stage3_4[32]}
   );
   gpc1_1 gpc2640 (
      {stage2_4[71]},
      {stage3_4[33]}
   );
   gpc1_1 gpc2641 (
      {stage2_4[72]},
      {stage3_4[34]}
   );
   gpc1_1 gpc2642 (
      {stage2_4[73]},
      {stage3_4[35]}
   );
   gpc1_1 gpc2643 (
      {stage2_5[41]},
      {stage3_5[15]}
   );
   gpc1_1 gpc2644 (
      {stage2_6[48]},
      {stage3_6[15]}
   );
   gpc1_1 gpc2645 (
      {stage2_6[49]},
      {stage3_6[16]}
   );
   gpc1_1 gpc2646 (
      {stage2_6[50]},
      {stage3_6[17]}
   );
   gpc1_1 gpc2647 (
      {stage2_6[51]},
      {stage3_6[18]}
   );
   gpc1_1 gpc2648 (
      {stage2_6[52]},
      {stage3_6[19]}
   );
   gpc1_1 gpc2649 (
      {stage2_7[51]},
      {stage3_7[21]}
   );
   gpc1_1 gpc2650 (
      {stage2_7[52]},
      {stage3_7[22]}
   );
   gpc1_1 gpc2651 (
      {stage2_7[53]},
      {stage3_7[23]}
   );
   gpc1_1 gpc2652 (
      {stage2_8[55]},
      {stage3_8[26]}
   );
   gpc1_1 gpc2653 (
      {stage2_12[73]},
      {stage3_12[30]}
   );
   gpc1_1 gpc2654 (
      {stage2_12[74]},
      {stage3_12[31]}
   );
   gpc1_1 gpc2655 (
      {stage2_13[42]},
      {stage3_13[22]}
   );
   gpc1_1 gpc2656 (
      {stage2_13[43]},
      {stage3_13[23]}
   );
   gpc1_1 gpc2657 (
      {stage2_13[44]},
      {stage3_13[24]}
   );
   gpc1_1 gpc2658 (
      {stage2_13[45]},
      {stage3_13[25]}
   );
   gpc1_1 gpc2659 (
      {stage2_13[46]},
      {stage3_13[26]}
   );
   gpc1_1 gpc2660 (
      {stage2_13[47]},
      {stage3_13[27]}
   );
   gpc1_1 gpc2661 (
      {stage2_13[48]},
      {stage3_13[28]}
   );
   gpc1_1 gpc2662 (
      {stage2_13[49]},
      {stage3_13[29]}
   );
   gpc1_1 gpc2663 (
      {stage2_13[50]},
      {stage3_13[30]}
   );
   gpc1_1 gpc2664 (
      {stage2_13[51]},
      {stage3_13[31]}
   );
   gpc1_1 gpc2665 (
      {stage2_13[52]},
      {stage3_13[32]}
   );
   gpc1_1 gpc2666 (
      {stage2_13[53]},
      {stage3_13[33]}
   );
   gpc1_1 gpc2667 (
      {stage2_13[54]},
      {stage3_13[34]}
   );
   gpc1_1 gpc2668 (
      {stage2_13[55]},
      {stage3_13[35]}
   );
   gpc1_1 gpc2669 (
      {stage2_13[56]},
      {stage3_13[36]}
   );
   gpc1_1 gpc2670 (
      {stage2_14[86]},
      {stage3_14[22]}
   );
   gpc1_1 gpc2671 (
      {stage2_14[87]},
      {stage3_14[23]}
   );
   gpc1_1 gpc2672 (
      {stage2_14[88]},
      {stage3_14[24]}
   );
   gpc1_1 gpc2673 (
      {stage2_14[89]},
      {stage3_14[25]}
   );
   gpc1_1 gpc2674 (
      {stage2_15[44]},
      {stage3_15[30]}
   );
   gpc1_1 gpc2675 (
      {stage2_15[45]},
      {stage3_15[31]}
   );
   gpc1_1 gpc2676 (
      {stage2_15[46]},
      {stage3_15[32]}
   );
   gpc1_1 gpc2677 (
      {stage2_16[38]},
      {stage3_16[24]}
   );
   gpc1_1 gpc2678 (
      {stage2_16[39]},
      {stage3_16[25]}
   );
   gpc1_1 gpc2679 (
      {stage2_16[40]},
      {stage3_16[26]}
   );
   gpc1_1 gpc2680 (
      {stage2_17[48]},
      {stage3_17[13]}
   );
   gpc1_1 gpc2681 (
      {stage2_17[49]},
      {stage3_17[14]}
   );
   gpc1_1 gpc2682 (
      {stage2_17[50]},
      {stage3_17[15]}
   );
   gpc1_1 gpc2683 (
      {stage2_17[51]},
      {stage3_17[16]}
   );
   gpc1_1 gpc2684 (
      {stage2_17[52]},
      {stage3_17[17]}
   );
   gpc1_1 gpc2685 (
      {stage2_17[53]},
      {stage3_17[18]}
   );
   gpc1_1 gpc2686 (
      {stage2_17[54]},
      {stage3_17[19]}
   );
   gpc1_1 gpc2687 (
      {stage2_18[81]},
      {stage3_18[28]}
   );
   gpc1_1 gpc2688 (
      {stage2_18[82]},
      {stage3_18[29]}
   );
   gpc1_1 gpc2689 (
      {stage2_18[83]},
      {stage3_18[30]}
   );
   gpc1_1 gpc2690 (
      {stage2_18[84]},
      {stage3_18[31]}
   );
   gpc1_1 gpc2691 (
      {stage2_18[85]},
      {stage3_18[32]}
   );
   gpc1_1 gpc2692 (
      {stage2_18[86]},
      {stage3_18[33]}
   );
   gpc1_1 gpc2693 (
      {stage2_18[87]},
      {stage3_18[34]}
   );
   gpc1_1 gpc2694 (
      {stage2_18[88]},
      {stage3_18[35]}
   );
   gpc1_1 gpc2695 (
      {stage2_18[89]},
      {stage3_18[36]}
   );
   gpc1_1 gpc2696 (
      {stage2_18[90]},
      {stage3_18[37]}
   );
   gpc1_1 gpc2697 (
      {stage2_19[40]},
      {stage3_19[29]}
   );
   gpc1_1 gpc2698 (
      {stage2_19[41]},
      {stage3_19[30]}
   );
   gpc1_1 gpc2699 (
      {stage2_19[42]},
      {stage3_19[31]}
   );
   gpc1_1 gpc2700 (
      {stage2_19[43]},
      {stage3_19[32]}
   );
   gpc1_1 gpc2701 (
      {stage2_19[44]},
      {stage3_19[33]}
   );
   gpc1_1 gpc2702 (
      {stage2_19[45]},
      {stage3_19[34]}
   );
   gpc1_1 gpc2703 (
      {stage2_20[113]},
      {stage3_20[24]}
   );
   gpc1_1 gpc2704 (
      {stage2_20[114]},
      {stage3_20[25]}
   );
   gpc1_1 gpc2705 (
      {stage2_20[115]},
      {stage3_20[26]}
   );
   gpc1_1 gpc2706 (
      {stage2_20[116]},
      {stage3_20[27]}
   );
   gpc1_1 gpc2707 (
      {stage2_20[117]},
      {stage3_20[28]}
   );
   gpc1_1 gpc2708 (
      {stage2_20[118]},
      {stage3_20[29]}
   );
   gpc1_1 gpc2709 (
      {stage2_20[119]},
      {stage3_20[30]}
   );
   gpc1_1 gpc2710 (
      {stage2_20[120]},
      {stage3_20[31]}
   );
   gpc1_1 gpc2711 (
      {stage2_20[121]},
      {stage3_20[32]}
   );
   gpc1_1 gpc2712 (
      {stage2_20[122]},
      {stage3_20[33]}
   );
   gpc1_1 gpc2713 (
      {stage2_20[123]},
      {stage3_20[34]}
   );
   gpc1_1 gpc2714 (
      {stage2_20[124]},
      {stage3_20[35]}
   );
   gpc1_1 gpc2715 (
      {stage2_20[125]},
      {stage3_20[36]}
   );
   gpc1_1 gpc2716 (
      {stage2_25[60]},
      {stage3_25[30]}
   );
   gpc1_1 gpc2717 (
      {stage2_25[61]},
      {stage3_25[31]}
   );
   gpc1_1 gpc2718 (
      {stage2_25[62]},
      {stage3_25[32]}
   );
   gpc1_1 gpc2719 (
      {stage2_25[63]},
      {stage3_25[33]}
   );
   gpc1_1 gpc2720 (
      {stage2_25[64]},
      {stage3_25[34]}
   );
   gpc1_1 gpc2721 (
      {stage2_25[65]},
      {stage3_25[35]}
   );
   gpc1_1 gpc2722 (
      {stage2_27[84]},
      {stage3_27[27]}
   );
   gpc1_1 gpc2723 (
      {stage2_27[85]},
      {stage3_27[28]}
   );
   gpc1_1 gpc2724 (
      {stage2_27[86]},
      {stage3_27[29]}
   );
   gpc1_1 gpc2725 (
      {stage2_27[87]},
      {stage3_27[30]}
   );
   gpc1_1 gpc2726 (
      {stage2_27[88]},
      {stage3_27[31]}
   );
   gpc1_1 gpc2727 (
      {stage2_27[89]},
      {stage3_27[32]}
   );
   gpc1_1 gpc2728 (
      {stage2_27[90]},
      {stage3_27[33]}
   );
   gpc1_1 gpc2729 (
      {stage2_27[91]},
      {stage3_27[34]}
   );
   gpc1_1 gpc2730 (
      {stage2_27[92]},
      {stage3_27[35]}
   );
   gpc1_1 gpc2731 (
      {stage2_27[93]},
      {stage3_27[36]}
   );
   gpc1_1 gpc2732 (
      {stage2_27[94]},
      {stage3_27[37]}
   );
   gpc1_1 gpc2733 (
      {stage2_27[95]},
      {stage3_27[38]}
   );
   gpc1_1 gpc2734 (
      {stage2_28[58]},
      {stage3_28[31]}
   );
   gpc1_1 gpc2735 (
      {stage2_28[59]},
      {stage3_28[32]}
   );
   gpc1_1 gpc2736 (
      {stage2_28[60]},
      {stage3_28[33]}
   );
   gpc1_1 gpc2737 (
      {stage2_28[61]},
      {stage3_28[34]}
   );
   gpc1_1 gpc2738 (
      {stage2_28[62]},
      {stage3_28[35]}
   );
   gpc1_1 gpc2739 (
      {stage2_28[63]},
      {stage3_28[36]}
   );
   gpc1_1 gpc2740 (
      {stage2_28[64]},
      {stage3_28[37]}
   );
   gpc1_1 gpc2741 (
      {stage2_28[65]},
      {stage3_28[38]}
   );
   gpc1_1 gpc2742 (
      {stage2_28[66]},
      {stage3_28[39]}
   );
   gpc1_1 gpc2743 (
      {stage2_28[67]},
      {stage3_28[40]}
   );
   gpc1_1 gpc2744 (
      {stage2_28[68]},
      {stage3_28[41]}
   );
   gpc1_1 gpc2745 (
      {stage2_28[69]},
      {stage3_28[42]}
   );
   gpc1_1 gpc2746 (
      {stage2_28[70]},
      {stage3_28[43]}
   );
   gpc1_1 gpc2747 (
      {stage2_28[71]},
      {stage3_28[44]}
   );
   gpc1_1 gpc2748 (
      {stage2_29[36]},
      {stage3_29[24]}
   );
   gpc1_1 gpc2749 (
      {stage2_29[37]},
      {stage3_29[25]}
   );
   gpc1_1 gpc2750 (
      {stage2_29[38]},
      {stage3_29[26]}
   );
   gpc1_1 gpc2751 (
      {stage2_29[39]},
      {stage3_29[27]}
   );
   gpc1_1 gpc2752 (
      {stage2_31[29]},
      {stage3_31[18]}
   );
   gpc1_1 gpc2753 (
      {stage2_31[30]},
      {stage3_31[19]}
   );
   gpc1_1 gpc2754 (
      {stage2_31[31]},
      {stage3_31[20]}
   );
   gpc1_1 gpc2755 (
      {stage2_31[32]},
      {stage3_31[21]}
   );
   gpc1_1 gpc2756 (
      {stage2_31[33]},
      {stage3_31[22]}
   );
   gpc1_1 gpc2757 (
      {stage2_31[34]},
      {stage3_31[23]}
   );
   gpc1_1 gpc2758 (
      {stage2_31[35]},
      {stage3_31[24]}
   );
   gpc1_1 gpc2759 (
      {stage2_31[36]},
      {stage3_31[25]}
   );
   gpc1_1 gpc2760 (
      {stage2_31[37]},
      {stage3_31[26]}
   );
   gpc1_1 gpc2761 (
      {stage2_31[38]},
      {stage3_31[27]}
   );
   gpc1_1 gpc2762 (
      {stage2_31[39]},
      {stage3_31[28]}
   );
   gpc1_1 gpc2763 (
      {stage2_31[40]},
      {stage3_31[29]}
   );
   gpc1_1 gpc2764 (
      {stage2_31[41]},
      {stage3_31[30]}
   );
   gpc1_1 gpc2765 (
      {stage2_31[42]},
      {stage3_31[31]}
   );
   gpc1_1 gpc2766 (
      {stage2_31[43]},
      {stage3_31[32]}
   );
   gpc1_1 gpc2767 (
      {stage2_31[44]},
      {stage3_31[33]}
   );
   gpc1_1 gpc2768 (
      {stage2_31[45]},
      {stage3_31[34]}
   );
   gpc1_1 gpc2769 (
      {stage2_31[46]},
      {stage3_31[35]}
   );
   gpc1_1 gpc2770 (
      {stage2_31[47]},
      {stage3_31[36]}
   );
   gpc1_1 gpc2771 (
      {stage2_32[40]},
      {stage3_32[16]}
   );
   gpc1_1 gpc2772 (
      {stage2_32[41]},
      {stage3_32[17]}
   );
   gpc1_1 gpc2773 (
      {stage2_32[42]},
      {stage3_32[18]}
   );
   gpc1_1 gpc2774 (
      {stage2_32[43]},
      {stage3_32[19]}
   );
   gpc1_1 gpc2775 (
      {stage2_33[24]},
      {stage3_33[11]}
   );
   gpc1_1 gpc2776 (
      {stage2_33[25]},
      {stage3_33[12]}
   );
   gpc1_1 gpc2777 (
      {stage2_33[26]},
      {stage3_33[13]}
   );
   gpc1_1 gpc2778 (
      {stage2_33[27]},
      {stage3_33[14]}
   );
   gpc1_1 gpc2779 (
      {stage2_33[28]},
      {stage3_33[15]}
   );
   gpc1_1 gpc2780 (
      {stage2_33[29]},
      {stage3_33[16]}
   );
   gpc1_1 gpc2781 (
      {stage2_33[30]},
      {stage3_33[17]}
   );
   gpc1_1 gpc2782 (
      {stage2_35[0]},
      {stage3_35[7]}
   );
   gpc1_1 gpc2783 (
      {stage2_35[1]},
      {stage3_35[8]}
   );
   gpc1_1 gpc2784 (
      {stage2_35[2]},
      {stage3_35[9]}
   );
   gpc1_1 gpc2785 (
      {stage2_35[3]},
      {stage3_35[10]}
   );
   gpc1_1 gpc2786 (
      {stage2_35[4]},
      {stage3_35[11]}
   );
   gpc1_1 gpc2787 (
      {stage2_35[5]},
      {stage3_35[12]}
   );
   gpc606_5 gpc2788 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc2789 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc2790 (
      {stage3_1[12], stage3_1[13], stage3_1[14], stage3_1[15], stage3_1[16], stage3_1[17]},
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17]},
      {stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc2791 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc2792 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[4],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc2793 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[5],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc2794 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[6],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc207_4 gpc2795 (
      {stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24]},
      {stage3_5[0], stage3_5[1]},
      {stage4_6[4],stage4_5[7],stage4_4[7],stage4_3[7]}
   );
   gpc207_4 gpc2796 (
      {stage3_3[25], stage3_3[26], stage3_3[27], stage3_3[28], stage3_3[29], stage3_3[30], stage3_3[31]},
      {stage3_5[2], stage3_5[3]},
      {stage4_6[5],stage4_5[8],stage4_4[8],stage4_3[8]}
   );
   gpc606_5 gpc2797 (
      {stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[6],stage4_5[9],stage4_4[9]}
   );
   gpc606_5 gpc2798 (
      {stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[7],stage4_5[10]}
   );
   gpc606_5 gpc2799 (
      {stage3_5[10], stage3_5[11], stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[8],stage4_5[11]}
   );
   gpc615_5 gpc2800 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[12]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[2],stage4_8[3],stage4_7[3],stage4_6[9]}
   );
   gpc615_5 gpc2801 (
      {stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage3_7[13]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[3],stage4_8[4],stage4_7[4],stage4_6[10]}
   );
   gpc135_4 gpc2802 (
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[2],stage4_9[4],stage4_8[5]}
   );
   gpc135_4 gpc2803 (
      {stage3_8[17], stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21]},
      {stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[1]},
      {stage4_11[1],stage4_10[3],stage4_9[5],stage4_8[6]}
   );
   gpc135_4 gpc2804 (
      {stage3_8[22], stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26]},
      {stage3_9[6], stage3_9[7], stage3_9[8]},
      {stage3_10[2]},
      {stage4_11[2],stage4_10[4],stage4_9[6],stage4_8[7]}
   );
   gpc606_5 gpc2805 (
      {stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[3],stage4_10[5],stage4_9[7]}
   );
   gpc606_5 gpc2806 (
      {stage3_9[15], stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[4],stage4_10[6],stage4_9[8]}
   );
   gpc615_5 gpc2807 (
      {stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[2],stage4_11[5],stage4_10[7]}
   );
   gpc615_5 gpc2808 (
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12]},
      {stage3_11[13]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[3],stage4_12[3],stage4_11[6],stage4_10[8]}
   );
   gpc615_5 gpc2809 (
      {stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17], stage3_11[18]},
      {stage3_12[12]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[2],stage4_13[4],stage4_12[4],stage4_11[7]}
   );
   gpc615_5 gpc2810 (
      {stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage3_12[13]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[3],stage4_13[5],stage4_12[5],stage4_11[8]}
   );
   gpc615_5 gpc2811 (
      {stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17], stage3_12[18]},
      {stage3_13[12]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[2],stage4_14[4],stage4_13[6],stage4_12[6]}
   );
   gpc615_5 gpc2812 (
      {stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_13[13]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[3],stage4_14[5],stage4_13[7],stage4_12[7]}
   );
   gpc615_5 gpc2813 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28]},
      {stage3_13[14]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[4],stage4_14[6],stage4_13[8],stage4_12[8]}
   );
   gpc606_5 gpc2814 (
      {stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[3],stage4_15[5],stage4_14[7],stage4_13[9]}
   );
   gpc606_5 gpc2815 (
      {stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25], stage3_13[26]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[4],stage4_15[6],stage4_14[8],stage4_13[10]}
   );
   gpc606_5 gpc2816 (
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[5],stage4_15[7],stage4_14[9]}
   );
   gpc615_5 gpc2817 (
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16]},
      {stage3_16[6]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[3],stage4_16[6],stage4_15[8]}
   );
   gpc615_5 gpc2818 (
      {stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21]},
      {stage3_16[7]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[2],stage4_17[4],stage4_16[7],stage4_15[9]}
   );
   gpc615_5 gpc2819 (
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26]},
      {stage3_16[8]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[3],stage4_17[5],stage4_16[8],stage4_15[10]}
   );
   gpc615_5 gpc2820 (
      {stage3_16[9], stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13]},
      {stage3_17[18]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[4],stage4_17[6],stage4_16[9]}
   );
   gpc615_5 gpc2821 (
      {stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17], stage3_16[18]},
      {stage3_17[19]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[5],stage4_17[7],stage4_16[10]}
   );
   gpc1163_5 gpc2822 (
      {stage3_18[12], stage3_18[13], stage3_18[14]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage3_20[0]},
      {stage3_21[0]},
      {stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[5],stage4_18[6]}
   );
   gpc1163_5 gpc2823 (
      {stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage3_20[1]},
      {stage3_21[1]},
      {stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[6],stage4_18[7]}
   );
   gpc1163_5 gpc2824 (
      {stage3_18[18], stage3_18[19], stage3_18[20]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage3_20[2]},
      {stage3_21[2]},
      {stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[7],stage4_18[8]}
   );
   gpc615_5 gpc2825 (
      {stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25]},
      {stage3_19[18]},
      {stage3_20[3], stage3_20[4], stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8]},
      {stage4_22[3],stage4_21[3],stage4_20[5],stage4_19[8],stage4_18[9]}
   );
   gpc615_5 gpc2826 (
      {stage3_18[26], stage3_18[27], stage3_18[28], stage3_18[29], stage3_18[30]},
      {stage3_19[19]},
      {stage3_20[9], stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14]},
      {stage4_22[4],stage4_21[4],stage4_20[6],stage4_19[9],stage4_18[10]}
   );
   gpc615_5 gpc2827 (
      {stage3_18[31], stage3_18[32], stage3_18[33], stage3_18[34], stage3_18[35]},
      {stage3_19[20]},
      {stage3_20[15], stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19], stage3_20[20]},
      {stage4_22[5],stage4_21[5],stage4_20[7],stage4_19[10],stage4_18[11]}
   );
   gpc615_5 gpc2828 (
      {stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25]},
      {stage3_20[21]},
      {stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6], stage3_21[7], stage3_21[8]},
      {stage4_23[0],stage4_22[6],stage4_21[6],stage4_20[8],stage4_19[11]}
   );
   gpc615_5 gpc2829 (
      {stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30]},
      {stage3_20[22]},
      {stage3_21[9], stage3_21[10], stage3_21[11], stage3_21[12], stage3_21[13], stage3_21[14]},
      {stage4_23[1],stage4_22[7],stage4_21[7],stage4_20[9],stage4_19[12]}
   );
   gpc615_5 gpc2830 (
      {stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34], 1'b0},
      {stage3_20[23]},
      {stage3_21[15], stage3_21[16], stage3_21[17], stage3_21[18], stage3_21[19], stage3_21[20]},
      {stage4_23[2],stage4_22[8],stage4_21[8],stage4_20[10],stage4_19[13]}
   );
   gpc606_5 gpc2831 (
      {stage3_20[24], stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[3],stage4_22[9],stage4_21[9],stage4_20[11]}
   );
   gpc606_5 gpc2832 (
      {stage3_21[21], stage3_21[22], stage3_21[23], stage3_21[24], stage3_21[25], stage3_21[26]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[1],stage4_23[4],stage4_22[10],stage4_21[10]}
   );
   gpc606_5 gpc2833 (
      {stage3_21[27], stage3_21[28], stage3_21[29], stage3_21[30], stage3_21[31], stage3_21[32]},
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage4_25[1],stage4_24[2],stage4_23[5],stage4_22[11],stage4_21[11]}
   );
   gpc615_5 gpc2834 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[12]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[2],stage4_24[3],stage4_23[6],stage4_22[12]}
   );
   gpc615_5 gpc2835 (
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15]},
      {stage3_23[13]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[3],stage4_24[4],stage4_23[7],stage4_22[13]}
   );
   gpc615_5 gpc2836 (
      {stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20]},
      {stage3_23[14]},
      {stage3_24[12], stage3_24[13], stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17]},
      {stage4_26[2],stage4_25[4],stage4_24[5],stage4_23[8],stage4_22[14]}
   );
   gpc615_5 gpc2837 (
      {stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24], stage3_22[25]},
      {stage3_23[15]},
      {stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23]},
      {stage4_26[3],stage4_25[5],stage4_24[6],stage4_23[9],stage4_22[15]}
   );
   gpc615_5 gpc2838 (
      {stage3_23[16], stage3_23[17], stage3_23[18], stage3_23[19], stage3_23[20]},
      {1'b0},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[4],stage4_25[6],stage4_24[7],stage4_23[10]}
   );
   gpc606_5 gpc2839 (
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[5],stage4_25[7]}
   );
   gpc606_5 gpc2840 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[2],stage4_26[6],stage4_25[8]}
   );
   gpc606_5 gpc2841 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[2],stage4_27[3],stage4_26[7],stage4_25[9]}
   );
   gpc606_5 gpc2842 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[3],stage4_27[4],stage4_26[8],stage4_25[10]}
   );
   gpc606_5 gpc2843 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[24], stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29]},
      {stage4_29[4],stage4_28[4],stage4_27[5],stage4_26[9],stage4_25[11]}
   );
   gpc606_5 gpc2844 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[5],stage4_28[5],stage4_27[6],stage4_26[10]}
   );
   gpc606_5 gpc2845 (
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[6],stage4_28[6],stage4_27[7],stage4_26[11]}
   );
   gpc615_5 gpc2846 (
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16]},
      {stage3_27[30]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[7],stage4_28[7],stage4_27[8],stage4_26[12]}
   );
   gpc615_5 gpc2847 (
      {stage3_26[17], stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21]},
      {stage3_27[31]},
      {stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23]},
      {stage4_30[3],stage4_29[8],stage4_28[8],stage4_27[9],stage4_26[13]}
   );
   gpc606_5 gpc2848 (
      {stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[0],stage4_30[4],stage4_29[9],stage4_28[9]}
   );
   gpc606_5 gpc2849 (
      {stage3_28[30], stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[1],stage4_30[5],stage4_29[10],stage4_28[10]}
   );
   gpc606_5 gpc2850 (
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[2],stage4_31[2],stage4_30[6],stage4_29[11]}
   );
   gpc606_5 gpc2851 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[3],stage4_31[3],stage4_30[7],stage4_29[12]}
   );
   gpc606_5 gpc2852 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[4],stage4_31[4],stage4_30[8],stage4_29[13]}
   );
   gpc606_5 gpc2853 (
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[3],stage4_32[5],stage4_31[5],stage4_30[9]}
   );
   gpc615_5 gpc2854 (
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22]},
      {stage3_32[6]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[1],stage4_33[4],stage4_32[6],stage4_31[6]}
   );
   gpc615_5 gpc2855 (
      {stage3_31[23], stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27]},
      {stage3_32[7]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[2],stage4_33[5],stage4_32[7],stage4_31[7]}
   );
   gpc606_5 gpc2856 (
      {stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11], stage3_32[12], stage3_32[13]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[2],stage4_34[3],stage4_33[6],stage4_32[8]}
   );
   gpc606_5 gpc2857 (
      {stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], 1'b0, 1'b0},
      {stage4_36[1],stage4_35[3],stage4_34[4],stage4_33[7],stage4_32[9]}
   );
   gpc606_5 gpc2858 (
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[2],stage4_35[4],stage4_34[5],stage4_33[8]}
   );
   gpc1_1 gpc2859 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc2860 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc2861 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc2862 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc2863 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc2864 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc2865 (
      {stage3_1[18]},
      {stage4_1[3]}
   );
   gpc1_1 gpc2866 (
      {stage3_1[19]},
      {stage4_1[4]}
   );
   gpc1_1 gpc2867 (
      {stage3_1[20]},
      {stage4_1[5]}
   );
   gpc1_1 gpc2868 (
      {stage3_1[21]},
      {stage4_1[6]}
   );
   gpc1_1 gpc2869 (
      {stage3_1[22]},
      {stage4_1[7]}
   );
   gpc1_1 gpc2870 (
      {stage3_1[23]},
      {stage4_1[8]}
   );
   gpc1_1 gpc2871 (
      {stage3_1[24]},
      {stage4_1[9]}
   );
   gpc1_1 gpc2872 (
      {stage3_1[25]},
      {stage4_1[10]}
   );
   gpc1_1 gpc2873 (
      {stage3_1[26]},
      {stage4_1[11]}
   );
   gpc1_1 gpc2874 (
      {stage3_1[27]},
      {stage4_1[12]}
   );
   gpc1_1 gpc2875 (
      {stage3_2[24]},
      {stage4_2[7]}
   );
   gpc1_1 gpc2876 (
      {stage3_3[32]},
      {stage4_3[9]}
   );
   gpc1_1 gpc2877 (
      {stage3_3[33]},
      {stage4_3[10]}
   );
   gpc1_1 gpc2878 (
      {stage3_3[34]},
      {stage4_3[11]}
   );
   gpc1_1 gpc2879 (
      {stage3_4[30]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2880 (
      {stage3_4[31]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2881 (
      {stage3_4[32]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2882 (
      {stage3_4[33]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2883 (
      {stage3_4[34]},
      {stage4_4[14]}
   );
   gpc1_1 gpc2884 (
      {stage3_4[35]},
      {stage4_4[15]}
   );
   gpc1_1 gpc2885 (
      {stage3_6[16]},
      {stage4_6[11]}
   );
   gpc1_1 gpc2886 (
      {stage3_6[17]},
      {stage4_6[12]}
   );
   gpc1_1 gpc2887 (
      {stage3_6[18]},
      {stage4_6[13]}
   );
   gpc1_1 gpc2888 (
      {stage3_6[19]},
      {stage4_6[14]}
   );
   gpc1_1 gpc2889 (
      {stage3_7[14]},
      {stage4_7[5]}
   );
   gpc1_1 gpc2890 (
      {stage3_7[15]},
      {stage4_7[6]}
   );
   gpc1_1 gpc2891 (
      {stage3_7[16]},
      {stage4_7[7]}
   );
   gpc1_1 gpc2892 (
      {stage3_7[17]},
      {stage4_7[8]}
   );
   gpc1_1 gpc2893 (
      {stage3_7[18]},
      {stage4_7[9]}
   );
   gpc1_1 gpc2894 (
      {stage3_7[19]},
      {stage4_7[10]}
   );
   gpc1_1 gpc2895 (
      {stage3_7[20]},
      {stage4_7[11]}
   );
   gpc1_1 gpc2896 (
      {stage3_7[21]},
      {stage4_7[12]}
   );
   gpc1_1 gpc2897 (
      {stage3_7[22]},
      {stage4_7[13]}
   );
   gpc1_1 gpc2898 (
      {stage3_7[23]},
      {stage4_7[14]}
   );
   gpc1_1 gpc2899 (
      {stage3_9[21]},
      {stage4_9[9]}
   );
   gpc1_1 gpc2900 (
      {stage3_10[13]},
      {stage4_10[9]}
   );
   gpc1_1 gpc2901 (
      {stage3_10[14]},
      {stage4_10[10]}
   );
   gpc1_1 gpc2902 (
      {stage3_10[15]},
      {stage4_10[11]}
   );
   gpc1_1 gpc2903 (
      {stage3_10[16]},
      {stage4_10[12]}
   );
   gpc1_1 gpc2904 (
      {stage3_10[17]},
      {stage4_10[13]}
   );
   gpc1_1 gpc2905 (
      {stage3_10[18]},
      {stage4_10[14]}
   );
   gpc1_1 gpc2906 (
      {stage3_11[24]},
      {stage4_11[9]}
   );
   gpc1_1 gpc2907 (
      {stage3_11[25]},
      {stage4_11[10]}
   );
   gpc1_1 gpc2908 (
      {stage3_12[29]},
      {stage4_12[9]}
   );
   gpc1_1 gpc2909 (
      {stage3_12[30]},
      {stage4_12[10]}
   );
   gpc1_1 gpc2910 (
      {stage3_12[31]},
      {stage4_12[11]}
   );
   gpc1_1 gpc2911 (
      {stage3_13[27]},
      {stage4_13[11]}
   );
   gpc1_1 gpc2912 (
      {stage3_13[28]},
      {stage4_13[12]}
   );
   gpc1_1 gpc2913 (
      {stage3_13[29]},
      {stage4_13[13]}
   );
   gpc1_1 gpc2914 (
      {stage3_13[30]},
      {stage4_13[14]}
   );
   gpc1_1 gpc2915 (
      {stage3_13[31]},
      {stage4_13[15]}
   );
   gpc1_1 gpc2916 (
      {stage3_13[32]},
      {stage4_13[16]}
   );
   gpc1_1 gpc2917 (
      {stage3_13[33]},
      {stage4_13[17]}
   );
   gpc1_1 gpc2918 (
      {stage3_13[34]},
      {stage4_13[18]}
   );
   gpc1_1 gpc2919 (
      {stage3_13[35]},
      {stage4_13[19]}
   );
   gpc1_1 gpc2920 (
      {stage3_13[36]},
      {stage4_13[20]}
   );
   gpc1_1 gpc2921 (
      {stage3_14[24]},
      {stage4_14[10]}
   );
   gpc1_1 gpc2922 (
      {stage3_14[25]},
      {stage4_14[11]}
   );
   gpc1_1 gpc2923 (
      {stage3_15[27]},
      {stage4_15[11]}
   );
   gpc1_1 gpc2924 (
      {stage3_15[28]},
      {stage4_15[12]}
   );
   gpc1_1 gpc2925 (
      {stage3_15[29]},
      {stage4_15[13]}
   );
   gpc1_1 gpc2926 (
      {stage3_15[30]},
      {stage4_15[14]}
   );
   gpc1_1 gpc2927 (
      {stage3_15[31]},
      {stage4_15[15]}
   );
   gpc1_1 gpc2928 (
      {stage3_15[32]},
      {stage4_15[16]}
   );
   gpc1_1 gpc2929 (
      {stage3_16[19]},
      {stage4_16[11]}
   );
   gpc1_1 gpc2930 (
      {stage3_16[20]},
      {stage4_16[12]}
   );
   gpc1_1 gpc2931 (
      {stage3_16[21]},
      {stage4_16[13]}
   );
   gpc1_1 gpc2932 (
      {stage3_16[22]},
      {stage4_16[14]}
   );
   gpc1_1 gpc2933 (
      {stage3_16[23]},
      {stage4_16[15]}
   );
   gpc1_1 gpc2934 (
      {stage3_16[24]},
      {stage4_16[16]}
   );
   gpc1_1 gpc2935 (
      {stage3_16[25]},
      {stage4_16[17]}
   );
   gpc1_1 gpc2936 (
      {stage3_16[26]},
      {stage4_16[18]}
   );
   gpc1_1 gpc2937 (
      {stage3_18[36]},
      {stage4_18[12]}
   );
   gpc1_1 gpc2938 (
      {stage3_18[37]},
      {stage4_18[13]}
   );
   gpc1_1 gpc2939 (
      {stage3_20[30]},
      {stage4_20[12]}
   );
   gpc1_1 gpc2940 (
      {stage3_20[31]},
      {stage4_20[13]}
   );
   gpc1_1 gpc2941 (
      {stage3_20[32]},
      {stage4_20[14]}
   );
   gpc1_1 gpc2942 (
      {stage3_20[33]},
      {stage4_20[15]}
   );
   gpc1_1 gpc2943 (
      {stage3_20[34]},
      {stage4_20[16]}
   );
   gpc1_1 gpc2944 (
      {stage3_20[35]},
      {stage4_20[17]}
   );
   gpc1_1 gpc2945 (
      {stage3_20[36]},
      {stage4_20[18]}
   );
   gpc1_1 gpc2946 (
      {stage3_22[26]},
      {stage4_22[16]}
   );
   gpc1_1 gpc2947 (
      {stage3_22[27]},
      {stage4_22[17]}
   );
   gpc1_1 gpc2948 (
      {stage3_22[28]},
      {stage4_22[18]}
   );
   gpc1_1 gpc2949 (
      {stage3_22[29]},
      {stage4_22[19]}
   );
   gpc1_1 gpc2950 (
      {stage3_22[30]},
      {stage4_22[20]}
   );
   gpc1_1 gpc2951 (
      {stage3_22[31]},
      {stage4_22[21]}
   );
   gpc1_1 gpc2952 (
      {stage3_22[32]},
      {stage4_22[22]}
   );
   gpc1_1 gpc2953 (
      {stage3_22[33]},
      {stage4_22[23]}
   );
   gpc1_1 gpc2954 (
      {stage3_22[34]},
      {stage4_22[24]}
   );
   gpc1_1 gpc2955 (
      {stage3_26[22]},
      {stage4_26[14]}
   );
   gpc1_1 gpc2956 (
      {stage3_26[23]},
      {stage4_26[15]}
   );
   gpc1_1 gpc2957 (
      {stage3_27[32]},
      {stage4_27[10]}
   );
   gpc1_1 gpc2958 (
      {stage3_27[33]},
      {stage4_27[11]}
   );
   gpc1_1 gpc2959 (
      {stage3_27[34]},
      {stage4_27[12]}
   );
   gpc1_1 gpc2960 (
      {stage3_27[35]},
      {stage4_27[13]}
   );
   gpc1_1 gpc2961 (
      {stage3_27[36]},
      {stage4_27[14]}
   );
   gpc1_1 gpc2962 (
      {stage3_27[37]},
      {stage4_27[15]}
   );
   gpc1_1 gpc2963 (
      {stage3_27[38]},
      {stage4_27[16]}
   );
   gpc1_1 gpc2964 (
      {stage3_28[36]},
      {stage4_28[11]}
   );
   gpc1_1 gpc2965 (
      {stage3_28[37]},
      {stage4_28[12]}
   );
   gpc1_1 gpc2966 (
      {stage3_28[38]},
      {stage4_28[13]}
   );
   gpc1_1 gpc2967 (
      {stage3_28[39]},
      {stage4_28[14]}
   );
   gpc1_1 gpc2968 (
      {stage3_28[40]},
      {stage4_28[15]}
   );
   gpc1_1 gpc2969 (
      {stage3_28[41]},
      {stage4_28[16]}
   );
   gpc1_1 gpc2970 (
      {stage3_28[42]},
      {stage4_28[17]}
   );
   gpc1_1 gpc2971 (
      {stage3_28[43]},
      {stage4_28[18]}
   );
   gpc1_1 gpc2972 (
      {stage3_28[44]},
      {stage4_28[19]}
   );
   gpc1_1 gpc2973 (
      {stage3_29[18]},
      {stage4_29[14]}
   );
   gpc1_1 gpc2974 (
      {stage3_29[19]},
      {stage4_29[15]}
   );
   gpc1_1 gpc2975 (
      {stage3_29[20]},
      {stage4_29[16]}
   );
   gpc1_1 gpc2976 (
      {stage3_29[21]},
      {stage4_29[17]}
   );
   gpc1_1 gpc2977 (
      {stage3_29[22]},
      {stage4_29[18]}
   );
   gpc1_1 gpc2978 (
      {stage3_29[23]},
      {stage4_29[19]}
   );
   gpc1_1 gpc2979 (
      {stage3_29[24]},
      {stage4_29[20]}
   );
   gpc1_1 gpc2980 (
      {stage3_29[25]},
      {stage4_29[21]}
   );
   gpc1_1 gpc2981 (
      {stage3_29[26]},
      {stage4_29[22]}
   );
   gpc1_1 gpc2982 (
      {stage3_29[27]},
      {stage4_29[23]}
   );
   gpc1_1 gpc2983 (
      {stage3_31[28]},
      {stage4_31[8]}
   );
   gpc1_1 gpc2984 (
      {stage3_31[29]},
      {stage4_31[9]}
   );
   gpc1_1 gpc2985 (
      {stage3_31[30]},
      {stage4_31[10]}
   );
   gpc1_1 gpc2986 (
      {stage3_31[31]},
      {stage4_31[11]}
   );
   gpc1_1 gpc2987 (
      {stage3_31[32]},
      {stage4_31[12]}
   );
   gpc1_1 gpc2988 (
      {stage3_31[33]},
      {stage4_31[13]}
   );
   gpc1_1 gpc2989 (
      {stage3_31[34]},
      {stage4_31[14]}
   );
   gpc1_1 gpc2990 (
      {stage3_31[35]},
      {stage4_31[15]}
   );
   gpc1_1 gpc2991 (
      {stage3_31[36]},
      {stage4_31[16]}
   );
   gpc1_1 gpc2992 (
      {stage3_35[6]},
      {stage4_35[5]}
   );
   gpc1_1 gpc2993 (
      {stage3_35[7]},
      {stage4_35[6]}
   );
   gpc1_1 gpc2994 (
      {stage3_35[8]},
      {stage4_35[7]}
   );
   gpc1_1 gpc2995 (
      {stage3_35[9]},
      {stage4_35[8]}
   );
   gpc1_1 gpc2996 (
      {stage3_35[10]},
      {stage4_35[9]}
   );
   gpc1_1 gpc2997 (
      {stage3_35[11]},
      {stage4_35[10]}
   );
   gpc1_1 gpc2998 (
      {stage3_35[12]},
      {stage4_35[11]}
   );
   gpc1_1 gpc2999 (
      {stage3_36[0]},
      {stage4_36[3]}
   );
   gpc1_1 gpc3000 (
      {stage3_36[1]},
      {stage4_36[4]}
   );
   gpc1_1 gpc3001 (
      {stage3_36[2]},
      {stage4_36[5]}
   );
   gpc606_5 gpc3002 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc3003 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc606_5 gpc3004 (
      {stage4_1[6], stage4_1[7], stage4_1[8], stage4_1[9], stage4_1[10], stage4_1[11]},
      {stage4_3[6], stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage5_5[1],stage5_4[2],stage5_3[2],stage5_2[2],stage5_1[2]}
   );
   gpc606_5 gpc3005 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[2],stage5_4[3]}
   );
   gpc606_5 gpc3006 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[3],stage5_4[4]}
   );
   gpc606_5 gpc3007 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[2],stage5_7[2],stage5_6[2],stage5_5[4]}
   );
   gpc606_5 gpc3008 (
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage5_9[1],stage5_8[3],stage5_7[3],stage5_6[3],stage5_5[5]}
   );
   gpc606_5 gpc3009 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[2],stage5_8[4]}
   );
   gpc615_5 gpc3010 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1]}
   );
   gpc606_5 gpc3011 (
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[2]}
   );
   gpc606_5 gpc3012 (
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2],stage5_12[3]}
   );
   gpc606_5 gpc3013 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[1],stage5_15[2],stage5_14[3],stage5_13[3]}
   );
   gpc606_5 gpc3014 (
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[2],stage5_15[3],stage5_14[4],stage5_13[4]}
   );
   gpc615_5 gpc3015 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[12]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[2],stage5_16[3],stage5_15[4],stage5_14[5]}
   );
   gpc207_4 gpc3016 (
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[0],stage5_18[1],stage5_17[3],stage5_16[4]}
   );
   gpc606_5 gpc3017 (
      {stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6], stage4_18[7]},
      {stage5_20[0],stage5_19[1],stage5_18[2],stage5_17[4],stage5_16[5]}
   );
   gpc606_5 gpc3018 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[2],stage5_18[3],stage5_17[5]}
   );
   gpc615_5 gpc3019 (
      {stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11], stage4_18[12]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[2],stage5_19[3],stage5_18[4]}
   );
   gpc615_5 gpc3020 (
      {stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage4_20[6]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[1],stage5_21[2],stage5_20[3],stage5_19[4]}
   );
   gpc623_5 gpc3021 (
      {stage4_20[7], stage4_20[8], stage4_20[9]},
      {stage4_21[6], stage4_21[7]},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[1],stage5_22[2],stage5_21[3],stage5_20[4]}
   );
   gpc623_5 gpc3022 (
      {stage4_20[10], stage4_20[11], stage4_20[12]},
      {stage4_21[8], stage4_21[9]},
      {stage4_22[6], stage4_22[7], stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11]},
      {stage5_24[1],stage5_23[2],stage5_22[3],stage5_21[4],stage5_20[5]}
   );
   gpc623_5 gpc3023 (
      {stage4_20[13], stage4_20[14], stage4_20[15]},
      {stage4_21[10], stage4_21[11]},
      {stage4_22[12], stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17]},
      {stage5_24[2],stage5_23[3],stage5_22[4],stage5_21[5],stage5_20[6]}
   );
   gpc615_5 gpc3024 (
      {stage4_22[18], stage4_22[19], stage4_22[20], stage4_22[21], stage4_22[22]},
      {stage4_23[0]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[0],stage5_24[3],stage5_23[4],stage5_22[5]}
   );
   gpc615_5 gpc3025 (
      {stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[6]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[1],stage5_25[1],stage5_24[4],stage5_23[5]}
   );
   gpc615_5 gpc3026 (
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10]},
      {stage4_24[7]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[2],stage5_25[2],stage5_24[5],stage5_23[6]}
   );
   gpc606_5 gpc3027 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[0],stage5_27[2],stage5_26[3]}
   );
   gpc615_5 gpc3028 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[1],stage5_28[1],stage5_27[3],stage5_26[4]}
   );
   gpc615_5 gpc3029 (
      {stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14], stage4_26[15]},
      {stage4_27[1]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[2],stage5_28[2],stage5_27[4],stage5_26[5]}
   );
   gpc615_5 gpc3030 (
      {stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[18]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[3],stage5_29[3],stage5_28[3],stage5_27[5]}
   );
   gpc615_5 gpc3031 (
      {stage4_27[7], stage4_27[8], stage4_27[9], stage4_27[10], stage4_27[11]},
      {stage4_28[19]},
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11]},
      {stage5_31[1],stage5_30[4],stage5_29[4],stage5_28[4],stage5_27[6]}
   );
   gpc615_5 gpc3032 (
      {stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {1'b0},
      {stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage5_31[2],stage5_30[5],stage5_29[5],stage5_28[5],stage5_27[7]}
   );
   gpc606_5 gpc3033 (
      {stage4_29[18], stage4_29[19], stage4_29[20], stage4_29[21], stage4_29[22], stage4_29[23]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[3],stage5_30[6],stage5_29[6]}
   );
   gpc1163_5 gpc3034 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage4_32[0]},
      {stage4_33[0]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[4],stage5_30[7]}
   );
   gpc1163_5 gpc3035 (
      {stage4_30[3], stage4_30[4], stage4_30[5]},
      {stage4_31[12], stage4_31[13], stage4_31[14], stage4_31[15], stage4_31[16], 1'b0},
      {stage4_32[1]},
      {stage4_33[1]},
      {stage5_34[1],stage5_33[2],stage5_32[2],stage5_31[5],stage5_30[8]}
   );
   gpc606_5 gpc3036 (
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[3],stage5_32[3]}
   );
   gpc606_5 gpc3037 (
      {stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5], stage4_33[6], stage4_33[7]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[4]}
   );
   gpc1_1 gpc3038 (
      {stage4_1[12]},
      {stage5_1[3]}
   );
   gpc1_1 gpc3039 (
      {stage4_2[6]},
      {stage5_2[3]}
   );
   gpc1_1 gpc3040 (
      {stage4_2[7]},
      {stage5_2[4]}
   );
   gpc1_1 gpc3041 (
      {stage4_4[12]},
      {stage5_4[5]}
   );
   gpc1_1 gpc3042 (
      {stage4_4[13]},
      {stage5_4[6]}
   );
   gpc1_1 gpc3043 (
      {stage4_4[14]},
      {stage5_4[7]}
   );
   gpc1_1 gpc3044 (
      {stage4_4[15]},
      {stage5_4[8]}
   );
   gpc1_1 gpc3045 (
      {stage4_6[12]},
      {stage5_6[4]}
   );
   gpc1_1 gpc3046 (
      {stage4_6[13]},
      {stage5_6[5]}
   );
   gpc1_1 gpc3047 (
      {stage4_6[14]},
      {stage5_6[6]}
   );
   gpc1_1 gpc3048 (
      {stage4_7[12]},
      {stage5_7[4]}
   );
   gpc1_1 gpc3049 (
      {stage4_7[13]},
      {stage5_7[5]}
   );
   gpc1_1 gpc3050 (
      {stage4_7[14]},
      {stage5_7[6]}
   );
   gpc1_1 gpc3051 (
      {stage4_8[6]},
      {stage5_8[5]}
   );
   gpc1_1 gpc3052 (
      {stage4_8[7]},
      {stage5_8[6]}
   );
   gpc1_1 gpc3053 (
      {stage4_9[0]},
      {stage5_9[3]}
   );
   gpc1_1 gpc3054 (
      {stage4_9[1]},
      {stage5_9[4]}
   );
   gpc1_1 gpc3055 (
      {stage4_9[2]},
      {stage5_9[5]}
   );
   gpc1_1 gpc3056 (
      {stage4_9[3]},
      {stage5_9[6]}
   );
   gpc1_1 gpc3057 (
      {stage4_9[4]},
      {stage5_9[7]}
   );
   gpc1_1 gpc3058 (
      {stage4_9[5]},
      {stage5_9[8]}
   );
   gpc1_1 gpc3059 (
      {stage4_9[6]},
      {stage5_9[9]}
   );
   gpc1_1 gpc3060 (
      {stage4_9[7]},
      {stage5_9[10]}
   );
   gpc1_1 gpc3061 (
      {stage4_9[8]},
      {stage5_9[11]}
   );
   gpc1_1 gpc3062 (
      {stage4_9[9]},
      {stage5_9[12]}
   );
   gpc1_1 gpc3063 (
      {stage4_10[11]},
      {stage5_10[2]}
   );
   gpc1_1 gpc3064 (
      {stage4_10[12]},
      {stage5_10[3]}
   );
   gpc1_1 gpc3065 (
      {stage4_10[13]},
      {stage5_10[4]}
   );
   gpc1_1 gpc3066 (
      {stage4_10[14]},
      {stage5_10[5]}
   );
   gpc1_1 gpc3067 (
      {stage4_11[7]},
      {stage5_11[3]}
   );
   gpc1_1 gpc3068 (
      {stage4_11[8]},
      {stage5_11[4]}
   );
   gpc1_1 gpc3069 (
      {stage4_11[9]},
      {stage5_11[5]}
   );
   gpc1_1 gpc3070 (
      {stage4_11[10]},
      {stage5_11[6]}
   );
   gpc1_1 gpc3071 (
      {stage4_13[18]},
      {stage5_13[5]}
   );
   gpc1_1 gpc3072 (
      {stage4_13[19]},
      {stage5_13[6]}
   );
   gpc1_1 gpc3073 (
      {stage4_13[20]},
      {stage5_13[7]}
   );
   gpc1_1 gpc3074 (
      {stage4_14[11]},
      {stage5_14[6]}
   );
   gpc1_1 gpc3075 (
      {stage4_15[13]},
      {stage5_15[5]}
   );
   gpc1_1 gpc3076 (
      {stage4_15[14]},
      {stage5_15[6]}
   );
   gpc1_1 gpc3077 (
      {stage4_15[15]},
      {stage5_15[7]}
   );
   gpc1_1 gpc3078 (
      {stage4_15[16]},
      {stage5_15[8]}
   );
   gpc1_1 gpc3079 (
      {stage4_17[6]},
      {stage5_17[6]}
   );
   gpc1_1 gpc3080 (
      {stage4_17[7]},
      {stage5_17[7]}
   );
   gpc1_1 gpc3081 (
      {stage4_18[13]},
      {stage5_18[5]}
   );
   gpc1_1 gpc3082 (
      {stage4_19[12]},
      {stage5_19[5]}
   );
   gpc1_1 gpc3083 (
      {stage4_19[13]},
      {stage5_19[6]}
   );
   gpc1_1 gpc3084 (
      {stage4_20[16]},
      {stage5_20[7]}
   );
   gpc1_1 gpc3085 (
      {stage4_20[17]},
      {stage5_20[8]}
   );
   gpc1_1 gpc3086 (
      {stage4_20[18]},
      {stage5_20[9]}
   );
   gpc1_1 gpc3087 (
      {stage4_22[23]},
      {stage5_22[6]}
   );
   gpc1_1 gpc3088 (
      {stage4_22[24]},
      {stage5_22[7]}
   );
   gpc1_1 gpc3089 (
      {stage4_30[6]},
      {stage5_30[9]}
   );
   gpc1_1 gpc3090 (
      {stage4_30[7]},
      {stage5_30[10]}
   );
   gpc1_1 gpc3091 (
      {stage4_30[8]},
      {stage5_30[11]}
   );
   gpc1_1 gpc3092 (
      {stage4_30[9]},
      {stage5_30[12]}
   );
   gpc1_1 gpc3093 (
      {stage4_32[8]},
      {stage5_32[4]}
   );
   gpc1_1 gpc3094 (
      {stage4_32[9]},
      {stage5_32[5]}
   );
   gpc1_1 gpc3095 (
      {stage4_33[8]},
      {stage5_33[5]}
   );
   gpc1_1 gpc3096 (
      {stage4_35[6]},
      {stage5_35[2]}
   );
   gpc1_1 gpc3097 (
      {stage4_35[7]},
      {stage5_35[3]}
   );
   gpc1_1 gpc3098 (
      {stage4_35[8]},
      {stage5_35[4]}
   );
   gpc1_1 gpc3099 (
      {stage4_35[9]},
      {stage5_35[5]}
   );
   gpc1_1 gpc3100 (
      {stage4_35[10]},
      {stage5_35[6]}
   );
   gpc1_1 gpc3101 (
      {stage4_35[11]},
      {stage5_35[7]}
   );
   gpc1_1 gpc3102 (
      {stage4_36[0]},
      {stage5_36[2]}
   );
   gpc1_1 gpc3103 (
      {stage4_36[1]},
      {stage5_36[3]}
   );
   gpc1_1 gpc3104 (
      {stage4_36[2]},
      {stage5_36[4]}
   );
   gpc1_1 gpc3105 (
      {stage4_36[3]},
      {stage5_36[5]}
   );
   gpc1_1 gpc3106 (
      {stage4_36[4]},
      {stage5_36[6]}
   );
   gpc1_1 gpc3107 (
      {stage4_36[5]},
      {stage5_36[7]}
   );
   gpc1_1 gpc3108 (
      {stage4_37[0]},
      {stage5_37[1]}
   );
   gpc1343_5 gpc3109 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3]},
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc606_5 gpc3110 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1]}
   );
   gpc606_5 gpc3111 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage6_9[0],stage6_8[1],stage6_7[1],stage6_6[1],stage6_5[2]}
   );
   gpc1163_5 gpc3112 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[2]}
   );
   gpc1163_5 gpc3113 (
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11]},
      {stage5_10[1]},
      {stage5_11[1]},
      {stage6_12[1],stage6_11[1],stage6_10[1],stage6_9[2],stage6_8[3]}
   );
   gpc615_5 gpc3114 (
      {stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_12[0]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[2],stage6_11[2]}
   );
   gpc1343_5 gpc3115 (
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1]}
   );
   gpc1343_5 gpc3116 (
      {stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[1]},
      {stage6_18[1],stage6_17[1],stage6_16[1],stage6_15[2],stage6_14[2]}
   );
   gpc606_5 gpc3117 (
      {stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[2],stage6_17[2]}
   );
   gpc615_5 gpc3118 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[3]}
   );
   gpc606_5 gpc3119 (
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage6_25[0],stage6_24[0],stage6_23[0],stage6_22[1],stage6_21[2]}
   );
   gpc615_5 gpc3120 (
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[6]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage6_26[0],stage6_25[1],stage6_24[1],stage6_23[1],stage6_22[2]}
   );
   gpc1163_5 gpc3121 (
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5]},
      {stage5_27[0]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1],stage6_25[2]}
   );
   gpc117_4 gpc3122 (
      {stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc606_5 gpc3123 (
      {stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5], 1'b0, 1'b0},
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5]},
      {stage6_32[0],stage6_31[0],stage6_30[1],stage6_29[2],stage6_28[2]}
   );
   gpc606_5 gpc3124 (
      {stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[1],stage6_31[1],stage6_30[2],stage6_29[3]}
   );
   gpc615_5 gpc3125 (
      {stage5_30[6], stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10]},
      {1'b0},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[1],stage6_32[2],stage6_31[2],stage6_30[3]}
   );
   gpc606_5 gpc3126 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[1],stage6_33[2]}
   );
   gpc615_5 gpc3127 (
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], 1'b0},
      {stage5_35[6]},
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5]},
      {stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1],stage6_34[2]}
   );
   gpc1_1 gpc3128 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc3129 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc3130 (
      {stage5_2[4]},
      {stage6_2[1]}
   );
   gpc1_1 gpc3131 (
      {stage5_4[7]},
      {stage6_4[2]}
   );
   gpc1_1 gpc3132 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc3133 (
      {stage5_6[6]},
      {stage6_6[2]}
   );
   gpc1_1 gpc3134 (
      {stage5_7[6]},
      {stage6_7[2]}
   );
   gpc1_1 gpc3135 (
      {stage5_8[6]},
      {stage6_8[4]}
   );
   gpc1_1 gpc3136 (
      {stage5_9[12]},
      {stage6_9[3]}
   );
   gpc1_1 gpc3137 (
      {stage5_10[2]},
      {stage6_10[2]}
   );
   gpc1_1 gpc3138 (
      {stage5_10[3]},
      {stage6_10[3]}
   );
   gpc1_1 gpc3139 (
      {stage5_10[4]},
      {stage6_10[4]}
   );
   gpc1_1 gpc3140 (
      {stage5_10[5]},
      {stage6_10[5]}
   );
   gpc1_1 gpc3141 (
      {stage5_12[1]},
      {stage6_12[3]}
   );
   gpc1_1 gpc3142 (
      {stage5_12[2]},
      {stage6_12[4]}
   );
   gpc1_1 gpc3143 (
      {stage5_12[3]},
      {stage6_12[5]}
   );
   gpc1_1 gpc3144 (
      {stage5_13[6]},
      {stage6_13[1]}
   );
   gpc1_1 gpc3145 (
      {stage5_13[7]},
      {stage6_13[2]}
   );
   gpc1_1 gpc3146 (
      {stage5_14[6]},
      {stage6_14[3]}
   );
   gpc1_1 gpc3147 (
      {stage5_15[8]},
      {stage6_15[3]}
   );
   gpc1_1 gpc3148 (
      {stage5_18[5]},
      {stage6_18[4]}
   );
   gpc1_1 gpc3149 (
      {stage5_20[6]},
      {stage6_20[2]}
   );
   gpc1_1 gpc3150 (
      {stage5_20[7]},
      {stage6_20[3]}
   );
   gpc1_1 gpc3151 (
      {stage5_20[8]},
      {stage6_20[4]}
   );
   gpc1_1 gpc3152 (
      {stage5_20[9]},
      {stage6_20[5]}
   );
   gpc1_1 gpc3153 (
      {stage5_22[5]},
      {stage6_22[3]}
   );
   gpc1_1 gpc3154 (
      {stage5_22[6]},
      {stage6_22[4]}
   );
   gpc1_1 gpc3155 (
      {stage5_22[7]},
      {stage6_22[5]}
   );
   gpc1_1 gpc3156 (
      {stage5_30[11]},
      {stage6_30[4]}
   );
   gpc1_1 gpc3157 (
      {stage5_30[12]},
      {stage6_30[5]}
   );
   gpc1_1 gpc3158 (
      {stage5_35[7]},
      {stage6_35[2]}
   );
   gpc1_1 gpc3159 (
      {stage5_36[6]},
      {stage6_36[2]}
   );
   gpc1_1 gpc3160 (
      {stage5_36[7]},
      {stage6_36[3]}
   );
   gpc1_1 gpc3161 (
      {stage5_37[0]},
      {stage6_37[2]}
   );
   gpc1_1 gpc3162 (
      {stage5_37[1]},
      {stage6_37[3]}
   );
   gpc223_4 gpc3163 (
      {stage6_4[0], stage6_4[1], stage6_4[2]},
      {stage6_5[0], stage6_5[1]},
      {stage6_6[0], stage6_6[1]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0]}
   );
   gpc23_3 gpc3164 (
      {stage6_7[0], stage6_7[1], stage6_7[2]},
      {stage6_8[0], stage6_8[1]},
      {stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc1343_5 gpc3165 (
      {stage6_8[2], stage6_8[3], stage6_8[4]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3]},
      {stage6_10[0], stage6_10[1], stage6_10[2]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[0],stage7_9[1],stage7_8[1]}
   );
   gpc623_5 gpc3166 (
      {stage6_10[3], stage6_10[4], stage6_10[5]},
      {stage6_11[1], stage6_11[2]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1],stage7_10[1]}
   );
   gpc1343_5 gpc3167 (
      {stage6_13[0], stage6_13[1], stage6_13[2]},
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1],stage7_13[1]}
   );
   gpc3_2 gpc3168 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage7_18[0],stage7_17[1]}
   );
   gpc1415_5 gpc3169 (
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4]},
      {stage6_19[0]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1]}
   );
   gpc623_5 gpc3170 (
      {stage6_20[4], stage6_20[5], 1'b0},
      {stage6_21[1], stage6_21[2]},
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage7_24[0],stage7_23[0],stage7_22[1],stage7_21[1],stage7_20[1]}
   );
   gpc1343_5 gpc3171 (
      {stage6_23[0], stage6_23[1], 1'b0},
      {stage6_24[0], stage6_24[1], 1'b0, 1'b0},
      {stage6_25[0], stage6_25[1], stage6_25[2]},
      {stage6_26[0]},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[1],stage7_23[1]}
   );
   gpc223_4 gpc3172 (
      {stage6_27[0], stage6_27[1], 1'b0},
      {stage6_28[0], stage6_28[1]},
      {stage6_29[0], stage6_29[1]},
      {stage7_30[0],stage7_29[0],stage7_28[0],stage7_27[1]}
   );
   gpc623_5 gpc3173 (
      {stage6_28[2], 1'b0, 1'b0},
      {stage6_29[2], stage6_29[3]},
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage7_32[0],stage7_31[0],stage7_30[1],stage7_29[1],stage7_28[1]}
   );
   gpc1163_5 gpc3174 (
      {stage6_31[0], stage6_31[1], stage6_31[2]},
      {stage6_32[0], stage6_32[1], stage6_32[2], 1'b0, 1'b0, 1'b0},
      {stage6_33[0]},
      {stage6_34[0]},
      {stage7_35[0],stage7_34[0],stage7_33[0],stage7_32[1],stage7_31[1]}
   );
   gpc1343_5 gpc3175 (
      {stage6_33[1], stage6_33[2], 1'b0},
      {stage6_34[1], stage6_34[2], 1'b0, 1'b0},
      {stage6_35[0], stage6_35[1], stage6_35[2]},
      {stage6_36[0]},
      {stage7_37[0],stage7_36[0],stage7_35[1],stage7_34[1],stage7_33[1]}
   );
   gpc1163_5 gpc3176 (
      {stage6_36[1], stage6_36[2], stage6_36[3]},
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], 1'b0, 1'b0},
      {stage6_38[0]},
      {1'b0},
      {stage7_39[0],stage7_38[0],stage7_37[1],stage7_36[1]}
   );
   gpc1_1 gpc3177 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc3178 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc3179 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc3180 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc3181 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc3182 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc3183 (
      {stage6_4[3]},
      {stage7_4[1]}
   );
   gpc1_1 gpc3184 (
      {stage6_5[2]},
      {stage7_5[1]}
   );
   gpc1_1 gpc3185 (
      {stage6_6[2]},
      {stage7_6[1]}
   );
   gpc1_1 gpc3186 (
      {stage6_15[3]},
      {stage7_15[1]}
   );
   gpc1_1 gpc3187 (
      {stage6_16[1]},
      {stage7_16[1]}
   );
   gpc1_1 gpc3188 (
      {stage6_19[1]},
      {stage7_19[1]}
   );
   gpc1_1 gpc3189 (
      {stage6_26[1]},
      {stage7_26[1]}
   );
endmodule
module rowadder2_1_40(input [39:0] src0, input [39:0] src1, output [40:0] dst0);
    wire [39:0] gene;
    wire [39:0] prop;
    wire [39:0] out;
    wire [39:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_25_gene (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(gene[25])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_25_prop (
        .I0(src0[25]),
        .I1(src1[25]),
        .O(prop[25])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_26_gene (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(gene[26])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_26_prop (
        .I0(src0[26]),
        .I1(src1[26]),
        .O(prop[26])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_27_gene (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(gene[27])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_27_prop (
        .I0(src0[27]),
        .I1(src1[27]),
        .O(prop[27])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_28_gene (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(gene[28])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_28_prop (
        .I0(src0[28]),
        .I1(src1[28]),
        .O(prop[28])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_29_gene (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(gene[29])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_29_prop (
        .I0(src0[29]),
        .I1(src1[29]),
        .O(prop[29])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_30_gene (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(gene[30])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_30_prop (
        .I0(src0[30]),
        .I1(src1[30]),
        .O(prop[30])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_31_gene (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(gene[31])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_31_prop (
        .I0(src0[31]),
        .I1(src1[31]),
        .O(prop[31])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_32_gene (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(gene[32])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_32_prop (
        .I0(src0[32]),
        .I1(src1[32]),
        .O(prop[32])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_33_gene (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(gene[33])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_33_prop (
        .I0(src0[33]),
        .I1(src1[33]),
        .O(prop[33])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_34_gene (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(gene[34])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_34_prop (
        .I0(src0[34]),
        .I1(src1[34]),
        .O(prop[34])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_35_gene (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(gene[35])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_35_prop (
        .I0(src0[35]),
        .I1(src1[35]),
        .O(prop[35])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_36_gene (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(gene[36])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_36_prop (
        .I0(src0[36]),
        .I1(src1[36]),
        .O(prop[36])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_37_gene (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(gene[37])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_37_prop (
        .I0(src0[37]),
        .I1(src1[37]),
        .O(prop[37])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_38_gene (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(gene[38])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_38_prop (
        .I0(src0[38]),
        .I1(src1[38]),
        .O(prop[38])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_39_gene (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(gene[39])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_39_prop (
        .I0(src0[39]),
        .I1(src1[39]),
        .O(prop[39])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_31_28 (
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CI(carryout[27]),
        .CYINIT(1'h0),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_35_32 (
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CI(carryout[31]),
        .CYINIT(1'h0),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_39_36 (
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CI(carryout[35]),
        .CYINIT(1'h0),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    assign dst0 = {carryout[39], out[39:0]};
endmodule


module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor2_1_256_32 compressor2_1_256_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9b3efca63c51239e96acb4cc372b3030f8ef75adc0c2cd4f1d9456a0795c079cae4e548cc6fbd8bec4b914689bc86fce47a3978c0d4070c3b33657207bdcf58f2049c6fbb90e2a230a04d9f74031c0ab85293e0dac4b87de8f6787d2c280cb0dac1cf11daadc9a1ccb6f5643996612d8a4cdb14ec76b0ac011824df14b4d15bd5918930cd6555dd590a964aef7b4168b07c72e57852cffc063c629114723e9746516f43395f1e5aa6067e4ff93462a5f64dce94a320ed26cfe0cd62bce081da246b96051da647c2895c8a9042b332b7cf14cae8cecdc47df806388f5a8764785a8a01ee0e7d01047aa87f8d0d62421f7fc0a21173a777d5f417da79a294934df19f2e3b134db0bb343badb7d4e766de02d90a4bc37003522f769891d4802e16854206e2a503cee76b28b6092fe9e8e65f9db16048130faeea28e4da879f9d69347717ec7998377d1ad3742901af6e783f439f0eafe4d9772dadd73bb44e106517c9239a5c9a7de92af20a7929fcfcf6aaa0fd597f3284938d663e0149054948c47e8e439746ed1a9589b982c783a1e419a249134f991c51450ede8548c23bf5b2397525478eb7351a2045db8619f687ceb82f0b24539465c1279fb83a4037915692fb3cfc49ca111c45bd81ad972dca4438f00f1252f7cf324b3ea4bfdcced54465448296df4aa825024140547555c6cd75aac5e2774556c48c723fcfad8ef451ea28305c7a4d99e6dab90d74d9693bb1768c97490f149654f3315d8647f5d2ac38bbbd670f6b9ff43c4921b2f374f98eb75c85a47a27b01ccdece969f48676fed8fdbd92054cb8abb9be4544099dac3bbfafe6e38924aecd1a006163782230b4ad827e8b605fe1828485dda67b27f7f0fa3808d76e5a2620bf48f8aeda9c2b3bc110affeea66969ab65cdef03236547ce84889c9d9e32d18c4abc605c36368bc811d9023fec6ff7de37efc0712b69a849e9a97f0dd58614e8e49c2237e67c3b5211e3b51f84ff15e5bb808a022d486e39914bb4ee69fa545d1c3a6f2813421582a9cccdb3839ac076017cf1c57cb68880ba10d22a9744d9ba88f42ec2c0dba0e0a6b1165e35852d1865037bebb2e392c0300699d6783c9bbe798c62a3e56dabd65694764131252a449bac58f970ecf6fb8cc8dbc3ac196d2cc1f01394230da22ced11a80070999bfd82ad282de5f82c18944a9c6a82b9948000c02c103137805988d1a8eb310a3e961781e78abd65277a8edb0433a53eebba0b4d38ee74da21a899847b29fa5dd68f7366f2a65edd2159d37c6eabb6bc6a2681c32076d19108b8c298da35052a8d752d72f6eacc2bddc10ef36e805c0d558ac35ca3e603d8f816f002ba3627a1380b6d9a9f05c86c1f4d9c58f30c85305497ce9d4272468c53f0cb3185112fb6b357de3b7ad44716fd51b24d08eb09eda12296ba8907a0cf2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfe88152dee5c1606a9720890c53406ace8d5eeacf16499e3c3b536922d3375dbd7508c9b2d8eddd354b536e38230dd9068328ec74e2cf4156c5c591570f8e05d18bc19a09e3742fe4b917d1b60322f012229060cce062a5dba25a66d170430c9422eaa2fc6876119039bb0f2b6240e5b4a684e05c5278615370eb96b3d6b4135d5c893f78e0f99b33d29ace7f398d49f3492472f826c64774870c31f131ac869efe3b8e3d2b74f337bb9dcc1993915cf72193f26854097d97f26c87b6186bc452567a95f434917748841ae5d7c949e9f3bddefebb648494484ca661a3fec744da32b879e4c1d6a818ab094d88d48add03d6bc4e3740d84d43e246f89d5eee6ba61f3748b31a74e8611afa1c5f0b85195d3eb5ca6c18dfa49900b507e34ae7c89893db031c0f6ef847442bdff2eae99d0e7aaa8212771fe7006ce22a7d0f0b06843622b503b43052a994ce7c366f846c5886d05ccbc7938708aeada527bffb57cfa208921fd7f04bf309cb0b2c4f3b6a4812eb538418e73ff2e50f19206813f6d04f8b7b7799b85b9f2268a8dfa316f95a8d2c93c333cc7ca4cf51ce8af2de4290ce9a878340946712320565857dad4bbf055b97dd0262d54243435fab8b4a5f9048054950ea508d98f6dec4259fbf4696779bee0bb6125a910d8f02e8895d0717e8aecad510a9dd007b70c56b31c24b7493b8eba8b4add2bd66e32ee518893cf4657948b7a88178bce0f573a97fd5038679f3c71e98a41c39ea1996fdb4b759c222cb2af2bd09a514b9986c5e1abbf1afaaae33393be4c51ce9674b2bf596a7322e42591add9e5acc8702cca68885d3c347dc688a39d57d9d812f1307ea9fc5fe626446f8586e5ed8a460f2cdb45e90e4341f999bee03b36e5b8d74d2eba92370a510949d8158a1968966d416e149de6134524c5542b8acc5c242c897b87b8132a41f8033423f8d652d8dba29a2893ace57594482965aef8812115e8b7609b334a51353a70d6affbac4bc339077c6d9bff0ccaefb039167e5ecc23f204510e09db575ed86669a0248a14e612843d401dff0412d2d274a210c14e469733fa6052ac84e7d8bd5baa1304fdccd2ba4f50f58c58b324e1d00736c32f46a6d2a1ed86719cdffeb353501486773c2155eaeeaa7a979521db52372faef9eac90f12c2ff7c68428dc567b22a144cd956cc6163862e10a0331163bfffd48808475c2147c72de983d68c71293c269fb174e25d5daf48c645ef7ee6ffbe2667d69c687b652169f8691d474477661f994a49b4fa7f9c0cabe1c16d1cfb9f35815705f4e895cd9ed5e372c6ad8fa52fe3dfe1a07cccbca2db0da3611f08cf1a25dfa6336b29d4187c3a9d29df01cf5997458c842cea1ab68b491de5994b5f873c618dea8d05d3a1ad96805e65e6edbf71956e3bceb7a84df1cd99c106904fd78ae34488897fc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc3109cb2a48acf770b6228810785bca168f4ce7c1bcd61f22b5f2cf719dd8eaaea50289240d3aa509009b42aef8511ed10c2a89dc14be7037800361e3be17dad18a5318d9b5bcc5db0e0f19db5e4e77191a844f199b1c4ac72bb18fd4978b432a7198357365bf51ccaf6cf72be6f9a19355affbeddd84a2908096aae3e280fd17686c71099c927030adb2e78f7f891d0db55c1ec3738ba808498b11262f78245bbc3ca1369a5e3ca5b8e58d4669a645ed74ada5c9dfc80f8e19910608dc82bba11ade0b96320c1f78c7c507c616acfbb38414add15545b0f6e4e5230caf252da023e028989ef1290a31dd052e6c3efa6dc7667fa8ddbb07f712aadf7ad57f8eec4f328615d9688d11c8905482bdf0c8a05b5911452547dc85c51fc749ec45f8e77cc4ebbe0228054f19e9f8f117f7d25ea4f3e315415a89094034664ac36dc9c7a02fdba65dbd48af58bedf6a7e46470c45f42263601794e929a6f8470207b846c081dfdb1610e24bd52c78dc27174333af5ad8eaddbaec1080b2f20505d21e40e0ad36f312d21e80308d44bd19577c6377874a181cf08f57ee2012cf3151c29e9a6861cf59fd60aee1487c11a6a371a5bbd444b5c1359e1de831aa567dd391e4fde4be6ea866dce835a1adfac02de00e9b78151a500bc9df0cadc405f409dbd328efab516b14774c4ce9a575c3f1766ba7ce336adbf3a75b5401fa7d32a728a444ae1378c013c99ea67752d769241eb31f70cf9f6b02f6c909915dbf2e037017ce8701910b39579c6aecc220fa4d1af06a80d68dcf8aaec081abf45e17093d77e169624841993071765010dd813f08c4ab591f2b8202592be79afcf65db0e1b06f4328783d90069713fb56e9dc2c2a07f1936a803992126f427f5861009f155d69e6cb236731cab6cdc73e42a043e25bc0f60e07f6789631bc58090e808c3015429abc5605e3ffd86813fc9c44710b74e186f15d304dceb77077d8e3c5819f6bac36fbe7f2fd24a117648f8fed7c6d78f3db4b5f2ad251376dd55c7e9fc2106340ad6836bd67af3c809a4393dd44e8120f4d742274ac02e786bff4d2141fd5d0dbc8c79c13a338e49da0edaaa62730b01441771d1ec6604660f6090229107e2e1a2d644185c9c605f050da30a7b630343d89a9e334120545c64936c12c808b33784c28f9bd8ae0737d544451fbb5a1f337d2cbf0381def18be569c167a7713aaea00ca0b4a2049304257715a32f769ecdb5a77c73608bc14d95c30eb47bfc9543ac5696b371715fd66b99f953d85789bd068693b7715f8649891ae0cfdfa22d535bc65129f7b0683bde0aa36ef40a2edaf4d1e36d86cb9a0117bede3aea72616d50cd036a94d8278e49a94a5d2902f66306eea5cb470e04e93cbb51e61510e56774a6cab43a89fb281836f4f7f080c813477a513b447c44c292d8f528f1dab5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3087da866f84b2046aa1c19c4e64aec816867b713eba29b2d5474c37447ee6eef210cf4507423de01c2dd8d4a8d6afb154f24d88ae5012b395cb26c2d6cf6d6f0c0b77ea7674d737a804d7d491c143f2e4af98ea5e81c93e125e1059ac928f895d67da70c6f38e6c6eb8f477339f48544c9393789be019e399691594c5de28e78d5210d2ed9c15257dfef5e535b534f85f6a375ece0d54fcab495edbeaba20c1860796ff3331085a098b0275d2bba48c40ddae26536d3c10c858bf9da446923768e9ec585a52834d0ae4bfe7b6be1fc1a909205688aae6f421f40c549e6b9f535d3854e2ae4fe3d123d2c0acaa3b7f11094a30d8b6730f4dd5fbfcdc2fdb6c046bfe3968b5c7a6c67b3a7f0bbd696243de2a8fd942a783cd7e6edc5aa81ae033fc0325461cec50a319e2de718343c75840655c090b976da66aef0a6032f4a7cb99d0ca589064f99a8380ae323097fd0a8e5ad9d7f197e3b519c2a2c52530a87724b7be992b428bf97bca3e4b950193c545befbfb7344f9fda717ec39d4460e67a253a38a56ce8eb58d476a3c1f170593c31666dc2256fa818491ffa370fa693090ec13c01c2019804b26afcc38658b93c131de381320eeb99fafef04fd55acc64311919328e31c3ae23a4ca960bd2d9092d2844425085490a0952f0b32ecc772714f65af05b2d1b1c3c6da79817f830258a930c6c608ca3d79f361491cd5dd5c19a8afeea9e4ec8dab9355d5fb1cfdc9732c3eca336edd83db968b58a1277cbb7f43e381c6ac308af06a784f6518455f681b47f049ac16129f5082e1916d8506ef3850407b997c7c02916de9962ca4a8a6ff9cb9738df502ac363921b9da8ed336c9b3d4202ede545b8fa2e8bc7b62213337b13cdbedc43b445f2211e7f24ffb831fb541f2d1c8bb7748aca96c60206418a7c8e0e7ef2872b90aa413b0f25cfaa96129b2258de90a9debd97d2b3c76c2b7fd2c7880c90e65c7052e2c3d95722d66a3394b85603edd1f55314bdb5832323d9d9d13cae381f5361e6ab624d7b0d0a2b0aa97e499663a6b42534eaa8fda3d88cc14ce84bc01938cf1689380b4c2949a9f0b0a8247b7cb2a0b59b5abfe761c5de474271504d55a01aae51ef3e432828efdb4309f9cd57c08a2b38d460e7e2c0af09ddea2de664e0eb34293da78eca0e8ec5cd4940c1500301dc496ea2abd343122b2d78baf6ed98a960d64b1fd9b4e28d7bfe2b72648cc259ec8f2f2fbd4f6d1b675625c71a36d39f0fe3b313af2a6e6f1ada9abb036ae105494397103b309d5664a4e8cecc8e56e19c14d034572f00c128694b55f80fa7638a129ec21e4787a8589d48d5210a1d4e57db389a95a97a2f20ecffcd4f1f42fc5a057bd30781826debde7f5c1ca333a903b6039f1c369b3324c4e164e2f37183780a2388f63d3e47f9d25565bdf21d235f165a3ed3cfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4050cf953a67326a11b0c514677cd51b6d0e27167ca48958916c0e85312100fe22b2b9d0db51cc5d0f270aa42f4e5b3cdde7a83ca82395aaf98d6cd00b31de7e00a39ad11bcd494fd469e05424e61b85e91141e46ef2fce6dd91d091af52b752abaccda4480b332cc418a65d6340b86fb8391658636cad3b52ca71bae55f585a02c425dba8ea1e844be83d1c1d2ec44796220dbb726c551be9b1c9977d54a821860efe6b0d3623617f4d77adcfd72ba6abe746fdc2142a7981eb9fc1ab51c8a331deb93eee611f90674e5c47c43cc8033b81722a0e9b55cd76f215d44723f2eba9074c0fd019f5dfbec785e3ee057de0c8149ec97cd81e090c9c0c25799aa30f0b75dd71439ca61dcd75177025fe11f99909d5746181462e85fa2699d909387111d1016decefbaf154dd05206995fd873deede4ad173a7b8a33fe33dd0001c34f4a6f00a11b501d687fdc27c84b8924d8020a3dc2a968639a2e82ec410a9ea8dd264ebbb74ebd6dc3384ed1e0ca7251c6a8561cc7f26441c3d86143bab842f2a41aba0bdfdb8fa32c312808ea1d06d3f3bf095d6cfbe22b23030ada792dbdd7940df767ea09fe26348f4d2683479d3f1860139231577baa3df6e61f8e843e06ae234d9cd1d5fa133e2d909bb27f46e2c10177a92df01f3b7780a7f5da93c167b1904db775da7bd80c49f7abc55dfa3adf3e618af409313c0a0ceef65293732e013c3b84fdca7ff67e110501824dddd811280083df564158073e2e19c7bcf501afb5847e601da70df6cd818673e00a639bbc2c72dfcca66ffa36d93431b9870e798c88d5bd97d627c293acc8eab7a22a0b10203b54b316f2071a9b87c4612b44274d40e5587306596fb2cd172ceacec11b2924e9794bc5ae2d7912dccb1050625f5856d09ee89328be68baad8e4ebf3c91c213404198b0481bd49462383c08a025f2c3b61f3137804ef985a87e4c6739f68e3c1d14f49e9084faece1acf2111dd4828ecf282fe192e766bbe5a037715c64762b758ecf6a2ea0bc7d92671d0bbb8b42925d075ec114c09151145b78290a4ec2ec3e2657715b7251865b9f4fe1d40339132008b1566f236798eeeba5c6c296d51d214da1ab78eadbe7d265ca4bef33ea662bd29343d3a7f2fecf32ec968472121f904de3fe15967be780ff4243dcd79a5b97f332bd2287110e477ef5f7c19a6f1acb49f41cf3679a627eb4ecb866c028e00a4a2f85db45aea1c745cea4a86bf12ddaa947724772981de52713e3e9a6ba9a18ec40236349057c519c260ef2eddb5f93af524e75d0ee8bd402e76601f7d1d8664f034880a866cdbd35708d9e18aed580b8332c69968f6da733862f52743b302b5637a2699a33934fd6d87a2f4f4dbf42ee52898ee68276be691705f09c487fda12387a7f1edc4f713e8e847561548851153ee482a80267bb01eede8c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7ca0356f242e9e8f0f4ed004019011dcf0ffbe445f64d344a9acc3ca1cfe7d3643b3b1db08a2e5d4177e37d01d43cadf6c727f9eb9a8fbfbc284efb9799f67a219d3396117c84ce153b91fa945dcdb59c66940181f70dfd51b08138aad0d3f0a145b5e94a95d8471fa285bc861522caa8ff4b1689b63e2622b35d966e44bef9c62946c12f2593da30007914b3261ab39fa4404fc29059798aa7d0ac54b083f5ae2beaaca95aadd13f0373e1d5a5331d6316c77cd3002503f4135111bee344e3536f0812b8fd97cdfda5352346dc41a1bb9e2e7fb40acee5bab73d4aa5a318c7eec042e7a9e60e02b72edf1f0e8ce3ee87fd453350387d2cfbc39d814b42ac668751bf0e73f79fb3e52df7e1cd081f05c5ce1678199116bc20c3ed3dc6b3884759d20ce6a154b4790f833281c5eb55e2d42c77815333a5115b4c48f45987d9ad31b4bdd448b5c27a08c32fc3f775508a8970f7d73cd7a054fc6da7a989b1f3cb3f9165ff9789adbfc03ba9007e3c3010327715a8a21b3d577369066cafb2c2d666e8be32f4acf4d9d927ff301e179253f30d79f490b1cd29c90730046caeac0f21ac5a325049f727e8f74af3aab7cce8958531292f92a30892d27917de6ac1728f1154f1d4415f8ad1778350b7b32d52713cc3535cde50ec63d1dbd17d9ea890dbd4dde1c469cbde126a07b076a9fbf179b730cc2404fc4b643e3e2a54a6ad674483f921d206b42b8b2c86ddb18693fab69320ecd023c51ee94c5f79f349f002d9facbcd149c3bfe872771a14ddfce38d7c9ab5d7970da9fdd4b2f123e94dd9c767d471c00b5a9c9907faf0479fc8663c125c45819ac484155055a4147b4833b7f08ff94b3471eb9d2ee0329f17fdfb19cf189e2663bd02706ffbe0587c3b929389e32dab399bfcb8c4fb99a44dbbf04b416e9b053e30a9508a85cabef6a5c80d402a16c01be544e6689721c4829f23510aef1a5ab7f0171fc8b7bc3df3f8f5cc579c04f670344f0eb9956255612d2cf8c3bf73f5da56d9c7c417cbdde975819646a0336b1bf4c04ecf9c391c29f5a3b65c3ae027398f6c2a6a55baa573f74c858efe34c57e1361502819aefaedfeee1979c53ff116122fa71c92732883ed98a2342b43f4c2858f33cc8207d1926db9f2eaa4e87624427a06ab48f2a4e9003a765c9a5e525819ba534a7476ed0f296024846be92cd951adb866ef6bbe9c5e7ab6ebf356fed4ec1a0fad25186c9314ccb996128f80d8b7bd614e6fc7130fa99771e27d5a8ac9e7de0b20359ee1600f4367a75241d82143fb3dc408a8f1d413edf5c5e063cda82acecb82ee1d3459c35ee43fb204c5a27778205e0aebaf137f10ac0cc2c3ac9983f0da1c924870cce53e12cbc1f2316643775c11d209b9233c724c76b175d25622a1124022790008c682df707128add3565a1c295f7679311a876f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hec2ec72bbfc7a2ff7cc210d8c129c6106f19601cb234ca9dfa3d41606c2aa2dd20dbc5dfe38867ac472288d196a7580bad27f2da4ab1e4f533ad457ed72e02f0982f2c55d5569507df8e6467a487fb106534f034d7c5c68d12ca022c6e0d7157c0bc4d04a4f797b69baeef585fabc9990f76a790e6d0230e6c5979ba7a860a3c6bd480b4869b09158aec09061ca5076b6a736a24129c6ea066fff11090cf90580e0c1670d5b081f2a9cd160d2181f8d6584ad558186653a7741bc7e248fb1cf51e43ac7873b0edda7fba30df599c125351d53614592f8d277f00e3a9abba473911f8232a55061515ab78e095ed34c3322a8669fcb12e8a9809b5852e0a72eb918136698e45cf3b12d8d0755dce31762d390c2ac329580d083f3f6caf78f9e1374ee0a239a7d8b1f28db847fe26b89f1ffdfab9e6eeed76ccb3fb1873fba36306d2a7487d2b3b6ba201a69880b2882fa2c3561884f5ca71e5099c18eef3b5e562b10e3fb77c5fde7e0cdcaa9009e2d3b0a09f3e474a57a02cc3e9dea97eb82351ad35d961d5c49a6f71696913bde80ff13ee290faa032584432e10abde6ad4f5916b13d63889e56b7ef96a2b1359d07dea47425fbc1d7fbbabbaf9d80fb9540322e2fae187be88cbcd1bb5e077d855928c742c2cd776e49f7cc43ff24c73cce3f57d0f9af3d01bedd6a617bc1f95b91fbf8508866b0442e500943375a05223559384cead6bb08a2194e02a25b193a8d6225fc20aec6c5835d35f038ca9bfb3656d36ab03eaf71d52b5504f0b110fc25ab375ceb522338ccc3ccec9883b96a9eef062c7a35fe6eefe6f869167a2303473946c4889f97fab0762264198f09540f39022ff8bf32b6d7d6c832024e74c7c863a6999a44dab2d097d7dc8cbc14a55858d2410951f40d322c733866a79cfeb577ca5edfb5de1afbc442bc1ebdef501aeb12d94843b1f9169966006bcfb4d1c78cba52ed541d0d471d97dec52ea07adff61b00c0ddeec75e2f18cf5db48feebdc882fa3886dfcd1e82387ed9f63b2f9d91d2f250c6ad705e9db0f5e9406ccb4f8d3ac52abfdb8d41ac8844789b06ff11b992eb701df22517c846997a64f0520ca6e39329cf5e1fc2527d736543373799811b63587c915acc32ba89be14e21dcacf15b75ab8a6b09e2d02a25632faf3f7f5b9685d30a1da0a84ede8a1f8d744581870ef35bd252bb0c415ffda6530c86128da13229693d317ea6eae2db55e6cbedc7ce83227f89b5d1b4600200b71f6242a3dfe1e71c1347ac8b4ac692771c622b9156c9d06ab69e7facdb7289b2611ee8a013a3e3d13e9936944b5c1992d4e15a5fe2aadec24b767062c60ffddf69d76de5498d3e807e923fe4450b6a0d10e08463102607ce77a31ad057417e51e74b67c23a1a36077d8cbf0483472d98035d89f7ad460e958bcccd04b8c18c4ff9efc2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h234d9118d48f54feb4ed51a5a55e2c4dba1cb1efedd8a15533c25fcc519b487e09cf16554c39bfd4caf10a40d08f69287c8a1ec3af7424122e0e002225d0827e46a502fcf432d13e82abcbf8b6a14da2f81733a5966c61c7661d78db75417051e9e9c92221938f4ef30af5d3d7b2832683a0773670e58b6db20d3422f7be43dbc6881ad39b69e377c5d02303a09c8340abf1f2455e0ffeebeb21d85fd83f52ad97fdc65c54362f44d5e19f75ff70eb2cbda31f5a81dd64944b792fedfe6deaa0775509be6cd3ac78b97d444aec2589e633980862c35de29166ef04cfefee3996d8cb31e55922841c23a114a07843cf00b1f6251970c6d0ccecfd175bf26ba7a1bfb3cf79d42597728221edaf0e6c1b8cd7f317a21d69ed7ecccec8567868cb28fbd3ca546c70a7afb204739fb64a8e435aa6628506327f039995c8bcb2128d49cb07ec766e93fb717df300b151838465d2b44233a9066db4a71d4e6860485ef55a1c74080b64e5e9b5f8a2fdbf0adb4e3125cf11c7acc30eabb58c002a9328ad15a9c0dcc3795204a6c4afb026fe4bd55606ab1d9d0e801f340aa2b0f81c12a2956bab93dffcb445e783a09f2c64cc20df14138a5cae4d82a600370d8abb6fe2fbd641865ab072791325611bf7bf7ad7e33dc53991721a8413dd9b3bdbba5f598ba1ac13c7397f41d7cea7dcf86fd3a91fe30090b084e6d643d5e7e49f0fe31a7b94179c7800978466656587c9496cb9e3eed740e4ce58abc414b7b1eb065bbd81cbde5e3b7ef97f89b1934fb7522b262e2843ef9717e685ddcd3f8f087978b456f39bb604a622686bca9c695bbb1b9f3740e5079e2527f2513d1176f0623c108ceabf9eba6b33703e0b5029c926f8057ef842a65e61f83eab2af6c801722b8064dbba2ca7fa8c5acb1fe5d3202e820c7e1105b1cbc6b759d5ed45fc0ce49159ca500f2523f1b06553d8a8d74339bbee89b491ddb1af424d49600bc74d32e4ce0001b123bf7eaefbf70e05f8341e5248dc5311994265f02fe8cc5a22ff11aa661a94c7d867d48342d974d45bc300a437d3ad289b8ed63eb86dd6a3bc977b3c992b7efdb45630841b4181286979bb51b9de8b7a3b34213eaaa158fef307ccb6688b237486fa266240e8141b7eab4b9b75f5177ea8218105d8bb83bbd168dbbc4c8190b8ca1adc7813279aaed3ceb5e2a495f6994d36935c8ee667e0769805acfe3b26aae1452882b6b306746604c0e0ab4739a21cd6bab449aa7ef1307d5df0d643ce332af9a6a1bfd24bbccaadadc4913d86287ccdccd8446a9c475a50ed0ba1f5a82d84de3cfa8f92091740992fd4b9a81bf40b15e50f14a7350a93f7d5df3e2c9ab8c6b373cb58a36bb8226a94e3bd10bef37a36748690e1e9a227a6e2391fb2ff5b567f113f27998a589b26c9d6e2e477bf5c3fa22f1af40773bceb60c2bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heec35e1fd7b280b2cf35e17a90fe5e0fe7d944543cd89d02dcb25c2e10946b9d2801acae52664d956f8fe69abfde1feb59950330b2913020cf78eebe63ac1dcb56920acd00c3531ecf94afb90f78ff54c62edc5c222c4259bcf868cbd3d27e2529c5d5eecab9e4c6ca7237e9619a2ea11b6edb5e0fef9a8ec20edc82aea7ed3fc8c7d8a052a1fd2754b30a1787a9eb968458275438a5de014e67294a1a38af43209c1a1f0a67c7d0032b5e9d8843098c08b318f08301a36bafad53deafb1b3e6c88153e696aabc8c084bdd4adc66bde5394881599edf4fc285a95e5fa846932afd6a55a3483d72058d5d09d6e2b614c3699286766d68b8c03e7928fafec0ebfd5303b31805781b5ccc44e85c3a3574e2a6af1c73a4aba18bfa6b6ba905c53b24f686aa1d23483adfcad09fabd3ef8bec55669783ca3278496e5a7d2b1367f55b9e6d52a041fa7a1d1bb95ea02646ad0dbbefd66f2fc8ccfe6e1e2889b7a48aa1273baa2cf4aaa1bca4c4fb73d24bab74a5e3682e05edaad21e850e10ccd6beadab71fc7b3446cf823cbf6cdcdc1a695e1ed7d129b55140eea543bb54c463ada1d84ad44bdf433f0cae942d84eff7cbfbd32ed354cf888ca068dd34aad66f73c9c4ac27718de3eb7844079b3d7da7c4d2f923a8ac2c076ee09bdabe54207a4309c176114ea32e2c3c9b54578a82eff1a73a9af20b315b3e4c716e3e5f36853fc8ab5533019c40db11964642f1429430579360ce21f6292ff5717fadd4e57554b031777892a8eaca5fcfb9c258f564d234a30a8985d713a8abb3828b5ae6c5774a08b3c208d2225f634ced2a60ffef3a982cb13b8a7d57dedd11b9cd1e0dd43fa47809fb1f26bde33c965edfbd2ef4256a90ed2a87a5199282671dee2e21b292071e057cf43b2475a35afc6b453c2e7d412968e8881c64dab8d41fecf5f0d71a8368856a7901255d3c15e2013ec70015f496e4893c5b35fbd29fbedf1c46ef9ef77002e8f3037616057107b6965c7e91b8d2cb5af34b32c11a21fd7b2ba22c76385eb421be7f2aa396cc1547108b2750a82ac7a54626082e5caacabdb5115b840fbd28c1c4caceb73c8576b54cc5f4619dbd58af852dda286fdcc582bc43abb12df2ef4c1d15cab3e8ca30fce14aa16fdec2a31ec71741c27cbc6bf522fc567ac64b0c15708fd534e1ca24aad0a7b0935a7f3195e3a352095e21e8bd305b5bbf3abfc0c51f5deb8cf8f25796f1d129809b5a4d4f07e7ed4201b9bdfcf582d926814f87a50a8a51ea16fe90c403f3f3ed74120ac5e0c81f9f523a2de2b27cdbef7e808f3f6384e70c16da9845d0efb86b1ff5f88f68281ff48628cfad8bfe18b75d60a5c0411f5e4421377f9a0f13a82ae385357d2f7f06689cfad874577973746f30e94ac52e5995bce50a333b4ebe2c46fe3c9ebc803f852e00b64d989b8919dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6b9a1ed5ce85d60922f66223b0934bcf41ebc04ad3fb1c9228f0bb5dfc094a5b01c741b67dac0f4f166474ec062815de6fdc67c92cf560838eeed648efdaa9849c747d93a38df277c9cd7fbcb6a0755f3ffb7472aca925e0ec76105d5d05d78aa58b54e4d3990581f2b39c24e022b416df11b0c38e7157993d9655339da58f45b9064d568fb835e907103cfac34b6563c5e6eed21a22fbf4ee4267c65a992e01525e805a8fc328794abbd2b68de08de78228ded624cc3e4f912d9a4d59a12fcaa178ff1871805b225eb74fdd13320e5a839c5cc0c1e0d4237b21a594f2a64a9b4d093ce3288a502fbeab765601e1cb955ff023f126e66c36bae68cf193f82de06e286f6b477692ae369ec5edae429ea05ee6f1b16c618208c3507c8b177887d83b5c8d5bf529029efdfc52bb0cf948229e081f2cb0ed11fb37443bac4dedcd2cc62c545c2d0fcd9b75b1ba4d6d8870629afc5481869424da96d7682e7d51489b15a20bf11a9c9d92beaf79fd332815f73247c0985001797952f0f73e5142f6e428b23bbd7bdf17097bb931c23438e07897b9b3c6c622e04e9963ec6933156cd0a44964181d0f0d637ab491811d0117910b4485db70801d781dce930c2ead19e8882d6376c0a2b0a33f5b40c2901473ecaa1a23e3c22f47efd6a31d37be63108996d23ae4b0ad153ad47c4a4d1edf48a0bd3ed5378b3d937fdcbdf138f4e031ed53c11e3ca9c5b0060bf2e08ceb13a3c7c47331da98424ed5eea134349e2ef4f43e02f82ebba3f3c9be211ccdded8be09813d86632083b807bcfe82cde66802faf5b54ee13c84abcd33670a87cef7a13209e839814a72de8c2f32806214ceee694abeaa9d80c986261e68c849ca16dcfd1d919bd441858966ec7a0a067ff135ac9e943d858c7f19c8101eda3dcbfd82948a38d6e3e2a5c4a4458ef827d792c590880ddb49062c9f11eb9abd6ee03a250b289efbc8fb7cafa1d92d0b3f6419a1145fe74dc4f06ecdecc3bc981f50b1daaa04fe6066efe04af91250b91765a7635bfccb514479f9246a3e49fcb9ff8e66d21977a78de8a80ac71ba4fe231f367c3523be917986f814ab18ee309b32fb46ba473bb081b37a3f73fcce34b36ee649d62a10a7b23aa36b63b946c4a0d5886e1f19d86d6627e9939c514b600de2836f872c563065112dc545c5fe39165c3f0456730bcefeaac60c3b5ddc78907a0a484ef53cae535c51e61340c056770cc96e619d2d7d85179cc8bc89470fdec99ef0f0fe17ccd8a2527646539bda7a78e0ea56b53913a9a3af609a9129d591ea86cdbb039a3baae1b3669129d8fc54f757823763c6637a6ad1c793e52123e830a403d9d1e33f113688b741a534b5c2b6f6dac1ef437e8c4ad6a956667c3994b6e073f656c4a0f416a0995dd32ccf1d6b4833981e198df273add1dd6a7460953d269b9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha7cbe1915c4cb94fc746e474525078a92d0fb6833fd533d50b2c5358fcb08910c098af0ac294c5e5ffff170b0e8f4b9bf7c46d4b8abfd20521ad03c71d99bd337576171e167bf520ab178dd9306cd0e4c2fca64d64789beea842b85d215000ff41f876c8a3989f0145b5111113fc383344900958b3d154d48894fda9c766205b6184c588ae11a67b6fff7072c113f13a998c2f7e53be5c92c3e08b4e0d1277fadc47c6a0cb5d4b72ed104d52974b0cebef71eaefef07dc2609615a7d5653b0176a5afbbba336d38ee3d0368dd1acfa5bba29b5b6bb82791f2b445ef2d76141560c9b853e66eb05dd6a87237daa2ff2a20303896cb1024286128378ad48c9533791e58a0832d5ecf4d93a7f4364ff82fa274d6ae98e420ed5033f0bd89bbb7f4e397007668094b7592dd703f9bc5df2eb128024c1983155ad0bfc8180002ccd720259ebc072ae3c7e568d9de8913796d1c2105d96e5a1211272d3236584fdfad251da3846bf15aae78cec96158470d540fbdfe3722ccb5c5a06b8433d24f424b9ca3f701374c1491ca5ae6c033a8bd8ab8b287556bf54d5bf37dbfea1c8cae13185ad3cea57fa818ea9a96a7bb9567f2242fc5ecae26d2afe38bca5d08c99f97d4dbea07acd8540e54dc5cf94759fdbadf822621b95dd93e21bd380a92b61a9dc3e17fa397518de273305fda5c653560415c7cced4c5b9599935a217f61d1984899bb230b0ec3511a8e64305551dde4cc29299c00c33eef32e38f42ad3958678e8b2d3640bd5f02b640acdbb1cd1e59e95c8044ca92be0f90a247fb11ee57520ea8630a958e67caa3f506337240fd77392e47bf2bb091f69b695c4b816859b0435ccfaa9cc5decef8b9d565da0bf9cc0bb504bd8c42a2fe908e115d7fb04078228d1f998755cada5619419e4ffec052705e7931a1475e6d78b03eafc13da362ccf090e1b1a36c4303c22e73090dbeb0c115a1d07fd5498527f99e4d237a1204c4214d852b753fc4237c5375b697ad0ea8ab68c88c12fc913ab20ba04b74fc9758d98e19ac2a349d08225c60acdaede024e44b6452927823aa96c01e9fadc347df840b6ba1ecfce4ac2c4dd86eb9f7542d2274532ca8cd85a8a62395c1e4776730daf8473d36723d73276e2b8e101aad0ee73207da402df433faa22ff8d26cbcade5c4cc33b14d99eb6283f6cb18bc033a8714694cb55e6fd14ab8f38b9607e31738eaacf73c01aa23e72c49a08e7fe022fac5142be24811f3357c2b8f47cef4076d2c1efdc18691ab32709bb61ff215f725053513db328189fa424d00ea4c6353a6e608ce2cbe2ee8e227a98ef52b48d6763c59577092a1d291e01809bdbe606ea35095113cf87c55f0d8243c488050a7cbd207018adaf197f76ecd87f96123a3325c309ea6eb4247b8f64faa8d2624498970d8f70034efc763215aea5044451f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h89f2410a174b18399b4eccee75640c839e5d20b324b3c5f0fa6a13e9c06a2bf92d590e78285123ba23d6c589f0ae3e293b6420932c50ae34a67fa61cb751ccf90821d69af062f965943840725a05385a86074f7507100790c45d51ff2e9a8d94df6df9841d928616512a54af0fbe3f5e6b601108f0a4a0a7eae8fbc650fb60746161e9679466b614ed39c33e51b125c3bde0c0d40151f58edfbdb50da6069dfc5d785da2afc54f9e185577825991631ec37b38316bfb93823f5cbbe18bad300d6dae1134074254ea2a021d5a55af47c2e89a20c086369ff2b676abde8b320314efcce4c9f91ff260f9e4433f7c321e409cdc9376fba4d9e6f4028f2bd88f9aeb94bb8ed53315db485e791343055d1c3d349546e1feda2370f55c0a256da6262070e832ecb5291a72b9e39b9b12b549f1ee92fb8be2170c53211ba9b348194dad04a50e661f348518d21cee471c82799492250f60d4ae72f5d67517871c106f4d6a0cb680886d4abbf8b1a777f3fa9c6aee2aa5a2c0f418000726ff461727940095adb8d5cb9f26cd985252346aef7646b9d884669a41960d436c31442ca4784bf04c075ae6c88a7ddcbbd860008a7f0dcfbd29d36c05c49b5be4ea8ff55b81642425932f3c7f6a84a70a205b949064f9448be053adb732ced644af5f087dd4c787b50cbbafb8739f7268fe12731ad2410641247404ff8a63abd91a527ad0379d8b3235be192175116f4c37b7d7a0e73f054262ff338c452e02f4eecbf1518ac3a8086f22543874bc93df54253a36370a56743811c348e2e28a50d5a4333972393cf3ad8b8bbfd9217b7c1d67a96ff100addc8374655db57c1ed81691b1f9de07851cd33bf685cb623cd366e0a93ff71c229c2290af79c6645fda906f313e96a2752c24249fae781265afb991d3e0a195645414afe677651b9b57bc391c3ea162fdf30284146e7e5c8656d98ca0e1322f83fa5971d43bafa1b5c772066a4bf90bcc2a12bb452a12ffd1e2d6821e98ce9b97a1853693cdeee850404ae262a2ca509b26ab8e039b2e0792d93dd2c3220e1f9e535c7319dbc0a0974d05f8c1cbdad145af311a0800e6d551a8a30f2c736e7fca80a5442f82b61e9a0b40bb7e5fd978926f95157ec1f02d6e721c5180037561159d5f1f005caad229c11208b9302ddeb7ebd898cc4d2d1dbac2d31da6bde74c9681dbcc230a8f24ea18dce622651beb7d204cd6a3ade72d39b29575be1255932189c0daa1767cb4e58b95c7056bb1cb88228498afc2b0cbb4739dfadebe007581514a40ffd7b96075e804176bc45d505e8139f61a58585138f4682c7fdff86b277864b67fe6fc0446494838492cc4c9a430e7053740955186ef74e30a3cb78c71ceca8ca56f5f0d81496fa6f20577c7fcca81179226e820005a37c7c6ffdac2d8f55581584797c2c7e9ca558313adc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd3a336c609eede1fc2e12d9f0bed346fbafc6c60eb372be41b1bff3d80d79289006e8ef3997d1e0c034766527c7816404dfda016b06f6309e336eb1a844a9ab80c5dcf65507f312a55b0327f48b364d666d0a9d5184d26f847788637cbfd3df3eff9c8e34f7e2091a3ec5596bd32d886c76bf8793e36686ae2964704eef4a26a3dce9d1153cf8ce9d680c289c3b4b87e94afb045ba371eb79ce1055cf1aee318035ef87d3b6d51b260e00351adfc19487d4baed658c01b0a96c20b1874e981619348effba5e47156a6e4b49dd50dde770f034dba4cdaa9826fb0461aadf314d169766d2fd3e7ed669a1af28453647694f4e768e0a893ca66e3f82cdf144ccc1c57a808e058ef4f3675fc3abaeed154d2200eea1ebd5ad3b3b4f482a00093d5a90ebdacf360896e35dfe996af0e481980994798e5eb5ae5a428123b9d1cf5aca72bac86e2dc03c4b72488ac53bf56e9727656b0df3131b96a73a96af81e13aa3b44ccff78ed99d44ed5f3d222943f6f48944543c41ead8f09888b4814b7d435baa45bd3d7108845e00bc400aed5dfd6d941e691d7ca0dc03fa73cb59a8d0ee536f0ad890bb557ac9218c3d59d437cb1662bfcc41257589fc14b98647e57bff3beacbd4856c308691e824704826fd2e638f8f9e9088edf9da2722d994de03e0f4f490674b1b677d0c1ddb920ef62525dd2a29095087f5af215be0ab8bb0632d68317c452aa0b969929d18dd9b368e2a5073a586e7c00827fc7547d0ed55f1336f8fb7ed041031fc78f1963ce59d6ae013cfe2e2b4328421660473ec869649d0929465a1f6a3350e49834674026f012b53e9bca47acfba8a7aff7bed53f9401964428bed9f68a64612826010c9437609d212c5c1fd9870f09f8e70d6b4b9438497d91f53b86c62aee4b497e8280a21ae1bb213a3fb6a698577bf79d8fe0fa80bbe0ca1e4bdab610a3e6d4cd5d1fe1921af17576352ec6337b41e2a5bf1387de4cff0a1276366056580c555750b41e3ba3fac309a0e7c8e33fcbd64c41b9dd03f2522bf2443d280e21a71862178423c9a592c4eb38cc52754bf401c5dd12d71938b00c1b1c9b4f14155fde3631fdb7dd85205d0d62c59caef26772a94423ca08690e1ddbe8bc037d5c2564da3d5e32b4a19bd0fe61916a85f57e3fd8ffb9bbc991f16503c0fc8f8d4c9024ed3d88ae7ea08b2564759b3cede0ba610434ea5481f8108f8d9ccac43487528b2b9f8bbe917cb8e8f23ad1c8603251f7ed8f21ea633ec340d792876ea045624337a157bd849d3d1860070a9ac3e27abc10f013c9807d3495cec3689583da37e9088237ff1aba6dcb29fcf7d4411658f7617611f1ce43a3d8dcd8973ab30ab303b9efc3532ecf7742e5aa510eea3cfe16685ddb74512ca03146545c895594685609c12b196e12b115fd4fdf31f9e4b6eccc467cf966394a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdb8b01ee2ba20391c733a8198ffca015f0492aaceea9fbd60b8405704de8dcafa8d10ef4db3051fc1c4fb31adef1cb250a2dbc5742bf743267bb8480c23fdc35032fda2edb3e6a956fa45e0185a2a56de28b20622c7d903bc16cb5fcffe01a6393834d9a1b46f2ab18023adb3f26e48c0ff0de9b9ea59cbe73c013c02bc24311cee2d7d89dbda4ef193b4e188d08bce4157e7df129cf73a50a792e8c91e4a7388ebd466c2669b66da88ebf35b8f35c72a23392eb47a43331b622cb9817db44c849e9cff09297bda4441f3b518c038c9b119e251e4455128f5e7381d0c480be4b16a6728c7a11292d6a2d34cde965414be44bca1a717f77bc2f7384e96cb45f3c3dbd21461f23923a789902d4a74eb99f230cc9b3901d04544225abdee72049bfd976c98a92ceb5056083e015c4d442eba084a4bac590cb9365b6ef54bd3bd942cf5cc8202ca0bd5920a6c4e822e35f0cedcf3e040fce19dfe563135deeb1fbe45318bdde30d6f16600dab473bbd32f34c42e5feba2283cae69a3b3661d4e6867e1e4057116f702e3ffcb0a14432caa7b88cea1d4514f627d8e57c5e174fc5002872eb4c4c96a1b79d393d1673adf9273dc838eb20f8de73953e4f38f4eef8220484885d1ad4b842db61ec3f7a967e196fa28d0ec9e8b52a896f9635c333ba449cddb4aa16be96d1a1c691db9f21e8f73677bf59aa87dfd235162162849bdf7c19f89fd1df2aad88b21039dc78b0caf04ce7ce705be9189a7893d9732bfe409aa5c086d3c1195089fa898c5e2db7d53895d0ef65fd0011914bc646812bb9130c5d2fa339a232e081dacf4c04300afe01f8bfb113a31d5c25fd393ae3cacd1c6307853febe5ddc3bc7fd5cdafb4eedbbe78aaee164f7f37558370e2dfbbb3901d8278917ad577b9ed5d773fed5aefa101c0862b610a221964dc54363362fb3d605e0c20a60b3f42b5801dea416302813738882ce1767251042f8fb19a7ff5f6cf2f529741473f5f41e9e25684ddc54a7295405e8f386887fba8447205b99e0bf96c8164a97f8aaf0811ca5280367db0de7e293792e89bad3e0e0a28016d10b7ab8d85fd88172d522ee63d3b34120fb1a555d2608256fbd339f70cf7e5cabb278192c402055cb6da4e116036f934b205d6572e3f2898fbf046a1ba94c35a3de15d8ca3b7de2ccb4d90e5d9a3042c69ffa24d79822ba47600b16795693846bf0c17fbcd6c66c3257243f2f6aff0bd7a3f3006b258c61d6e022a42d2abf2bd24933284c744dbef1809e0056fd01cc872f426c75c76ee9463d4d6f90ef87d78889efe275adafd23b533e5fdd95383364378aeb678d6d24031106951446738fd01b96ef3e17d3572108ffc543f3060596a5990f10e9cfa7a46ff38131ba1dbf2adb92e6bb7aa6a00970f44ea11585fd9dab89918972f332776f1c58834eae7134aa87c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h930c54c0631616d9c6d7b58b6dd07c08db04fa93bef7397c6f609f54b467f1bb1407e571505e009a39458230c7abc403a4a841d31edf527ae2b1aafc7f95b578861d4ebf2f0c46e1241faf574a467468580cf515387a7203cfffdd2c95ae974de5b0f280ac8567527a7bb0d79729a67bdfa01ca06204edfc21f9ee72871972beb0e1229ccfac1a1e4b9a9ebda8c65ccf3f29da95ea2db1a4c5117f5f5a51cde921fe48ceef6ee686668694c5cb6459b990d34bae1ef3d1a12c27ecec497e017194ecd465c7ca3d846b4497d23b81f4b33329c3b6adb14ce3ab0193c2d3ee2a842d66349b5a97997ce7a2b0eb3d3f85de7deb59deb321db5d06d74e6837e32a26defa63979031f86ec65a472e63b90bea2c63f0eaffecff3dac9f6b0bc4c1a17210b51d23206698eca3decc1b5f2db7021731894f67ddd0ef8ecf53457ea9f5d9ef1e2dd7c0321fcddd5c88a845f3fc1bebc123abadea44db9fbe5b719ce0865f50f58143bde5f423769166f20747a90068a6653b91f1518bf67e175326054c5a033e36f533e1a3f5e0814fdcdc7eddea215dd1e0bf23c5a50a0669d54e40493415a42675d41afd9f217260e3cdf2adfa89d7ddddaa3f8700907e3746125249851826f0cfd13e1c63b3a710d99f1bcae2ef638aad5fa8b8ae5abf00ce52c955f3ca2ad21e2025884b32e5d5329f767ff74c2c161e758ca5b16fa1d94de3ed51690c4227dad5ef8033ac733f80c51f6258d3b09e0bf1a9218ae4f50be7d72f653ea9ad46571c6bef4c910ccecb4be18eff37e3a9f6dcb993cf0488aede0911104e668e98bc06b434fbd1702ab9f03a054adb287f960a5cc2bcb74a0d564d523a6c7890c5d2664285b71bce79d4c8d6e04cadcecd64638dcd5b9e9c973dbd43614cdc7c809d4f16081b65b8b94cfa095be27d0ee120ac6aa54042e8b857bd42714e9e4c54f721e102bfebefb32d7b4295c50730b6d7fc35d4c731c30dea2161c026b6038b61ee55be4b4b642dbbd13c6db2f839a038e4f95f5e1917e515fa7fead16e1ea934d750cb1fbe07818ad827be9ed4f5824ee0354998e0d76cf1d12d0d904351ef60bc18e9697a34b6434f611c676fd0f5329e4284faa35109b2c869e038298d949b3ac84ce784a8a90c5863f0e544bf8b85380b1fff3256bd928c10b336598706e5cdbb9e35b2f31803ac5c76746ed2b035572d66bf60af705610fc839b2355c11ccd01aab88b0c61c76fa0a17c0765695ea408fe9beff15b14c1b0431197a83c3d4958eb3cc9eb6ee931682f216d213fc0ce4753583160ab5617faee795e2e7050a0079ef30d65c45063365524e958acd8ced1e38a43f72b0d292c60c3010f1b77d8b9ed8b736ee41632595f2cc5c83bcd686904600e5652e4f303be885ea01a6aa7339b9b5b4455ea2dd1056f7fc9769d43897ecba381e4f0a899ef8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h41f1baaafad3a0e476dd4426bb106533f02c30bef88c4d5406926329a4efe06502d931324cf074ad63bcfccf16aad53400cd94f0c163f3b96026328673e62f02d386e247000025ff4e7ac8604e90675175895388da641e22d00a0196168b5d150132b851deb7f071c3f564905747abd9f5166b8734300e66ec85051505808235a2d49e26f3bbdea8ccda51ca570dd38f46af7638adf7f07c60b7c50bbce3dace13721edb484ebf52b5cdc7203ae9be555a4e1eee8c6962eb276cb593b1ff7c96ce7e893d7ff4e6a8caa584fea7685b13ac432a82b0ad299c2f2f758f5ce8baa8723c0da89f1deecb5fe8d5360d5cc9d817f8dfca6bc92893a29ea576e19777e67f2e5800ec1cebfcbae1edd160258002d240d5aa4ef5546cf6cdc6a61624d38aaf4801250856788f91938abb5adb2dd50f2e17a97aaecd2e95fdab0574cdb73b024b3a2d730fea437033b0637b35931686c066a5e8bc77e34eb6a89f98d277838b06a65abb98f412b5f81ed4e4a63e104ae134fc2da9c8ef71c6a30fd9b22cda57f6967c6e781cc287c129e1e0dd6eaf7f6d8dad176a645a5417dfb4081d31c8cd6dcdc70b4baeb07ca92b3534b89e477038285c6a26c55af77d3fdcdb02b6f7574d3825a618bcfb905c7e31e6ff9a055b666c9b90e9e19c3fd4e186e50bab718a46758e490c58e0230badb790edfbf125984b8c5e2bf92c6e7004d36df8965572de821ec590cbc13ca716e733c18436e9876aadb742c3fe098d9fde352e6c33bf5b192cde10d5fb86ae4b632f1c1f6f219723eba58239586a7bfa96e3db349b3437637d85a2842372ae91b6ff8ed4a65f2d5009c0d6c4b07edcde91e734dac3949d72e9f3ac2f96255fcdbf97994873c53e3d76f40de7c8fd9ca47d686f2077c999e4a7f5dd6e368bd4283daef7a2bfa7c0ad69a9f4dd9e2e1c8235a659e6ddcea1001af9e42d8cc034a5a226ba0ce7708e44cf5f049ec97f82aa8f4d2b37e2b975a281a5bde3f79484fde0cc8aa3ca28e2205455c7e122a6c1f6c5a09f043daec5a6b6814e3e6caa7ca7166896c24755840f764ba16b3b7d75afe6979bfeaf437d0ca489d971053f24569e904b496dff722f54797e78ad06101f4ec0a9ebc0455df99fe2b855424bb90f7f231f05db9e124520e5e18360af77f3caa32a194421d7b8168dc97812361d8edfcfd6e17ddef2c2016e2951151455a0bb0896d3fd21d30d1670c2498d2efa4a1245cb489c9c217475acffa13ced4b23f32ecfb7d3f39d76ed492c45d92acb3bb7a62650337d6ac99968f61ccd1dd5fd7dcd67f02dbe74e682f9a370454a49a787132c827cbd4120bba39a4a853bdc7a64e9559f944ccf5957b2a0052fbabe927563ac23825dbf360529f9a48ce0648b83b20c8b8a8e0230963c06ac4d4cedf75b68688968988ce0606b308eaf1b4f0a337ee3cc31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h21f43858073c1c199a996871cebf3d1a2c2a7c91029ce3ccc80bcfd06700ba04b7ceffb6c394e99251d7266ba6dc9c043f2f72eac2adb224591392bedad4c799fe03656383c80f5d79cac673d41462b7042570a1a983bd9913b8894628e23568e13b5fd849396ac1f2b4a6d1402b501f0a538a64b1cc7d657740d78df42d13aab2b4454d2a0fcda3ee6f63b28874cd33653efbc35af8f8fe7e525d4fd7d652210ee023770d6362889c91715c3353e6ea80be0a08c40a72e687768f50512be72e40923f49325f4ee03799e89cf067deb7615728210c280c32403b53645a0745be28f2e1a96d68a3652387e9c5e81f95e933168e608d681d7f12dc6c8370a0e3287cf373216c35ca372f77ba13f3d9939cf878b441759e2be2a13aaa2e0c52e9c2d66218e695f42c52658dcfc4d0facd96583937ae8a257e57dfbc7db327b85a1755defe7671582277d4b9d6c823e484cdc2a10893228be7fca1e4a9049a046ece0630343610ec0f961fe086b2b8eec721ea5b466312e94b33494167afd04557c83ac0942266cfd0701facf25d8c0f710955049d8ff1b5b06dd2258fcc9d893a65925c4affe8c17fe69cae89387b117143184083a5e7c9ee861f8e40837882562f1c81ae6520be1768e61d3b9671513392f30a4af6f238184fa4adf55f6f47ca702f43f02746331cda7dc217a7d3aaef8b8b64b7c6d8d725a019dd4ffee4b8ca576bcfc98d105724371035ea313a3b4fcd7cbaf1d54ba9db4e233ae3fd63d49b42a3f59b81661c8825287a261e64f57fb1bfd95ab82266ae7ee8ca0a6e044c70e04d9cea7f4f21fc8d611848fecc64965cf74fe2e2423330bb2a5301ebea218b9de776083ea8102dc15694b9434f570b7f4912aa8d34a1b5ddeea75b93142fcdae3416599cc001268ee9c4ff00c8c50196576b610238ff43b89cf07b23501ebc81d4836c27557805d97e63b0826dd3c9e33368853c059d29108e25973e8e7f1af1973645247d9a8d8441f4cbc190684d65aa9fb79600b52ca3ec0815c1a3490ceea13db867d0e380fd7a976aa77ba1a3e18e488afd816e68aa8c0f11a26fc8b6cdb76a929a7985a14687ebe3978434deab883721173b14d4d21d523af1e1956e10768c1ce8d51bd21e375dab0d3d74587ec4cca821aca952463696907d35bc9133e8189d4e61013d960765a0688ede216e4d468615e701facdb12d9ff27625a36636d06048b475cfc44073eded611c29c8a5e5ae448c64f76058f36f6a60ed5bfe025d93ac8f67e039af8e738d7481fb367489de86c1f62935ce85dcdd0ff3671545786478f3182647c75c81d3dc9b7e1daaafc9ff1efbd265f446728f95d887893e4c819b08616c62c5de5b58581a7d8bfa61736bbb7c44ddf159b9183f293d657acea4ab35e96a33a4c69f4e6f5d3eb4d6a0ea34a6572fd67e30b3e77f3a09a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb2914609c1ee90c648d19bf14ecc289086d3250b980dcc2e37dd8426063c1cfb37103e000bd417285750632e1a0353da407768388fdecf420414f29756b8db012ce80ff270c273d8fd3b445717291bd8e2a25ce73b9d46768e5ea66eb795f9550e5df5d726598b24426b5b4849b29a06bf162dd72e949acebd369b52a9433fca08e4b6c8d8f1e79a712bf90ce03b8c4915367dbc5a983f548610d842965876292078dd745aed0dba4811c5d13092f322eacdb34ba78a8484c78c068e5d35b3eb1a5fb7fbda76a3a213fecbd3f644fbce86dd548d50c1cfe8ed8229182ee82f774416aadaf152a40c377c4b7c68afef2a3a3497db8f11c639e979f36da14cf5570ed12bfb8c2893c6b7e1a0cd9c9583e6f035e16c07b2f2f813a4a7d8322c2aa0e6cec23d85ed686b4f1d9ea1d5c6c3454390959a732ea579f22787873db8f7823940ad67056f4ea50172f2bf92bdc7e84cab7a65627524c5b6fa2531eadfbd70396b6bb107fbd0e5d92fef1487e5b336645aac639f673be80950025269f48e755c21a91812fe8ecbdd7423f6d642320943e5456f13ef87fa5c057492c72c8b8eaba48a456d741f9077db5e497c147db00cb8695c90a7e4c0d7ccc77d689780704751a3627339f01d1de7e6ca2623cbb1f773dfcba054855398964d23bdf4592f1c3928626a560100ab34f0f1f3e47007dec6a2b86615cc721977616fd6ae1e02be603c7b60c532d1ba6d15fe95effd89038eef1d4759daeb8be195ea749bfd4e40f7dc6c9fdf2c42fc2dddddbdb0ea101f52fb046a510d6d0307e6257fb26cb0091e55de189767e0dd46e4ffb6ab9079fe2a8e8a89790cda0cea987b5369ecd7c9dce6289688855f3f03c36d8c0fcd8114935ae7436bd377f4dd85c354be5fe2e183b7eeaada98f786415f384bee1a25895ab0e153bce0f56b69d903a1d4012e17a4c73e70ef33e082bb8e513f04b9d0a5b562968273817ae6af2839f5dc99a63a24e1bc00b67e7a693d20c44d702f610ae64607feb425ec855556c12b9a4e01e5a2a3532af65dc4eb7f1f9d978331732a9a73ccba8471b2e9d298fb3f2a7e26f6952be84ee205fda947cbb235af88898fe048868c899f1a4057fcb5ec833c72a5f1eebd5f752ee3a25f9c9338eb34b145230a4d99394d7858ea22d06182721cd04568fe2ee756049de777e8fa8e71c94eb8488f9531f35a3a134bcc6465aa760167a331314ad0210e3e30371471420ca2c3e55a5771c862bcbf587897ab30ccd4d3d9c3b52f9fcfa88264b6d1c3b0bd29000b3c5b3a2799798a1b738275c6951278ca202e763f1169552a804f2dab5caacfa1de5bbe50853fe514ec9e14a778427986980fbfba51b7832ff34e36c9964736d50b852aa14fa9c47377f7eef8ef1e3db279607abd4d776085475b079e16ad07ff24aa680df4d3e31b6f3be4955d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h613848afc16208122e535a22bca148e142129e1cc2a1194492bc75982e3d09c5e97c5aefaceb8be56f09efe4fdc6c523f296bc8c2cc324ff694325f54fcdf80a7d707e4b2a2a62c5b1b901591aa3a112edafb08640b92f9a018e2dc53e731f55d956231984c99da35bc442541008723539ae0d212967ab3442cd49249a2fb366c8e7b1819b9118f6501d2f96b7753780919a7ed38db7e4efe79f53954303ae8ce9bf89d6ba11960492dc0ef7ea7c85a8dc48494bcf0a23d3767021d832470aebe7502833e94107625c335fadea874968b5eef9aa909245038479d4c1fc676ec942aa4b49462ba9bd209309d4a0cff20f0370696681e1ca525924f412920696875c9ddfef417016eed1516b6a16f6467df9f5b362f366f267b368f2ca870467db6be6f1e1b7e52e6523033dcee7326fb5b82632bc8f9673863a90b276ecc390e392ca8e0825ec3dda270dd46ed7a0735a0bdaa673da1a57fc7d35f56be9d35a7ae9c8d94e1a4f94cb5eeb017360f583d0e71ed9cd2d721c7fa7927a13f8556ec5851b76a608b8406e80348c394d7081b26bb8af1c4db12d022913a7ce005d9f2f523b83644a1fc41edc0ee7989ff01624498e93756cbfa386f7c0764fa19a4c8354d759a2bd73738b88ce13b9594502d135e27c791eaa2fe394293829dac6da4818720f472eeb6cfa873da87f23f68de0b4f6f484a69f85b098b64fbec04f92fdd369608d14bc2be253aae0ff2802498ae3a99e7f3df8c2a82e7ba0059d7ce5e208296cf6f266f1fce3e9da12ff429cd5ec4a505d0f8e41836545f88792aa025c553ac9cdb2b4c10b9614b7c09f7dae385a67fcd1d33aa36d169f3bea43e9fe83f9a0b89c478ecd2503eb1001d9563bd342a93faf47db477968e4c5052caa6d4cddc07faf559895d94e10b08e6d162fd197426d501f6af2a659a10017eaa33254a8b6f815decca9a337d5a8c1a7465b64b218d62c0f300c7e4e5fdd6e89e84e656b208aa87fbc5183cf8f96ddb13f9e3ea5b2b17b84d36bdf81ce62623375a16b5a816cec6c187bb2aa42730abd76e23d4287474b8bc974b459c8a490e70a523ca66a006897103738fceff602f6c9abcb8134d454096e5dd4914eb304cf4c08b366e472d10377d0718263699bfc66917027fa51733fed8e14ed1ace7d54b2f8227f6536caa84b7ec19b08533101a2c0f503210bd51c0242a57f216331996bdd995bce979355a3b24c14c04ba5869d781f91994725c78aa76960c2428eeca1dcf6518ea14ad6186385a78a65dedc5524d8d9d5f58a61320df5f1b3ff0a33656970732f30227966488f609e2d71d32dc28cba5408e35413756a5c104ca86b7c6859201237a0e4bec7a85bc7871ee1fcd4acaf7a33c50c324b86f06cda8d70866fd927a16d461640f89f2c9cd09e3162d5c7f9167b443eccb6c1b4580a07adc488e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd300451a5d1963acbfd0b159c84495aa6b10a5c6456b1b9b4afd087648e37ab0cbd93fc0fea61d940533a1a16e9b828be75b9b19d891880bcb11a4077efc49a52e1294bb8a6982d83ccf631c4ef79df70952b1c6bceae86737759edf5827ec98e394fcf20a434cc17b6ef1fca9b06a66aa523d5b33bd4e2a21f6b2cd9ca6a78cc2760f73975f2490de6d77dcaa11679664d92d87d881c6534c939e4fa97bb4d3e3e8d0b34a8485ade0215405e84f6700eadd7873f379cc3eaf12d2146d8ebb8f31a8f766d14c1e1bf5a92cbbe01115b8e5cd9ac9b27a4b8f4f02823226b327b7461e2640773fea49cab173bc52111e395db511d9e4afcf8384a7eb1398821db5c6e95370d14b44f74c6c25d1ddee5dd92eedcbf7c35b57fe08ab2f067a3712dab86dc1df4520187190f0b86a08d7eee98c987b1ebbc469fe2158abc1e79c97484ccf64f05d1fd1b5c9fd6b8de2cd598e01afa95446221ded09b2eceab7cdda4fe6f43af7ca3ad434acb2c69e38696e51716f8b61db395ba5e156655cf515edeca04128b18eea4d73415e81f11a67d5c51ffa7581cda8264a88bccae2cb2023210cd5caee4ee2fc7b99c1f3ccc07539e6887db662abf8a8d66b9f8e8dd36a9cacc118938abe7f08d6c9a17333c21771297a4a5d3b6d330387b5638d041c299b91c031154290c1c20fbdece736b33ba62aa3f30a8574951c4b9b1f8b7b36c8f8295d045e3705a511c471bcc20ecf190fea9c99a4a1438f819087d6ed4694644eda577b74dc3b4640cfa04d22c11617983d6bb5203fc1eee3ba7896620e5e622c6ee26e68fd938283a3d020e68333a761aa4f956f36109f3e0f5a5ad73591dcb9ffbb3330e293cb4d71ed9791195d56f58a820e7188fc65123cf1b248f9ec114a85b2078ca93f2567e548a105a67a5d5143e866c1f7de979473bb5e9cf8e357413710c1cb1382ef61f4428f40faaf8f6e36007e7037fe6cef7915aaa2f8e505ee929152c2f7e5c23a6faa3f7139a55acfd9c81b672dae8f30b4a4b4e44a23489faeba38a7dca04c61f06854f6fab953e20bb2ef92078ba17589bf61f8267c36f1de4526f2a84f0bd25dfdef9e8752077c848ae99b26dcce0f266ed74934572232f5b03cac1fa046c0ca2858936ea4f092d7450e52b00b3fab0f5867efdf2cf4252499adabe470a8ea7c2008314b23ebb8e5c8c4a479b707621a18d91e55be95ba1c6f7b361c7bd424de0bc09a1d3268e2a115c89ef712a6ff9608ad77c8d428af68c576f90a411933ce9575a30e11cb8d9c6eb63780c32c560ca5b17a0ca94da2b108d361a5f6d73f69b9b7922eeb9830f370a99f5d2402530dba1bac5476dff7f260a31350951b7d33e32f4415f24d149751919e76d0add0d903300afe819debcc2950fcb21fd391467e2fef6558888fa289482643949b22353dfa4855431acf93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6f01408b9d1b3dbad2e5a7460141d1071a06fa7e4957ed18c587fcf313ae7fad329d95dde443cf3f492ca2ac2062447dd61694cbe4ece50e212bf9ef32b7a690d8a6332c49b9308c930154a2d3b2340b49bb98f2a56ea89b2295a9fd813a115b0fded27c12297b8090b1c80cd31e5966993e7adf30894b9ab6487d39639674ddc20e320e937e447230fe775fe64303f6e284ff53685b38f323c22d2fef1d95f20fecedea5d9217d50c93fd3a8beec3500f576bdb301fe0dba5b07009543a5b104124d198aca4824b4903039c702d1432ae1092ae58ea776034cc6364be3fc24892ba5e9bdfe0dd7d751bb077f8202a87764324407be8fc64c00d586dc904797aa3b41741f3c5b6ea676f07515ce6c77f3648fca57728a7ec795293ee9bfc228b038432ce0978fb1d89a66698c47edc6febafe43440591ebcb56b011c6de90b937e9ad8bb35a29f6d727339ce0ff6bb6d7eab7cb871abf2583d32e00b194db151edb71948f95d37563ebf0bc228817a05d6e5828e59b6e77627a3b51eedde4b480237d6a30bb918d9a0a080b909b371ee8e7e5a4532050db7e0f584d1ca2b677b46680a887a1894abbf788d6416d44c3693464ba6837d0bee68c917f0c9d84913b6b45debd60e1e0bc610089f9076ceea059f95f929525fb8af6d58c30ca8332d6ed265ac953ea66b2dbf7120e41a0635924ead0f00b85c0fb0558c090e3e9a3c6680f5658ef977dc687b871b7b5bb74748a53081752db7f1bd10addef549367d3915ab1058eabf34eb6a9e510e0cfc7fd9bc9ec30620c1ba4979d0c825f5b6c674ccdf4a8306d9ed3a2d1c3d6e64ebf837476a7999143a259622d1e93573ec33c2c55b08ae8497aa7e0a0c33bdc1d3404c336feeaeea6f2b062fcce84e74d4a83bfc5ac65b82384a58b8edd59880c7cc8a1a94f75204984bdccc4d24ccd684c410c16832be9178dc3e4a570cb4bfe12bb93ea976c73caf0112671cb716e345fbbf8cf15bb7da33820760ac5ade0fd56f1ca9befc44ced73c9b77c13aab95109b466e8d04266964536ed6584852c77514f879cf0117fe051e609eae50f565765aa267cc52ce70d8f17cb86cd63f913f45f3224f945f0b6afff53db6e36d7addbb9cf4934a3a7eca7d464fc84706c91b488e449188ac5f9385b23ca497592f2d28ccebdaef7943a5fd2737f82641d7af9a1c7eb61b35cf78cd6d42dae9893ac6a812c2273d07b68f5e19e1cd2c6b2ab3601d70d108835981ea11afca78d80ac04684f8c49c1e7764e7dc6815e76bc55e8bc7fc6a0ea742ceff2c074139f6c8d10244c3a4112e516731a3af8fc7f1794562575dc5515c2b882fdc01fb0c45f819520d68833fb13f23ce3f71ddbf52ef28af7c84d657b94ad44cdc6b04c8a6ab38d7afcfc1d9542c9bd7a17e31c5ec5b054075227b801eee399edbb05b55df3a04a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he815689be7bc45dcdde101327d332012bffd25d31b350462aec40b3b3c32806569a3315c91de0214496454f68aff2e01251657a151eeb919ec8441c0d2593ad6442bd4290a4e409bd8d5c059520d6deed5ba440203335fda3a449791450db1fed91450b0de8843e10657ffd8dcaf5334aaf1ccda7b89708f78ccf0ab2156d58009d1817f5c34a2752e26af8ca28c9c1c7ae928904a61009cd06ba64e63537bbeae00379416b4430ac587ea0118bc41c4e41ad03e84318f35a75cc39d3243f643c4f3adb47c34e2f27b88192cc7e79e65c3a20cf04be6e8952be287aa6e4df27885842cdab5cc64e74094d0dc14dd77e2a1c940b9245c11ddb2ddb57785c6a943381d5f5062009facacf1f073b1d60d7ec5a8e768ea304e2bbda2a1872e54147a1c2888e4510066814e0bbceac4c1a0f72dea7dd62e5d4ca9e72e5223dcd7950a112ceeb5cb4cd74e6531eec70bead405902f80d05b17b58f36606811dae1d64a60242a55f92d7bfe4be1ca6a86338a2ca3efd02f7e621f8cc4dd436217e591f4c0d035738f35d41dd2755a2c4ff48236dd5bc5c6d8e641827c980be7c2919b188338fea2e688e2a30599a423f6fc2b62db8e7e586abdc108cc5ab2fc1904a71809704eab0e848e4498677d64ec21f3ae553a50557610da22b58f4a5d754bbc838d8258552192e1cdd9189eeb28de213370f9717268667c1efd6147e34a7d5490d216f93770eb7d74369cc56e01ae71ebde0a43785893e880004322c1cce59af622dbff5479071ec005e8407b0b7df569da2b9f6240060f00f1732643b3762ab6c6b67a8b2f718caa8abd67846f5633232c371be41a5651905337bbe329f56abc022ff185bbbe59e0b01d05be7cf9e47b19e24a212c128353309a3056e2519dd06a90e1c4c72967c1f6a73944ac3a411a9c1c82378c328f43f6c3993acfeb7c418ece64674548eb88a0b99eaf90851807dc29e7c404119669e0152b385ef6170de43eeda0bfc8a120ccda36e7a0b0399e6212bbf1dcffb3e21a6d17ea70db31a7b74207d6e594599b94a2d9973abfd8b1eff72cb50b8c4924dcea40f05b54e10b4667660508db12f7f257401dca91491403735aaddad0b6410f291933e318e2bc6c03905ae5fe339613fbfd99fbf450a8677dadee8b2d27e10424dcd4f74da2f7f57ab5f950a1e010f41f3e64ecfef99655b61596c13ca4e7b18079dfe7c52b3be603a6922b44b6e70d9bf6fe7746ad8ebce583c8b393605838c5b1a36281891e329df94408b1d7f27d8fa02c882f3277ad422e6d9d49f44945b51c3fef5da60ae04c6d332bca6b4a0529f438c332303d84a949e315086d692f42b710b19d99090eb3dc17c2a847ef8716d3b56e10c0e016bf83efee6b45ba08ba098b3c8497ec49b932a2b35413ea371819efaf24e3220c4dfa6376e9794b0618336c988b53d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h17aa80c5b1c73d55493b694027fcf9dacff62a136b6a26d054b24a206196f0f6aa42b1f8461e9f38c067a41c7673485d2fb92d15a1b468ad6824e67a88594edf07a11d7f496b4ca7007e89b5629863ade0acc674cceda155bd4ff47471fc7703d7c077e09e767b350b68d1d1c004b76627955d1d99e3878e7a894d3881a64c121983bdef790ca3d8f5ac231de3931153b7eaf6e100fba4b2fff6b73aa2516850c50757386ddd8816fc45ecefaf058adeb645bb8128b27145e2aac892926153bf67ddf337213e91ffa03b924c6dd81c9aa7446fda6634a64f4d13167353441e4d7b91c68ceaee7e5542f5a72c86788e7fa5df96c77c0c93ee5f3d6cd8d21e6b3ede81396c21c93dc4f08571c9d8460d0b4fe4cdf09040fd774d3fb913d17da90610e39d54de4c9e959c55a290133e63010db96650cea82bde03a0ad119af16ac0b51e250ee5c72b58521387ef67280924f9588454e10d9e60a755faf1dd288d9639f231f40883bb6c914ed4c86526f23d3e2532ba409c2a48331563e3845eeb378ab06d97453067b65bcad39a196baa7da6b81429d2a267bb6a9696f83ef1dd2494bb31b8fc9534f40861421691977c1151d1df1204cf50c277aa16e3cae6de2b185e5cc0d8a041ce3ebd40fb1c79a26731db3c6e67ea01e13e222e96d98632bdb1e20ecf0626cdd5407e3476bca7db79bc78d4a2d33c3c38d711f0657090d3da839a700a43ef087810abb1290d2be8c881e3b1ac938f60a273a9a73ef0dc5a8bbdb1a72d1e07401b31054405adbeba1126df905976a437543058cd12386705428ccdab3d033d3054659e45b54c9ae2de7cddc1163e14de8abc338898c9b0f0c329a377b72ab19c5e903b165734a49b518075473d0684417f88340d5ffd6bc44ca80c8bbde6bfbe2a95f9dc747ed1efac5a92cb0bfdbd7441fdb4c840b9ab3865f7730958b016da4dd1c91cd7912bc16f26b58029f674e6426e9b14d8eda524fd6cb6dc341c3fac18ff8bf982085a42013a5535a44d9f2069108f777ecd6cf703476ea69b8f2544a5c5590f70b8aec77bacf556f879626bca39edced915bd68432d5e2f320177f5762b2777c15edd154a13fed924e5b1b5d719a106a25d7152ea3e2e6511656cc970574665318cd5272b3d147dfc33980483ff233e5001ac3409e6c2b950aab5c96c85bab0b4f36bc437d74739be680bd74819597a62de28ae088370e819a812aa8f724069e82629ddc450f9cb2a771b2ab5251cf96c8b15ff9e388f6007cb6b605689dad9fea24f1a6e3ef9668a81822034cf1c5443fb5731d5c151f3ce65532e462ecbc208dbfb086919eb56daa9d4bdec2c2e9e3245024d2a3183ee58ced7cbb503a730b1ae4cbb3a7eb8dd5984d5c9d1467ce6148676cfd75ba1b5eec81e64d8283b5e25e71085eeaf9bbd05e447a33b9eb7baa9fc1a563f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h78e1f60139f16181d77d19756d7261e90534b32f77d6509e04f9ad317b999585987940887c8f19a4b3595adb528e76ec59382e3f39b13be132bb7befe6d37bfc6c47a907785a3577825178e0c6bce2403676b8c2327d00f5dbb8cc8ac5d2e9754594d88a1d1adb50b24985100b78f3726699d307b5557e636b3b3be436b6a7db75b956bdc3332bffcfd895e332a7db826faffba7bec376db06a6f031fb25a904cfebd76149be97944f86160a251076afdd418649fdb2ce6be93b920a9851120bd5f44a08a9f3e134a191ccb29f03840a1c89a600f35c8a3ab3a80148272cd0752d512dbc9e9733609017dcdba520f705db4b8d59a90b945fc9b323e48e07ea775e86f502a0887b6a704565b009fda46811571f1ba3624b7e81bcaf2935008b9121c44bfc3d4ec8635e424227c78f41cea0eba868c13992820c53a111878cb3d9f737faf393f0fe28e047c5f3d879e9374be5665f687fb23abe303789292b5dd38be37af8cb88dd26b95ce46e6774fb308a01e725869dc40c7e7bb2c06633f3889f805ff66148f9c6c68aa6232a56cea7a628cac2a6be3a72b4dc45f39144dfcebaf29a47a6f426f0f4e63065e26a02679b53867785f596efa9c958beddb977cb02852cb0c7530bbd2d83d75e7e3c05bbf6cc7f7125b38e5d744fe166685e2a8fbf871701e9ed9fdc74914653382bf84ba0f2d9ee6fc3650b17a7e4e7a6f0d87bd38ff4fd202a756d3014e5fd317bfe689bdafffe116cef6beb4e7a5e42176fa75596f934c0e1bbaea2c81cb250239fed689f1c510c605f1d0af490fd5fff5edf08164b3e7530eb92e86658cc7e0e054476bd99adf16bcc151e9ac7b8d60ff477e9134d18539b2699e897583793739c41e4fa861d741be3757844762428755afd07d27d6791d0b46896848494c326a28ba6756ddba225504f1e15074b0032fc5e702446220261f55eaa5b40ff66627168c750a30909e1a1b5d35200ca1557ee2cc31f8fb25b74f08247e52781a1f6cded25d3a56587528ad3b01340136e4a2597616f068e3f7c5194de2643bbf10e9b16c9bbe177359c537f7ddcec3e59d050aac0ed2c15e3d7310e6141919ae532cadc267920533ea6aa65d78823088d8f89fd9d3f4cd039575ca14d4fab8eeb150d02c4f06bba4477e38eba3e9177d2d31fc8a2267775e5c7fc6ad21a126fc9ce6e1953a0218cf9bfaa2ceb9f817ae1ba74be7f495e873f8e1979dca06f88a7f013979411b24795b9f90c7a669304a35e0c16bef515a7679ef1786d4cab0344c9ca1b7a9a1ba5e930a3292d6d39a8b1b959a9d9c7c25c56d6de7198ca1d5466c3115ff0dcb0a3ea418dbf62a58f13b39aaa33c615f9e54b1e86bd08ed317431d70ba55761c249114780723789974bb3d4bb6a21e9fbbf5776c6632183a81893e4c7c3dab8736a12750a6e4e2b43c63fd6f0e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb025b43ad684d18b082aa0777c42d1092a396a69d9cd5d69d7cc660f74548dcc60f9ab07c35b8a3d32e2467730b02312d6145359be564400af4768b492ec632e69d2fad8353bc9f355185a1a92cd80ad61b3ee38b2e5702d70d520b2e00d244253f9cd634311ee3224e8bb62f68ce8e92882441b15aec8787dddc9a34ebd4aadb13063dd58070432e05e53d77985a70f0b6cb1f18334fb0cf00136147e265af09df1efe42bd92bbcb314c6970eb690319bd8d6ea7531e3b1a139fe2fe4ebcc8e299bfd91fb89060cc4e26d5a030c42b27db59487100ef1a3982fa7833bd29481140f28218eae07c279fb88a2e9a878923dddb28746ca91fa74cd0e269b6a84d8dc78bbd9ba275f6075b0a1cb511916b7a1a9e07c4058cbc12a3b0b708525762cab641ccababaa13fd8e4a7aedde1f7681c682b4394dc57eda956c67e831932c382dfbf00e2375db519bad06b6554f7640ce92f188b59c9dd31c7131fc475fffe15eb25f2d6970175957ba3feb08cd7a413bd04f02d7bce51d55dc33593dbf52f77b311c734f2880b6cc7eff2587eaa69941433001b46df84def0360896a79920d4c2673f4501d47db9c6d6ea2e4fa52755eb11d800afb04c28d4f2ced3c0f1c7539809feb766c7ed5621cef758bb8a70b3d63ca7eb637bfc9fe1996dc546f8c8fb1ce89214775272b45111473a15014f320da61f8b4d9b046c8d8f2e3e104fcbe686095e8ea598eef9db175dbf18f10df53c591fd0f1fd8dfd965f42aff43d7c1ed81ce7abd5a7096ff60f48e27ad3e594ebec172ddbb0476ef9d2c6365919bff3fb86369e3d4648b2522c634c92c6ebf80e848147daf7a1c06e1aa57bb9d1d4c232cb433ef09e507bd94db61b2e99ddc9417dff90078713ca3d0361221bb4ea593c4efb16c098ba70c3f29fc7e8107e0c24cbf8102705466fc1ec08e3c4cf75a16c3ef23929ccdb205481a8120a21e9ed9ef49f74077fdd3ebc1bd5960d4e0d8a3e4512d71e7d9f2c102478493d8d38f8fcec020fdcd69acc66e7482b2a22b509baff9934b91ec241512ef8f6d159003fcf8a31836726aabb77fbe1cccbaaa668e570c8bcaa32b774ca723d3a8a70a53300770876de21e7d2b1abe7060257c3a3ccad9bfe22d770f03d1dd21c813cbaff06845b4c5527f29cf2b7f8176b47f1bd37f9e948de2ffbb22c194176b071facc8dc9cec505b1c3f7fac865efe8299cdcf9da8c2b87efe5de9f1b20527e428d8be21f61df398fe57d5231dbaf0562e186de8c35b08348ca0f6fa654735f45c3e087c60777ae123997c07880a095bd917a884754c0a35feb60a9255b46b7281e17681303ce4d32ba1e5223e36174c0fb63488e5c5396de731acdd7297cfd601b2663b92bf52866bd5d2744f5c4f0403282ae5165b0aaf78d4b0d20a973003244474d16767e7769beef4a48a2cbd39ad7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h637ce7eebeb1b0f0a4efc06cbbf793205b924b12a1cacf129607c6d4920ba9b2cfedb3ec4e3cfb0c2a4e533c5f81f2740750a860d0109c9ff6ffb88bf479baaf91857f73c46712d0516f7dfc6ea01af1cb5e6bd9e3f0e2a7303fb2e194716bd2b1c159a8d67998e5a4b918679ee16b12b03af58aab176620ce900c8556e9dc737e27fb4555e07c6b633f13a75d244f236911b5ddd517ae37c118ff7a7959274911444e9c7b7dff8f3c54fed313e24fe9e1867cf508ac5f96b4bfa5a25e889582404b24c7ef839834b44ec6e02c6aa503e33469be3a90d4bb33ae787dfe3727c9299328d84c4059ee55d3e2b54ee695574eeaed996ac0e4073bd5ea2e94e5f9ccd65952740cac5efb4f27f3081865998db96dce60773c3526a7c3e229057cc0bf958fdce750109b26208f4d2c591c88ff3b06f6ffab0e02fd63909131e3577bc404c8c404fdaff9f88514e21b1f9afc212389377c92dcf073e0f2ecbc80732a9ac6ab29723f50c97026213c0981086267507cd9972dc06520629716c7f83dbe7605092e7355850bf5d804ad32cb942d839ab094b7fb0ab229db503846d18c1fe878584c3fcdc9b45312a3a2af553a468af44981d68b8000503f47b3a27b78ba86c633b9458b5b328f263b7b23d2682f37ec4300799e4fa81446a7118f0226039aaea10d2e79d3a3dd8f6750ead99f5ffe903181a0ca5e1e901e9c136ecbe1558ebdbd6b14dfcb81b2c8caf98981db4bd7389330732fa7d2e492cabd890cd5f39ceb6ed10796d63c2a374102250f389e28decb5deabfc7771764ee4094af9855b47a1c6969676c5d58b17cfafb2c300a406b42c0a1f378f1f4f20670c9ab802c57c3afa6c436cae41503c93e9556d594c9e9eb07fed20dd7d677bd4c513e6ba1f0707744ba6cfbec13a4f03d7141931291a20a9ae69a3335ed2213e8e12d8bb3dbaa3549d4edd0b903f3e2cc3be7a1cfe74f8af033d5fa92d3d88dc412c654ed12372c1bd944f37b09d09c31a6f5d98c00473496dd112291cd8d6f577e1f99be35b63b1346173567d72abd231809548e889215e0aa46ff897cd29a28a84db1061a196f9e4c618a48d9ab4c5837666cf608e2f4e2e5609dd9edc662a1d2ff48127d239351e3162ec6ab11f113511a1d3636b484c4351e488e8c99d1a7f7510bb5203014d2b74c139b882af98a273e6399cdd349f6571b5477c4e07f34622e37a41654158ac9eaca75382cfa2a54e90db405d3b8f62464ebf7c16ad1b13260cc6bd9ea619d27ae5bf09ec1562bd7bd64ecb50f10c400f21abb88e7a6243f44d0f2c3de079467cb2b99e0f1aca0b72bbc117ce2019b41fa792c4c46cb1c372a2ac1e7649ff103a8f9432b0bb04c3a088fa48b8d43e062719fa148fbfe0272f9352322fa04e9bcd319dd27f9c4893c7aba11c2bbab0fc805e99148b1f67336cb109110;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he96dcd9a00abaec6327c74187e4321dda08f8b64d3df61c3a421dc31d9b891a2dfed3730a10cfe7d146f3ff6ca4a41cf1f62e01d954b43aec0c8266f6744b32fa6387982af05399633d6e76fe69883afb7368be3aea41257f68ce29c886f2c107aa97421b480528ebd9c5199a678bec2a8b41615b5b182a83816df825940b49de00de7189ed32a43167e54180269c32d27199a52a963504b665775849a64bbad07d46d5823b187674338a8fed9800aae7ee208856313a9320b1a3d58d8cb3b58dfde96b9890df97a19465b2de999620256699c11d144f91a57171f3cdd66f326f55913b4c8ac70de1bc10091751ca0c183bfa048216ca735137b58685a748972b3f7fdcc162f26df47053ed5ab7eed4b4db574e203b33cc07c6c9afb6f508e944a2496160da2cec579ab7f1e60363fbc22d62ae18246be5b36dfe3ef5ec4a87ec12089440a28bc667ad05d28e925702a508c70fc490fee6fe5e2c8876670cfccd7c697dc86b88034e25a29812dc3e4995fe815bd5a178cdb73c8873192937ceffdd74fcf5b385ef8b9f16a86c7210d61f57a4b7e8e1f1ebe32b62b384217ea6319a5e93fb21ec31ee27e0aaccde3d48a98c5f8fbf08c122b67619011505375d21d958a96ab16dd45e6f4b132a8daf420215c92e6d1595a39537c18435aa64351cbe5b749c45e3130e4be582f6066a6917d6f5b6917ad4925a83374618e9a758626b17f163c38ac2db27092c6661cda8789a2ce692ae76f629043a000452c0214a3b47a5d39bea8170eaa147ec40805be5952ba5c32031a6b1387c29e813c6c7ec6c4ecf4515b7c61aac9ff9559d2b06fe533dcb22cfb2174cc4b4541376b9e6c588d8987650e7c85014970f6a6829f44eb951fd02c0f5e32efcbfd9567e1d198d0af7d20f48c8bf1a20636294c2eda9eef7b7361c2b61edb75a9bdcb3dab1fac6df8cc0ced5a3358e27f56402bb94998614c7b1bf0f8ecdec15e915edf9c39eb2244a3f1422c72702a188c83c485668e7815cfc84c18fd30abd33b0bfbefba85ea5c7435bdc83d31024f5ebb7bdd97011aa8e9181c84b953872c3328bd3bdcee9db2c9f25476379f6d8ffad8a77d23f19e5b07c127ddb3093b7da24920cc0e52bfa74fa4bc323637ba395a9ba33eb7669b7d7f96423f93913ed21d831a186563f48f1e2c97ac5b4f49b9ff2f79ea9d5557131776607bd026f7378edae2651cf3821e61816f75cdebdfb495507583c04dae7c2e42fea9cb71433ccf5b70ccef8f9fde504c1e77ef74f91701faa93b5ee24a266f9563de54c18b9f4ecc0fae80fabe12e62225f944008b39913f288ac4a90ab2969473b4511098db6d2d903a4e9b6195d47af79e748381577d12b75dfbab8322ce2b0e4d0e22c0d9c1fcd8b3703af8995118789d3adae1bdead6acdf6f2e35af7908fa8cfac2922927167b5996fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfe9075b80806e923361407bfd9d12e386fd01a5204467e9e19a294944ab6f19b43b7c3526c56383279e474d08de93b8e0f4225ed40971a62da3fb76347d2708150b698e3f15277a915510639a7a6a19e1fd100fdac7462a996af7040113a28165688002aa99ee94d79faf113b1f9c175982ebc6400ae47059a73489e827b320375d8c4dc54d4e53a5b00cf109f60f6300ce52ad400a949f2a0e9d6972c3c20e6712aa38e89325520977a78e31abdff00a61aaa63f2193cc6bbe87a9574629eb0173c774d61e11dd3c8cf450e8c66a486f8f322759e0e0c663efcbdb59e470edde25c14ee91df988e4dd7e65c4e2ee8a9f2c12bad4b1ecb9c273866a738f4580c9c716bf02196c8a86a4519352e852dc73ed63128d10ff0784c00c2d93b1b5eea54282953a24664ccbfec0f559fe84034ab5e6bab9b06cd13af1aeaa17ce8a2e25fc633df19b2df233862dd9ec2f70962ae663220d3a8a7fdbc5674d5770e74b4b208ddc32e117b111db7afa71b291c54205c383a8acef80b48738d34ce2de00c8ba30e040d72137a1d448eee1c60ed86a26bb602595817c58ce34693a44b026f43958ca9d75b8333057253f4d3f9256bf61bb472c31357d00c2c36340b9fe00f496a08e6aa29b216a37d8658c02f487159e18c58e2ab1e31c65ef1bbbbbdc76b2f982796bf198679e0312d1a3a8eb31c26f5a5bae113426627f57ecb0b65e1f3eb725211c9dcd610548bdd902e5ff5de08874c658f945d8a6d037ad7ce67ba86a86469141fe19700d3f702104313a41f7d7f78e02c016cd10cdc23b1e3aeb46dcaa747a48e7510c0844788257d645f58e318d610d67fccb108496dc6ec7e5799beb516badb42e2922b95489c249525e87d72289d7e16a9e788c0c671e21bce7145e267f27fda4e29f5e70ee2b572835c6afa22c5a16498315f5b47b09517de6e4ce79810220674ed0143bebfadb855b37be9201cbfaab26494280e1916b64c0fd4aa72824cc06d34903f117d11a78c56e9e422db5583e1215247b9dcc854ed268b344f28590546f78b30fc14e73ef7d0f048259919ac6e6fc07ad913a0a600cf24f5defe0b5c285ca47c8c75f9112073e9fe804f04c98de120bef61a1a17018ccd0ab3b67fb455f70f39c9831c00effc8925f8cc18886608522c6b4d4212e349858fb0b22864aada62eb4b8b1de3cfbb9e8786236882e4c47ce7495195f6d1c9a26f8c6c1751b43db93d643fc9204b85aea6e55250a1bb674ac65fc2d5de25ae995b5b5f5740d42e5ea0249eb34ba48397bc5a696adcd1eed5ca624e2f44c4fe367f37978e38dbf91a16a4abd5cfbd727e40cab04484f83d8d0f956f3cb400c3c95048935b093d2380263aacd0032f2979c8c3f98084005c410ddaa0d72adedbe12a3a53569161cf0849780a0b98240a4d8cc3084fae55a099901b7ec25de5c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb40e952a125cbddf922563e745a7d01173ffef308c2070a2bdaafe19c9e5c0bc2e07001a512add20b96069e8684b0cc6ad68f814a5a3c24910c74f5cc7fb99c73c48d5dee967b56872a054519a5df939dfc630c3e45656976fa598a27ba292e42cbfaf87fb10a4b62ecae22cec7966e4355c0655683a5f7a9dfd3f24e3ae6537015b8cecd0e2b0c2c5176628f4e5ff85298b681633331a88e74f715f6c86ec932a9f822ecdc8b1f19e38209f3ff1810d5eb36320bf7c9637ce9aba46d6dc9a9b3e5d398d026f3373f50d65bda06f88588bd9266fa889b3ecf9a2ab1525c502a67864480d121614cfc2caef311fc0d83b1531928bcbd28e764d6dd95e311b97851439ba47f7f8d7a4b3bfa7e71d608ba9bb18868ca4669b0581f22181596c482a63bdbf7a6b38a8d93aeb796355c58ce8b42ed0bb80edb3facde0088f4a99a3d5ef1c87e7ed356571d7caeaf6cd305ce5022ae8974d1bcd0a1c51d503e7fe30866bd9a07b5f83f2ce558fbe67d5152f471de69c0575bbd88882dc75efb30387efed5f4234c6a41e05021164e08d7007fc69ba645b98451ff7c28b84dea599a05b36a72a20e41f793ad2d004a07805324666c3d665184c37846b0aa3d83f1459a883f8557fd3f219bbb5d4bf0875bf902f9d14fbc8ae55fc6198464e5259a70f3b77508bcf5093c310b2725b5bbb7ec5225437faf209d3fe3db3f696f02130612cf45667effe70eebdfe711b85f036e88b76e1df9c3ff4a0a71dbcc783eb52b4c190a8f9cde1c69614be244f68eb5949ab29a6832ed04f7d56d7740bde3e85df7b28382c2f3e65e88cd83913e1930a3452aef945403aa74934b8d82eb7fa69d34c696ff439eec786dc8c14820f9b653934a7ef320cee1ce294217c59ca689992834db1827d0154e8660b54635c7a0e9840e0098c4b319535b92735b40bdf7a77aa3245a2eecdd1ef88c8ae35d35c14a5c43f150c37ad62e72f140ffbdfab3df2ca57effb5d98e804488ff02428169ed281699d3407fb3f13dd652738ae75152c98f1a362e35a070c36c6c9a80a88f64a961c91274fe088731effaf4990144c9d2dced3434bd15ab9e25b77e57d5278ab8087b955c2cb633b78cf6b8777753195abe94cad8f4ac9a0ca85f111ef208cca00a9b1e59812782a71dd3fc8f0abf3f824724290a2d539d9b63d5b17ea7c30e6fcf0a482e614d9723c275de6ff2899077d09599ded213a3872b8c5b799a1abc3d8e63d12ded63b47c1f593bb537a379709aa5c8fd8df3a48802eed6f131e1b7abafe7c4d895480bd6126b779fe6457e44f445cb34a9effe889a7303743af1786360c588e3d2804dfd8483c62f3f35644e6ea9d30b28d6356cd2e2e0c7f028c637fe2a53094e314de1d2c23849e8badd191efc44dc812a3797edd71435b36bc44a9911858f4159453a3332f3cbd654eda21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h61cc0f6425c3004f1a5c7099ac350b7fb853449b3c05e0f687c32515b66543c6114170554b5d4fd59b7e7514020acd2b47714087b6c10e7b821eb7463b52987707ca24808c6aaac9aca130de44438b39692599fed656388904003046b0526cc8dd6bb0f9250bd87867276d6d5ed46a0757b33069dd22ed4d571882d0919b769496ede66ba547cf40a393d6b7a21b7bf1661513ce8a8d3ae4569ba07ac5d1b73ceb898f17594d688cbfc0d0d0b31be6ba225fb6884036aaa2270150d11748af6998b01d54c2c0e4ac1843ebb39f028e1ff4af024cde192d57f6fbfb8c8fa13d691a704185ccbcc2a2133172cabf4479272a105156083d03969c0218592873afab822ee80731d4cc7b9877b88e6180f48391c9726c1cc10a65be343d19bcf95b7fbad629749dd8727db32244be14791cf1ab3ca4c312b768979ba1b91a3e4d2181283fbd9297195ffd464bbff8c5d5c275ad1972eeb507bcffe06f8f80dd9cb7f1b48c8a81b6f88b2e0af493b938e528134b010bca61cd7f31bfbb9df9f710f46e555b939179fce87e86d304df8b0b5010a2b1e54702b123833ccd9cbc4f44c569682b65b0fc9f800430f67767878bd7816e538cb6ed7100d37e37d9c0d29ef26759358bc627059640dda6c59ac0595aeed130f0808c5bdf0a3b73ea795033b38e963991f0adf63cc0ac5e5a16dd8dc1dd71ae9c3cb131b456594c0d53b9210e54c88ca11f31b2d2bae1178172e8cc3ba74f43b6dbea67b3dd6b2eb665455dd0340b91b980c3774cd6130830e1149331a89ee62186a3291bbf23011dd4d082b42fe5cb12d624bd332740a3d6ab5736cec91bb3da13453bd262821d3dcef2c66e1f24dffffa001b850cfd59f20d62b5271825a7b499283de14002d8af130be3e6cb96eae89f4770c8a6f2c45cf77b7d9de08d4312baa13f78d7291f29fdc6f0e0a2f7a19b619b8d0e3e34dd2a5ca19caab4faab9336b70f4c7c88c52d03b42cf4b5c342298b95a961bf893123f9340a0dad3b6da386e95d16226f370a90365104824111c5d781d248c8b06cab0543558305db4fe993a9af661ef6d94decefd4885b27f9018defcd8162711243bae3be9845375717393b565bfac4deb064fa11b183807d36030fe0137d166d49c95494548e38b95730dad155ab643ef160cc9fb5a71c91aa57d2afc9612e248324dd22e612da73a8d7c42ee10b58fd50e9a9353e78fff0027a37d92429e67a681d5faf9acd38ac8a1f17d7e53a30a54253fe24f4c85dc6024d09bf9e8d7fe751f941c538f3267fec7e3d1f6053aeb4aec50e0a7d3926e17ffa7f4f90bcc99095e4d107f4d89994913f0bf9453e89d6ae3cd9d1000503a95256fc417e10faf53c2c3602c1837c9f10ebb93b832e1c05cded41399802fa032e93ac6f8031d507683306d155d6179f9319002fa54d6d5e0ff2562eb925;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h104a6a174573dec97efad14b3ed9385b202963fcffb789626a5b62bf95d8a7f5e2d769f9e14902c6e98035155861111f0d9e169dacf265b477e77675d111aa5818958a8a84f26e0d8cf38cb186d7f93f7ff2da2c345beb1fe1739f0f983723058a6d14a37d1fb474a2b836bcffb38b2e3d3b13840ff49f9320158f80dc83d0ca208fd228578a6ed73cb2e195c174146b336b598482bb45ef46b59c7fb06026d0721a724ee794a590a6c8822ac1437369962273083056671c479a26224b46cc82f2803d5b3e4393d258ba90390159e3c5da07586281483fe1c685544cc6163dbf240d3f958be94dab878f9a3a9c879e60d313b34ab7d5fadcefe518f52280719464b8871aeebaf159c885a1514cf81b72b20e16ad8464ee37eb7c860db4c74376edb34226e715dd18123620f895ec0dd4458a2eb1a1b6a2c3a57f87089c4aba58b8a52ebf2c820659ade0a7f9c562b9f986442c9bbcce935b5d422786d392870a716692f8707bcdc4491325269943855054a14393fa4e421bca682a6e7b0fbb9c21851b2720da561c7d74447887227b131faa1e69ed90879d076bc597bb35072e5f570c64b1997aeecb624c0804b9740a38b2c8eec81d26efd12c3e65d5f5810c4a435886eb893e31446e3c5af96323ded7269e2eef18de5d7da2317f35d722256dd36f9f2bfc2f3ca3b9e11637c79f6ec55c0e7d2a4cb6eebb3f5ae7f4f9b9a6a268700817c0e111ac5a5486a21279c5036732290c979d81646219e3ef116b59d48e12bb335c3f86d691bf277ae838b57cf9acefead38617b7afb9d768fbf11ac7674e901dc963f0337a7ffcd8457f19ec34ce2cc00073f692c52be21a82c5962b6dc4920e3994bece9dea9bc1001f4fd6f3f84f1bcde292d251608b6b3f06406a11ff91da932811e52189bb1ead57b5cf6754eb7240747cb21e288d66b71e9bfb49969d20c9a6e973b475e7358ac22e7aff1c63ae9e220f77afe4b46cc6f3469e104e39aad0071822b4e725a2d7f41c16f31fee9d0dbfdbcbc4dc25b60d832bb35bcfb870f9354eafd50399245afa9d11f9bc34feb648947b241f2337f6cf6751e45f56c3e9b6bdb0505a3e99c7a67858d1eb165c82d2ee9111ca16271a7ebaa7d9e82e2a8fec5463990f99aea0180e2c2419df56a6ba0918260ae93dde7fe0a995de472fb9f9d011acbb96a936719948e8dc55c47fa400191cf5502cec860a4d06219380c07acfe48cbd9bac1fe0af12525a47c35443972d239152a140b9cf607cbd219f867fe2137d2f07c89180269856eeaf26aa41765b9e7a46bb361ff212b0d79aa2ce0caf4ede171b2e45a1d318f612f207d66888d610f53c475f97fa575d039fabfb42e45ea42917baf4bfd6985624a41f663d5a02bcdcbbaae4b5826e274cdb3028ce934266a7d403f5a367515bc0b2ed76bd3e61c7fd486dd54c33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7d57f25ce42a6fb4330da602ef88e824f52822f40996e2322eded062ccafa5ca8da6d4e32dc981395275b522822f2bd01093b2ca99eab098c7e2c19b305eb3b57c1d433678639eb7e4bf0c90aaba2e2a2660c3f5f6fdbfcf5f40c9945f6219e3aa9315b6ff0771810c0513b1785e8e323d9d36815a86d7eeb07415f811efd1b41b9cd31a75b73969aaf8d3e40c60df7b31bcf327ff0e5357ae3d8301e421cb8ac6b959f1860c10aebb74a41cc3a3275c693b7d3988989bd9679ecd28a608b70b3a292843dff15a3508a86a42dc65a52cc08df3215b72d944bd6c5e1e01ba3ab04b2d931fa5eb6a826ef599eaa0b3c2d4acedf779e2c59355e4e9aaf9a137599c3fb951d1063ac17b04eceea7b0df80c64a72015e885fead62dffa4ecf49ccba9190ac904344feb66d490b57dbc716178f1930064df07a0c4bde0ab5fc6accf47ab1f3b15d63b0671b49c1ea4e7283e8f138109442c31a54528c28e53916e263bcdeca5bb2d434f20af3e260dff79e12630ba9a5308a5262157caa5f6d51822421c314a478cfd0a1e4d928db64ee160ef747002b5e7213c3d6c90ac37d9c16cc061e1b2da5892770fa31b5536f03144b1c63db5ad057babd90c95a76b949ef9eec67f7c75b63efe9ef44ec223300daf1f9e956661e4853b61c60e2a8f7d0370e226ad7c0331a2ff53c81a35f3598502c0363cd3cf96694a0b424fea6433dec996f94e9820aa8723d435499232830ce5ed3fedcc2284d955b829d89d932f765e876292944f13049e9e34a1b72c423bc78da35f57d3a518f6b60a7928077292b44f6b707fd5aecb5c22c7d71a09f12745a87a195edaad76381b16339ea93ca2a652a76b54a5f30dd12e72836df148aef9f0fd9ed00db10546d82db8ff9048c80d0e22aeab56e68d7c8efbe817aa6f6113a42fdc907c40e2508c79a1c98b3f500c98534e124b22446d109cb0dddea95f839a434ddab78b826dd947ca28a0f25adf042402a9a0a5772c1725ddf25dbabe2de920b79296038d149dab4a2f72196e905970cd70eacc15a1e974bcaa7b1e92e5a81398d74350eea21b5cc3c5b5e33e0b0d156e9a2ed9e2e7b82de1a482f7aa0c9b66df89483875b36c88b234722718737bef38b4b73b3f8de279e1267440f343dd5d9ba9f5e281e9514dd1c04a6e1f20d0deda815796ed3d9e786c6fa5db6ee4114d58b8c4d0012e66bbae060c79f48cf51efb5414ebb2efc4e549781b64cae46b35708a5f985aaec9233dbf1227b65a9dd87ad37bb3d5c3282a5744ce1bea50bd7f836f3cb4d0cb95541e1b6ad9c2bc4e5337c76638694daacc406b8213a21bca41aff2936ab61d72655131bd1314b8276cf1bd8d80174db9635fff3a1dbd9e2503eff406dd32e13df9b7e6ca3d360d122119e7827c89f99416ea0627b6fa19a071d05533f1f51ab39dd1eb67f43c73b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7672ae49902e5eb18c7bbaae1704fc0667511083dcd2a881e1516257358554ca1f8690d992e9f2095aaa9b088779541e357ce06913d733216b1f4f795fe64474c3210ce3f618e667e834c653fa1d7cdd62e0f54656808e1c983c961d378f4044f4362db2006fd1af56090401af076a5156bddc803385ae04db7ae91002c50eee8bae5ebbb4f239e4e8e699153330f636be5a6682015532ec849e3229186c4bc9608730ac4f8c3e98e927a0bc3de19bb7e0d24fcf98b8ed5b30ce2645aac41027e879c5d146df9afcbc8bbf818347e0229b39afd93fb6c56fb398be7b8bff46efd991feebe391aa446b03ed3dcbcec3122456f35d6bf06e7f457d274d807db0758805b78fc458641afda75c9322aec8e8aff129ed9c71c25a42409edb94b38da8e2ec5a36ced1b3232b2f92e8ce53f7152ce4174ee6e92a056f4bd157c36f91b737e8e707e110074d89b2a4a36a544c1342e1931e6a5dc695d376554d60f1edd517e2418185d2fd6ccef589410c253c01b67350e4c731632bee0fc0a677ca34a5d52de507e27eaa1ef1f7c77d45e52b29235653d977d23c8d213e9fe3e2cf557840523f02f10dbb25eb4cf942d6ef5a1e63f7ac65986163e158928a2202ec08edccf1bcd78bc039711cf3d2de9cf5432275c395d2c779071ba7c466b04a39cb6a34cc119fa09b1d877d6b293173801cf3a4bf5b6cf6c601e3db79be34b0f8cbf15561173d5e7afddc436ee5246e10501c31b30bf22de4631680ebbaed6f8aa298e64259e199c7e08f5ea6659f8bbc77415595d427c714c7ea29d1f2d340121067990da282684a27d279b170c21f3dc5f407eedbfb0ab2e4d4ff6bd3ae1a60223caf9bacc8a66727e77e3aab87c77ff867f3d90d044f614d26352cdd97217734207c80716e96dd1e7b4a08ef102447c2c968b9b000689e2ca10e7128b91b993c98539933059c2a79c4ac4f1bb19f5b2c834087e7a85d49ad173ec14cf9a0d3580fdc20f8fbb214044fc620152935049529c42ecd75cb5a171820422c3afa287f5979140fc3780eff6c734274384954d496e15e32022e0d758648e79b712022e2d19b2675efa9379dabecfc2856996ee75276b3db19b30f867afdbc5848ff6be55538d1ca643f5430d06be3ba1d25b9149cda4111e760c806882a4fb148524cfa891959ddac5a3d0d63a1499ed80bbc59c12644f94848192cc88caa997e7527d30b2c2a1681fb475945df4d834c9c037fba3ced6cc7815be3f3c3b90f4adfd86b8ef53a8415ed10796bfc6a755372dbc85e876482bd75b562a5b5fa74324af18d4272e830a680844028524294410156a16027e7ed8176c753bb5aff1483bd7d5501ac0d842b0eae4fd382022418b9a7a475351f64b257540fc7c6d8ae6cc18f62e4819c355a4d222ef37180f4bf62e6ee544525090964bca5a24763f2cdb8078ac6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8cbe4330ca2fe68978f615238b61abb44c4bb8860b12d7bcd857f95d6ce1150f3d0575e56c65761d84d68c13def928e809099d73d6c57a1cec4c29204d6badd99df6981d82d1a27893dfd7d06757fa3cb36b5e50ba6b94fd37a5e9316984ca1e8b3163d64ac62b76fd539645aeaec72dd1a0fd3a7988dbc85d10fa99ad12af7c37f987b69e1e4f4cf645ad3ac46afc6b0c9886ed0d46674d3d38a98fb2f84f238d4f239b2ddbda6431543c179e32066e49153d04e8bc7003b83fe64003ba2173451f895c171bd52a368ba2c2b15abb54a5e487f4ff7d32d09b89af63b6c3f10126d5156c3f87fd40ce837f609e9ea20e0df77b7a4fdb5c50f882c7d6d967deb359a1fe986713ab17ffbb63b377538274547a017c61f0e0bb92115c2a3686340e64a41463ccf4cd224312f9f775e8742334420259f7bf09d33e89806b6d0ab09b75c30b8a0120fdf065c92c4d332921fb65e99307c7c62bd5784f672da2acbafd7b989eaa025aefd885723e43325a43e902c44b3c268604cdae539ae34fcc483f22f3dffe1da4b67c3e29e5f08b0351ffa1b2d63c10e0f9e3d79b0e8e3fb46b7a30fbd5e7b9f83205560660b2de74e577af22c3d9dacb473addbc02370fd01fbc8950f534cdcfeb5b2eaefdb5a2c9ff427983dd5e4483a26d12d65a2f8529a575f01a28a3ebb93b908a7d17788a7ad16cc01706f8fe1bcb5183a162fcbebaa51afa4193bf756fab3f3a8e335e733137e488926e565d66056dd97950245af0a3ad61ee59db54784a61892e7775afeee8e0960cb21716ab9c3b36de489aa0f4b39624707e19abe45966363c7bf95fcafff79afdaaf5db174dab5426739fe6491bcc8e18dd961692df3065872a3f04f5a9a7ba1c8a82b1fca6b308be7ab006130985c3ca6639d65cac024d7c154ebfd458dd617d9856f6e21a5348b0e4db33f1d38e9fd3432a9a39a06457d073dfeb8f0e488a74986f90639d22758047613fd40d9d3bd6debec1aca5e762ed4039f9a4862d3ac62f008c2a577407c3288b610fdcefb6c5b3de8a3dfc9eaedda82ca1f496aeca83e518988269277d65959213f8f2ee39262dd26b715189c15225d17b4ca6f58e5d548f9b52c20b41a684081e45391ffd2975107a9956ea81f43c42411b75d78d250b827eb6793712fe97a95ae5929360ef4b940ec6180d3542f4e11f9a86fbe9ae8912f83dd22e727298a2c079c4575f11bef2681df2d36c21aefd0e3a2e217273acb8d1b5399a2d3fa25a6eaab1db43409dd99a6e8b454a64e38ec1c084ec8c0c34a6c1b4901eeb2bb89ada67458c5d8bf182687c41d9b41d279b424ffb171076f0d691b5561a1d101f8f54ab4a0f4c6d020c51a6844af0d028deebf4761577297fbd2790e0334c0c9f130eb788dd1fed2a2cc252ff5b30f1bca69034fed08ab4dc91f8a33c5dbfb24896915595e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h34948479807707969d8ccc79563599e3fb499cb54dbe72f3d70620fbc0185ba40c1cf68f3c6765c6b05056bd6a48cd43bd0ee05a3358f5a5d2cbd62b9d7d44c5591dba4ddf594c31d1381ef0d4af5f8607ef40e55dce176450a9a7f3076b68f83bca8faaa3b871c8ea08c89bc4c672b802f817c8989c293ad59ec366999542467d8a93e202d27c4b5c05512d9c94207d375779345a5a86765a6874aa6b281ace503bd614e6f3cdd08e0887e1e0e1fd82e2b8b022015111da7350fe215b497067949f91b60953699a8ad8260b6ae75330a367f5ae23c6c2c7dc0332bf0c663300ee727d072c12ce1922bc940b202406929feed4c170c528d87b5cb13cd0cde77cf74d945376020115d73524db349f874bf548bf76cfc04a7d247888ab60ac7fcf73084fe72f4ce5edd87d6d7799d0d0524e4607e0d226cc29427a2e6d81b415a2fd8e0e416c8b18848df4399543377dd1845cdfacfaa593ec8cca3f2f04431dab72155c10639e1254a699bd2627106503a7ac7b96d488c1b3b60b370bfa666231f53e978641ba06e334226ae7af8d9710c434bd55ab72e8b6acb69739f5557a2f336d4b0f8e85d79becbc168e2bd7a58578874722327ead80fd24a96eed730a1aab6a623ee9c6e192021bb8c75bad24a26319bc66ec84695a9d7575658c5e11a2588ac6d9443c23d6777c3164c7fd2f9d088e7659d2feee125fe5fd61747c977fc0907ddbca6618f13c5359eb555ba250b5c5f96c539683779118e8d83b5f2e5fedea47c029d936b88a1c6215048fc23c3b54bcd90fd0ab5a562575961fc096b1bb6c528a6fdd58cdf0413c8deea52dfbbf4832c5884675b8c109348e0aabcefec096679d23cb6ba269e7142e87cc06141525895108b3a83441a1f5111dae406219890c21351c559eab832663d10cc46f7371f8fedb9f9f28eb54ac6aa90b83362ea2d7a9f523f622729ff511575372d170c6575cf972c79e8fd925e2c47223d1da81a5a534ff211426ecc043d5a62069f5fd6c575113a5183d12d979635741f932f4c50e77d5a625b6597c5477339b887fa5e699919388fa527a17753ba7a4ef75b3004fb5488e0c5e6bec340b73bf7a42846572683b23d8710a81e127366b7d44e6d613ca27d0a731c3ff60c649a04797941f479285fb3553d13054157b59aebce989191442c4ef9a6d4b427d0d8795cc5898b2ec8782b737235420d0d4201ce51cc3bd7b415423f0ba789f501ad48f348464808a7a1af4e2c5ba0f3a5afbf14c864ded8de1e4d5c6dc2d7c3b07ac6895429811c4bdcb9ede0f24d85983f9877b0fed2ed331b63983bc72d5511ebea4fd18d730be47c0cac98a17acd7e328711e3d5d0993c037e9a07d172db6b88b0d802072530082ddf0200edadc6f203f77f633cfed8587d37416d85f9210ec5dddec02ba8d07b42680f36b732b96d6ec3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2167ceb7dbb5d18fa9861dc7309da3637ea80cea796aadb2fba82582bbd602ed8ab929c55df40dfbb517e80b8c39180e7ff238e7298b416dcdd238dedee57ca1be467515874077395b74a1a4d32ff0efeffa8d98f51725571568d588ff3388f475ba8ee9c0af58b5ab6e46184057e9fc9da9d152c5abd24d30333962fffa9abab6496ec1572d01e8b1b41e5a071f540c7667dd24a3684be3a955d0cb517cbe7540f6ed19b4c95806620f6227f1f3f59c876cd7402e7b66572ae46de9c2bd8ad83bca5fd7bb332c55c033a2b2f9c079516a271cddc064a1e3e4f46578d361ab44c3f68fe955767910ee74950156463e07a503f5ef77fbe1db63644c67d607115ec07793613918baf2c805ab9cbf8a6d8eae32ee809514533e08c24bd123d8914a354e7477ded6ada8a93a7d71039dde0911e51b894877c06788a87d8bb14e8b693ec54a5441f0d58aeabd1488706afbb425aba2038ecac759de1dbf27f0a680973e84f29c887603383c9d9ce87e155631490d7443e5b627720eb117f0e46e87e02c5ab22fd86fa2504bcc2d9fdd67e9c688cb84c1d01d6b1a62fe9c463c237cbe8e4790f8eba3f035878c618a3bd7028886eeee9c151d39f4bc0eb881eb05a956055b6ed8fc9f700496550d44751cc0c8aeb5f11936ce15c7982fb7c3238145866e1616cf7f5901a3652b343faf42cbc528f6a7a7fb684b88e4693bd51901028881c504bd4383ff2ccd19b80a931196898030ebe202d4eaedbad76ce7cfd14e25bc2baea471eb6fc4074d482286b6600ee6ea137d4958b0a642947039eabbb28ae979872ed5c41dcc6160b6d41872f5237b6a5bd57f199f73669b0f18eabe5439cc43f7d121524314e0c0911e4d075f478123e509580f2a14526b229644b9f67a2411385c1b105b213cfd8bf4235b575c420b004fc5f5d07578a5356d928d63203efe6b0ab7893953adf14de1877a1fd36cec2198520d325474e8e478ff8bca77b74d9a562657aea72ddfda8e07dfbbb408efc07e4e5bee9d170f03bef19b24e83a995dfe5eb9359e20dfa3988be9af340da2d8c2c7824a5c82f68b68db820a3ff1aec6a0f124be0ce2aec089ebef3823c9d9cfdc88dc2d89bb6b0cfc714df469aff87dc4e7a259a3b178ab99bc65936b2dd0a47fead12059a928046073a57b6d18a49663b7b602ae900e853635dbdf773fe909809304ae75cf5619e5f64ade9d8bd72362f28cae84ccf8bbcc7be9a166c04e521735084a261d6781c3d11f375fd6425e24ac75cfd15149e51f3cc7b2be752257d7dccc926633158fc9dbddb00c82406b0fd7ae0e900fc18c430f565809e6b8d84aab75e6561641f9a20189e6646dc162c941d7a0a8b1663f119705277ec7f59a21a59349ba45ef45b15054c24d2d7f92d7a5ccd9be72da80706a875e268c1bac8c37f4f35dcf0c351438c4a967;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8d4af6b6b251d46853c78acfd3135906488754f23761ed3ae60ed4ff2c6e828112926d546acc36170ca7400e1dd21dce739fcd03d45eba700b7849820f1597c7f36db6115b2d0d25cbf95c467dbfdfeaf90ecaa18100987e4fd31575b7c0ca60b58132904752d62302d9a530aff66251cbc45e0737241a1b03fd2014da73cfda20c0d30e586d794088ab92dc519cc9803031889dfc883dfe4b8631bc630757dfa6c52255a16b374a59921dd46b798bde627bbc897544885703af8df57531c55ff1abd06a8b6729995486fb00d9458a765d41944ce27c853b3e4750f0cd1f4c2b567735e4709e935fea2589f93b8e15e430a0b9453e33e1e1b5cc7c5f4ff28974a1b23917ea85031611a6d403ac223f97d39d3c87396b49dacfe57441bd20774a7cf7caa355bdb49e7c6e405c205bc4a95d6f9dc09d1bf39804492787acccdf0be18396bb4a6a13079868aa728f3d727c09058fe0f792e6a4d3819dead8d6f5b45987bfc5cbfeff1011cf9690dfbcd481f72892273bfd49280e0fa79b418f7f4559a3baa4f62dfd852e6f4dd7605378db25e82896dcd8edf7cd61d7e0070f41f142fcd4cc811b270fea48b546e1b75b2129e4aea9ff8ff9156544b604d270f32815165487bc56421dd553c518d01d6906bcd30e831966333ad9aec1e2992d0901d769229c153a4d257c62c20f0fea4b0ffc477bbd6981a52ff3748db6fc2ddc1070d77b021ed96574ac07e984d9aa798e1b8ba9ddfce8086c6be94696459f891c3795ab5a1ae9ca2f23c294a21610d6bce3185a2fffa388b0de3125e9522727c186943503f302daf90fd938beebc521d62f65e7a142494e4f89eb856fcc5c87a76ae37d52069e5ae14f37b7407178286226f3139fd0198aaab04beb44f8c61f8e9b937008ce616fec957b43c70d2cf4e02438daf1f51be5e200bec1edd91ca3b46aa67917c523830e2e41e68352554f2ee6d3c606b5fb751bc415610f19ece60aecef1ea2615ac725a215033fb94f28591162e3c804455fb74b2f6846ddf6980be568c4082ef58222c9e16bcea6382c348d8b45f546c4f0f87ec8af5dc4c8dcdbe6236efd907e792927e68b8fcd7f4e9e2f636f630e5fbe75f48551c2553d396718e0950317e3ab769c46a2375704b59a172d80f046166b1c76bfe7d72f58bd08b2c3363f41ae7c41c99fe66e7846e5d9870c595aaf77775455ca4f2a60805390fc68eb3357daf11f7911b085a757232ecf88e5dfeb0c4d4eadb30745a49e01b42921613dd598f4389b96bb56dc6da5e88ae5dade2833d2b573f606021426c8d60a4bb3ad6ef146f0c4e5f184c2763e74d862a2e9a1f0dfe451672545bde57d26fd654dad46f7327b659ab1bc21d9cd6636b37e7e0d90b948664e1443b5f18e7c750d383b700a08562781fb3f8d6189f6590f7335236849a0da7ed5d6e4f6a777;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9f19037565a885272b171c1e1e4fef49ff586cbafba526b3a51858905727f34f73c6e0312ef83a24793a836b398ae751b02ff52d2ee92ab4dc758440696487449abf5ebeeb90a84a16b9dbb4a6c90046c189917de0009df724b008453d16c0863b0361fb465dfdc915f80336973778268c4c1352aa29dd3ea9e1978d02cffcec357ffe1902ebad7f02e65e31b6f34fe601c3f412aa520001714661fe34b862cd6126967485fd48530a27c1a61478ad10b64b136e811ea952fbaac6ea99837a272929df39b79ca22deb6f6893f60c491155f7b1079961c624ee513e68fff6612cf68cfde8cd386b09a5faa6898d79dedf0c1da5f4292190498571116d207172d674c82b6f0e9af26025693241b0b0613b1bd66ff873e332130b47319deebdf4dd2cca4b8e90fcde080e4d0a43931c4c6de2ff28b908954621a493a70a69741448dde089877ab1a2219ef87a44a5e62c317173e616582dc8bf6b348fd814afc94f33a3008e046557c403704d2c920c383a6d4a9fd283987d0469eec9b9ba80f51b2ce54f65ce63eddbfdf130973f5910f330ec2ce26005a890e2b22472ef92d0e161fb2f631b7ed37889abb8b6c582f5fc84e9b2357f794656c8fff363db4bd204baf5d867875297aac506796cdb836033d5b25f00515b5e31a8271caa0d0f3b6a0e94b6aca6174a6d2e1dae9e0ca224f0440ed4662721edf7193827255be70a4c2a87aa6820059a577f55ccba94060f5c5390e83b1fa3cb375d1b5faa7f696d3405fbde0cdba0cf41376d036eb63592f61d24147358517b0a65aceb2ac889f86f2c3479586efe50156d4be987dee037c00a6b8bfe0ac94e48171ac19f5aa40c72dd79646b23cbb33da34b6a3c5efc45a39a1dd26f5b25ce54084f6f57d3c179c739ef487e29b23b51a1d7cdc238e8c3a031ce1ac731d9b3d6477361296af982901d79161edcc5978db589b10867e81c47e5725075986a51c71e8b8abcbcf88b4cb118b573263883cf480896ea04177e87f7dbc2fe0db2bebd7d3def17ff08a6268e8714cb8fb2a22edf823f1d74e2f826a9f85221050f46d56f9a6026b6b0d14abc4a20c2953e9ccf32ada36c0d2c4a765941e136289aba9730752987e530f6df2ae0624df8b87698a9584cd0cbacff99b64822de3a87958b1203487475d79caa815252267273e805c73741ce6650ae62ba7e23f597c994ef5dc333345b5c370ea4731bc59d63b705eb0614a71d169fda24f388470377742c12989caf8fcd71e70de2085976c88130829603aff3665fbaf4e85f7f2fd091241c96ecf1b5d5b14832a194da40529b8c067a2742b02ec1f164e8450d293ebd105ddc7d28ac039515fbe3f40c0571e74bac5e510e7bc0dd81ec52ec543d9eb650a21aa214c0c317c99238c096d0960863d34de767bd5f2140aa7da6214726fd29466c306ecd5cd749;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb8e8df545d6311e1cf8b08fe7bfe1d8579001ea4928d6ec9f45eec044db3791ee9dff4b7f023c0f94e04023cfb836be896dbce3894fe9da0bb387bf46c2e826cf09b0eedaa46e832c8b8fcf17b0d47e61de48caf8230bfdae1b93819076eef9396b954ad2c1c3a1bca7d672e8c590159a885e0945dbec74c358c077d33715d89ea7bd354e2d07ad51f2177be8fc458de9934099a1799670ef218ba783de565c2e3dd80238b1f75151c925f661d7053676449e2159f9b1ae6291a5561d1eb1124e06cb6789af956d81916f9154c1b2cbd3fa3fcd1c2f412d47601987eac29a8cb3173fd5cb23ee63a3b382c7c5c74eae2016dd04a9a846b10f988f9c69248baf7b6bcc2b976f694187c2f899e58787a6060d80e081baec564aa4665a9e5d904b3aaac34e350cd350e6ec7ddb52e98d9ba50f11754c232452119e6c27a57d1c1d961880249b5afc5a0df2df2698e31b30829e1be43bf3bca24c8898f2b7ab1a2a442602fb3bba57c8c0d6ce4bc4315d039fdce67c3c743fbeb10b6301175db2d3f49ac4c033ef82606024f4583890e7889d91e3c605c63ebe45bf853a3b939ea0fae2d1506704528eea3e6cb7ee824c12521f1ebaaad77a16c9d089bced374546cf6562eb4b3df7be1f6b13426df8cebbd2fcf977e9fbfcb37d40445c3f557753e03942537ff2e7e1d23f95d12f05f148e7fb452f647b358cc5618cad8e99fcfbf308fc6c240848f8f2bc44b607cd11a3f3e93360a96b2c9fd12f93f1ff5ba4f3a37f636d9621729fa50f35dc153b49eefe34c740870e61c76362f2a271cacea7996a45f51b6989dbc878bf2f5018511a502779ba4ce9b8858312c3cb09e8dbb521b725257300252e1ee349d2e54d6ccac561670bbdab3ad0db59493e3cc510a6f8c644397a6daf55bc56fd788070f5bd536286a702253d0b9dd76abfcaab46170d15cbfeee74aabe809340a970c5937e8623b21493b9dc23ece50c90e5808467e5d76e672cf43211b185f112e5b611c1005c13b60907110be0bccaa890b002924976f36ed0c887505fdc1be5e458013c7cc2bce10222714a6b76e202d40c755876ddd0cd1489de153736527573dc87918cb53b4fa4f36482c9fd308b037f7a9d22d4563e493b55a86585a3a2237ae3fbe872f6618dc8e930a15bc20cf8e157f3c53086737d7b45174166faa6fc373ddb3cb126b56e51a4c08a5d1c1dbde96a4a606d6a87418016d8ebc51384f5cc9dae94a0da7437e4f052581cb85bc6383b194453f01317a7929e7eb46f7cda39ef15d746e64173394bdb1b8b64901a157fafd16437c61b8f524732f40869a1b825ceb2d8b40cc6ab639940b566393f867b285d51e22455bd6cb7f52ff69664a280e5638edcac9070431aff1f4ff7377ab5d598e711927d94fdccba79c5442c4bf051eb3609c9b6c293d859b2164cc330b64b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc20d6b79b503aee48a23089e0248229b1cb60b3ef8b14be5b6307f8448539bdc36537bf28dbc18561d258c4140358c264153cee95354a014b214ebd27b8fc0368d41773dce4179c67ee55a70de46bb9784cffda5fc883ded5708721d941d2e4df8f89550fcafa9e0dbdc227a96270f955f2d3324fabe6f07027c59ad926051c42621b4f261c96206a16e6d489d924ec45ee9ba3a4476e2da353264ee857921fc131ec1cd8e6ac44a0fe9ecb4b5c2354d5174162501263901e63ac6175f3f23a02b0b35cab30c5ded68a0e2f7f9037d1fdfd3cecb9b4cb481287695e606a66dcec764fd5038c0e2567a0764680f9e1e14ce55aea7f846e20e312b5c5d8d65ec29e4be8642b59ec843f5de1400194201bf487b695470748d49de0341e63871ee662b787077dace35a9553f3b55e97ed8635b39a75126684a0ea3e3d473403cfe51e36a70fa78b762d6f3104a1f529bd71466cbf194c71438d86ec9c832023568eb8be8db2c13561eaaa3208c687054c881b8f25eb25f9e65ea1a1cc8de194909aca25e32ae0fc5c72f8bb47ef8652bc18d2140d21594bd4ec0c1b991a344e42d3f2c941956ac94cbf319f54fb3ae56b06ad6d52e5050f56a04705b604e51c935eb7964a5d2798798b876c2fa24e48ce9bc9eda3113e5d61478e92a996def72d6a0d0ad2f7b0512452838cc64792df3cb218c1cebe85e70061089acc8828439b87a9b7bd76de0350e29d7f9b2c051a142839f4d1b9837ba251f1e684da86257a09f1377fbe99b3e77bb09dbafc9556b51d57fa98f74cdbb282d25645787e4f723e943f8cb80add9d473cbf5b10d1013ad0de347b2274b0e31cb7693765619241b5a7b7014ae908bb73d8fb850b1dedc75cd5a0ee5ca6f1c8f2eb09d699f3c8eceec5833429dafbc87f24c13e67f02c9f06fb04f632683d9179943ad6b725cd16c531ee60d3a6542e12c8b67a8e5efc534cafaf4995e517626eb186ea47c83a8d24f51cf8af4a569bd3837dc775b71e22ea9e34326bcb458bbb44544c852da46a7a689b482677a0f874ccaebaa3cfec8c8d4f84c073fe041b6e63bd899187328780aaaef04335ae700546903cf7ad68d9282efb589338a112a1257fad1de53c19821d955b0dc34b97411d08c052f98536f8c911fc996ccf5eb391efec1cd3d264b6383cba0fadffae73465f89ff766516741ed7bea7372454ab6702246ae32149697e4ef1d813e1066e75d3986f1e7df3def1ee262889e7754c0060ad086630c64a0542a0dfada6732daa36c9e396fcf070acf206420650e77b193948bc93d281d72b9df0bb4861b36963d98699e7ea0001d641448dc7e711e92889680924da187830b59c0e2b8102f29ed564ae65b6f11e94ba2caad16a6c73f24c6d405bacf679ac0a633a88042ad7d19090c2cdb68eb9f4e3e928543e0e3aeb9b872e570bdaf4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h21a9fe5a4811bd0285ef2ca57166b1967939c00ecc5b7212a6a62f0eccd01df3f420ecdc050cffc59d40acf6ff432fbf4d505483bde8d008d0a22d0f49d3ac1c79a0bef967ee6e556281b703d0ea59305fba933e0ab007787b39531c89988211a7e05f899889a764583e5d3789276e8535b85785210b61dc9522ee7a9dd3967daa8131519b712b4a5c09ec7130c578842218060303ecd0317337460045a65ec58eb708da48c78aa7ec84e2ed338a47ef5930336217d580b112b4784cd997032cd8a9233aded7c5702a2ee32926db1abe1af6165459e12fd2973ff3637e40136fb0c128a2fc1e530bdfd7b6fdf11e64739ea2ee4e898467d0217812db5ba074f60b2160be986bc33eaff8b3400624e319e7e41cb7bdc2c80e480bb725d18c4abb8fa17e77674a495267c7777b01c3286a00a0382b2c216339dfaa007151700a363868511276dcf0da0e5d35f38edb53b7fd0d0402aaf86fd7a04f1266f017cfbd8bb1f8fc71fcc72ecf5f553236d368b16dbbcc8c3ec7dbdbc66b77d45bf504f06dbe9d05543bbd78b2d820a979c5eb9fffe57f93ef46a418d2bd1438daa97df9d66b70a761c507dae91577d2458956560788292ee74028e37558e75bd63636dfb25f2fdeb5af4dbe4c32a7d9a94eb6f126e93dc650295fe2bbe9d77100fa67c79bc78ffb969e8ba578d1afee23019a759b2d7c35768b0479fd5d28ab79eb16f328ecfebb3bc6625c2073e45e9ff20712a1075280da2de021d3b71df06bae24c41e3e4ff68c424da1ebf48d81d9a3d9cc3be576a452ab97e8ec38e394b647c3a95bbf63fcf90d4ede2a5e6143b33c0bfa851e9a7324d387c860e0eddda539ecc032882331336752e4e3c8dd14e4c6b73f1b490693c59dc31ecb06f3218289a46197b0762e10e56fd1ab6143c36e0d1b76f446ba6715efb317cb7f84145da4f288e828496d65516b21a4b519bb3bdedde4c73bd45c83003f052353f21ff6a0673646e68c3f7ade8833d88a6e804a74fa22b05fc756ecaa17c9f59abefb541b93a036a398f34164952b396719fa8e6b6f573f7837b05a9ec000d1ccec8b57356cc8bbd357d1a3a5c3972d359a0955435caefa4dbfd838622fd500a976b4b816c2a2aaaf84125a28d29c2f7c7fe38a512b9fba55bcc4498752f503b1147559662f439bdc9ca444422e737d5c1ea16285602466b88e8cf8a8f7f66d65c53d33ab15217e527cbb95382e5b710a93290ac02763b5b78c776b5db0575281aca4384f898b6fefa515c182d716e33f8b815d33dd6d5a86c6e18bf6c6727bd5d2eafd94da674379b59fe88892639ab4c76c7e790c26d6f91690d2b6f6b7376aae9561bddf9a1335284961239163054ffd76d774ac9508029ac88e5dd791fea07adb0ea3a12f12f1b0a9f40192976e224ea83f173bdc3ad75a6374767a0f6a5f02c95cf97de3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he2147a2156b53d3400c056cc651cb70d22c00fedf7f300e1436b4ce9d44779a47a5f5c54521b01b7c60edb7b5a06b977cf82a90c48a19358ca7eb452f8fd9973ea9393c2378c545908f7ff1bba7abbe1a2ec538dbb1a12bed4e33cb4c87cd9452cb686e9165b5a86f6401c959f4da238fa902feb895fe6984c122958aee68ef9676e54747944ba384564c574cd98ac4d8c33a5ba9a6748f4bd916da19600bbcc944d5dbb1495ba1681007a2cec034c0242a2f6c0140126b1f85c70ee40d92432a5a7c9f11f1cfbc07a4248d3207f7cd9688682cdd444bd4d89b1cf8ed3182566b09f32b341bee7bdcbf46b5ed7620cd8d2df3033efb7c4ef30e3f1cef1e21d11f95606dd86abbd341cc142d3bf0146f52c65044bad48fcb7ee229835e5f6b0c27cbce949565ef7d241c64fcacbef7e9141449344471aac9d12814e119de8545245bac60aad6a05b3f041df4e681fe9df953c162f210d0f34465ab4ef3a0edeef8303fffe9f3c0056cd7b33883d817822afcb699c1ae0370170a2e28ced15da6bf02c129ffb34ae88d00131389afb14ad25194868b43e5ed4f516ef139ce9b62e53bd057461e63b8af34f01301346514554a8978a4d858b47345d58676059ad64defed076a14f7bbf70c12a2fb38eb5bfd81c7237f478e0933093e1b7923fbbc25bf9abfe9fab629040d9e9ed886bbb62784f0d80e2af8ace95b1b50c9492601ad0005e56fd54ed0161fd5b074b4e4d04ffdd641744cdc27e0f34f330a2a27805579b9fefad297696ec7890775fe473c69a4c6d9ca8270e258c63b29739e1c81031b9939ef3b3d052eee7130373a099f8f998a737135424a28f770b03b499b2b87eaeef9c603731abafea8b380eaeaa3efe3159cf25c5ac77d3117c58c52b7eeab24b5c53c67d086ccfc36cda24aecc4bfd26f352b7c8df9062c9e34a8e9d008aabc50522d39674f1fbac487673b5562d0440c4c5d2cf8fc6a478bae6b57c0f7678efd549bf13e2945b1b7b2a87caa6b963f3eb45dec9b1fe118c1fcbece99da3f81f0b39d46ead5adcdc7eb3fa37a9a4c2b4a3b6022e814a8acd29d868ab975c43e6c450db4f4ce71d06493c401be44fcb32d79ee018e272bf56c16d76983c46006254e1baf3423a9e4ee13c1bd4bab0838a00247763a21186ba0754f5220895b54cc1b85235d91d694fe618b4dd4a71faa99274402ff4ba9505ebf78d6a7e178760670abd91ac6339b0511c71aeab7c733293f23e25f2f8537f720af2489ef941d94c5c1559e596168fe75523e82e075aa5b73f041702d042ab4f047da2bd1f056f736cab81c54beca925e87a6181afb3bd85db0f5853db6a072172f0b02408119d297ac9f370abbc0418b211afa0692517a601f2a84588730cd3fca4bc6d0fead9e06f18eb2641a4d2ba07f977a505d0179adb884435c3cfd4ae62e5071316;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h788d631878ada871dda31720387e05113b5716125c1b1bd86789219ba3e41c46953f227776202a253fbcf42c8552140341d1edcb838a9b271d1d33b56c6730030ba4f34b7cae1bfdcbd678eefd49b76e4e336f4f46652af38df7fc0354a914d2097a2ece7d0760bc24abdd7072123da6414385dd91198f3ebfb9c9d3096b8e1ab9cba1912366efab48c41104b38bafadba964de89dfa5ae98bd9dd13448ddfa85c1e5f60f98ed2b3fed2abe3426467591c11ccad50ec40a5f04d9a69d8fab02e8ca7e8ba67e9c4c34004552ab81815d844d38901b9bbab134259edb7885dd412a9ff8288895c40fa311e653007fe2cd68d42b8efe661d8265dc8316ef5cec21a6f1ffbb1017e59dc69ec3d39dd5073ba3fde1d24016a95ef43b8d104a959d741c8f46ee70a8fb8b5e8fb8e4e17e6eb431bf558944f4a7aa4c9880e086b7ac8f819328fbecfdcc7ed3b054df7a19fc13ac1d01508122ec9b04e448ac9e13afd65819c80c095fc3b3cd5de76eaff585815e0d68130f196669724e74fc318b2c4fa318feb263a90989ae478a0516107681858344787021ff29c6237dd074231d5661090d3057b7d8b5d9bdfb68dbc5b4d370fce1aee2366ae880e92ec4b2748ab3102bd6015d4982d004369e94b27e20c13be250fc41365d5f0a58603d2067c2a2a9fd33947d7f1a7678ebb388e9c079ac19fb98ad8113ca3220aab5d925c8c082d5a1205ec1d36aac3a2aef2664e2a13e2c3b474f360e0117be073f55b786b07a5a10a8f473f9c4b84f1be09b7adb28e96d01c8185cd77c0551cc3fe6d1b2d090bb07fa937441319c3d7267aedc0bf4a39bc7b359561cbc4750e6e98bd46d353e95fe8c4483240a12338f5173dc1a484afbd3b778d9a573d68c36ca3975f24746ac3b7d0f7b0c450dff6570326708608582de0af8dafbc2915e706f990af860038e1ae30231a16c0198abebbc99401b99ed99fa090dbcc61b810af270e3a8b757a04dec9710bca56adb8684b1ba20db0309f8e0bcca4c180ac25c4783fd9ff7d8a975a565fd718c4b6f686328de4bdd2ff7095bcc25b0065e22f0a66e56d3b667b881a263b2cfa88b50ed13cd6070ccc0ce8910f54ccf82d78d21807040fec5f2200e8b3dacda858b6f3c1ee3a6580b9aa3a643ba8ea77fafbd933a8f329943366ff814f7f6234f15eb26cd320ec4c89d04041a703b6fae5fc552394e0e2e720f9e1f0e796ffbc53b0b4dfd036adcea1de93fd11d24bae97dd137092f90568ebe35204663d0f0d6fd25f0bad9d10eac9fb437091e0564aeecd6ed21836f11ec88184da0a7963a8fe5b3dad5a9e5f73e880acc3318b196dff277dc58ce125dd1725cfc58982ddd177ce68d2d1047bcc5204ef3aaecd1a07473eb4c49d65b53a2d3e328d3e2fa98782d243010a75ee3f17975bc7bffa23c06d8ee9b3500441881e38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ac70b44147da72d6fdd79217772cb31021f8af7a69e8cc245bf90b3bf2021242aa87256428be9fc3b7b83cd809167150853144d45ba02dc8c052dfb00f148562e67fb8b63b54be286eabf9c969a09ca7ec35a1c8977f9c84776105151e81774e9a8cfd82c0bba75c525a98b548995322ef13b7cf097eefb9f3a452aac570c410739ba90e7116e845600233af9d18152529ff70167fe40d48ac3230061da17336743cfe8bb896f1329ca5d829baf1dbc13fdcd5e7d4254ab0ee336d9ad6979245ac21ae1d2ee3dc94904a152f5677b5a0eaf1cecd79ad30b669d0f871072392c43a8704849ef67ecd4838d32e69551f405e7c24efa888cec0833188fa5c42ce06f836d66c8ab8499fc3065154b73d6729171bc580dab0217e40b4200497c9e5af400ae3839981c7219f6cf91802ea38abc5f2044ba203813ab9b97e85c58322b3a935b2ffebb2c4c65fecf38f24f0eb3a36165e31b59eaad62c5af6b5e39530a66bad5aa7b4cbdefb8a9082c037b0215e7cd5d6510af449c0e5959cb6cd5b61cf4df95d1b36e9281b4e27045ca9ec9a748a4510b268bef190b5c6967e38c611ac3787ab65d2b332b0f5cd711169e7b38cdae7a0b3623795f748f7fd3683d31431239c540230292fe6d8c57eaf490568a16e05c80972ff952edda40a63d647118ac70bc2bb8ee8faf606518aebae4e090e5e215deb79450d201579002b3f6f610a6ddb9bed87552345ff0962d67c61824e2ac9cc3a757bb2613af014b37cacb9ba34619f372ba74d0c880012dc8146d789133675ec3d5b74f87a0d8fe2b44f018aa37ac75a44727f1ce79b33809e614cc497f4b2bd6511b52c3ea34c779f9d3b726ca3c0392622ec43acfd2597d5c61141c852c7b24bb2b6600717d7bee3297af584dd26f068d29ea4f5627fd7a483330d2dae04e146312dc34e90e60cdbed71acec97c9b3cca3a76dc8876c8b05498f8133124b40fd40095b6b6f4b0e6c308681362c3fc2596fca70097675125c7abffeedc00478c5ebd77f5a1cfab59ecef954c9965b01dd142a4cdee9d30a20642afe8b14cf18fa169408806b1549a9b39ed31067feb7bba1df926ed303ccfb6d11f12c5aaa24b788788257d062c7c0b79704cfe655ea79cbc18125c65a29383fcc8c511b7064b277955d675593a244c4e83dd4ed31d12b6901ce67e5e02a36291333372270ffa2a3f95bdc3e672207113416aa48316db09968b054dc8f6755f146c17d2c5d4beecbacc7070255b444afd706ed86a1a00ae4e8ce0fce4fad6f10c935dd096b7150a34e4100a240228115082c3ab2b404d405e6b003220f820875f5b8b83bcfe5fdf2402d447eca0bc5ac7725788ae7d3496936361a54843661edcae654d9a6c7976ef64d75aec5873c3f03f2d02f82058266dae2abb091927e764ad6984ce2855cdaca73df66a295242ffbe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h52044262621cde384367e567189148b79c103a84e168a05750416876f01ce0962503933e6b26cde83ae7463f3f01ddfcee0d5cd7189d1c9dc330a612d88c05f0e4e17e8fd6b6f8301dd72b4de3213e5f7be8343d80cba9efe72945e8c32babce4f977f798c8794413318b9cbf1366c5bc4b1fff9d4dbee4f1755d7143bbc43d51d490949a72ba38035bb70fe7496e79d80c2e1061cb7b21aaab73f939c5453ce70e28ba1354d4e71e0bfba18de0a2169fc632bfb2e898f48e77377640e453976606e5683719afde5fe290337f250138cb4e8fe08e025a89e25e01fff84690a1ef2184cf0863120bdb0038825f5552ee62e23fa6bb97cc971596646c85213957f57ae783426809b1d297c20152b6a2652c4e32f67d3ee697e5c94d4cdfd9d41412b2a39bdd583b25941b52176b1c0cb469153358d0b36cb6c0c9a8e9f3dedcfba9cd4e537db212f9881b5ecf0ae9d375d2db7c9016250e29515ea87b6dfa384c7efb49d5ccd7ef7065927ef52d8eca5858ec879df036cdcafb684ee8bea85facaf86d48f80bb2d194abe9cebf7b16a23789d8ac146d14a45d3df900aee1c4952c4d71ae11e3b8c6f297aeb698880df6a4450aafa3900a4ab62dff12e24d54f36127ccd0af6bce4a81bfcb1bd5c2e11dd479453bc3f34390bb5155eef1d54e4eb8cbfcc9df14e266b2a01cd23bde8ec63a759938235f364d5ebfd12dbc27e1363f1d6bfb99d56863928404f98a6d88c96974d8fa5b72536cf524e178eb74d1c65de2a20171274eef2f19b753358dc33aa842157fa5a405571e523f92048d84d85363aeee14ec4c28c040f58fe1e29be3f76566bf92378f36e7b335ad84f79d0e9f8e1855df4715f16bfb0e45f50d08d56f9d17d3fac4f0d840c254e9e081a96e38a4a2dc8f2bba978333852fe61797c0f97b92433ec96ab46e0bc684c012725b9db5a96e7cab88a2ea25667ac4c69597326d60d5acc7f720bced06cc7b3d3e4ed362ff3437690f2a189566a14aca15cbaa85ae4a41d76b9267445167f352dc39be5694f2dd897307208a7cb9e75f07bee6abea16800a061dfb3a492b914a54c1ddf9bf61730c64f32371c2f3b492917d2b122106d75a5bad203d205b80f91480e2f55809ca4559f495f4ab93232af7bc443c4e7c441f4fec2bc6e2928d31a5a52b2e41cfa65671dd5abff5423f4337e659b82f35c54c6601384616486b7f5e83dd219a7504742490dc622d72c8989d6590e529c8ac721d43ae221b1831d7978847b17231114ec5db2e642ccb49900b1589b91113856e1472c32d3c0c48cf88feb83bc22e7556cfe6a95588bddcc891288e1b9c1d1653fe04e3f3066d64fa264119c2dd3ad4bba116d682a05d2976d1a5bcddeacc32ec458c67a7a07ecbc8a02fa8a29008168dbc477974aca1a0b822e3bcefc2ceba2bca7ee0f59d8afa78a81f47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc6ca2dccf130744079b056a454d8dfa49c0e38b54bad29d0025e0fa4b2419ae92332f2d60b17e2b3bb9972deac1691ad4d07e50447acc8555d56805b12d42e255e0d5a04ab1e1026513b7e7d214498dc88e7c87eda30dc61f30cc1cfb13d21a602a08ef261cf0305d3c5bd8c81aabe7cd759e645f05d48b0909065f9c5904a042d14a57d8a194f91aa8760ed67087a4b64f3bcc9779109c58c25f1d230e2e582e2330a40961ff3a6cebcaca5dcb8e19508692d1e4be0940a492b43b0125d9b0c80a9f1e78c50a9cc30b64d45847b5bb237dd099869f7dfea15eefd3386eef07d3987b096c914b56cf5c67316d22daac03264ce3c207f087fffda79b6bbf1c9937cefc9a9e6ad4ecd617185fcd2079a46523d35e2d8a91032ed06cea1c82f0b3fc3aea09a682d6eadd41f38db837e16513bf9cbfc5dfb93c1021a34e04ff4e923fdbbe1f2171cee7157f2908aed13f3f467fb61aff74c9da2e98e3602bba2d5f95454b16a72a144942f24ee6dc83d37eb6ed6a157038c02ff44a619088606304a740d3549e2bb49163e9416dc52fda20c643b4604c80cec15e5120d6afd4ede527ea88e70adb4181c7eb0d84b7b4301a5cb1afb88b584f85ab32d5da28efae3267bee2099b69820a4a68be472a15a1526bd163e2b3c6e0fc0600872f75411c61d3cc69f21a61852619a3d0c6144b3c33cefd6f8144be297792f2a562f40bf1bcdf3cc279e7a32582d24ed7c3c20842dc57ce91c9c14e3d9b30416ec0276b5b9905b986c1edf437d46838434872335388d7888d25aeec079412a83e5c7bbbc1b1c9a57aedc110afcbfa97272037928c7e94550dec2b74be9b60ad632f3f162848335c6b482c7c4969c64bb4ab7e3e87cad7c2f824a1d845275c7813b5231431669ab34d382759023615b591b0ffae9e8776e4a9722de432b23a18e3dbcfcd1c1103c32e405bbbca03ef11e6db0bfa5554e5a358e2ae27e74c6e0713d3ff8574237d42de4336a68a0d1b00ab1c2898e70282123efcb94de75b1f6f1d584bb6976da85bc48ffc0292266be848f7db73ed6cb490e9a2fde03342c33eba833da8d9e7e100639a6d84d1b22b4f4dfd0f2c17be11d4f604bb3726599974fa5745fbf119ee2f7c058b6aeefad9f9bb13cef8f8bdbb3e104e1f36ab0e48b777de6df580bbf500b94cc468556a48d8ba5b34b1782ca423b254e29179ac6bb56bfdf8ba00a520e05ba045a06a9cdde9c63ccf5a62ae7dcaf5d53f63d15227f9459324ce779d8fad8e1216e3350c4e38c22d17800b8c8c6f4faa2a111fe7d987eee664397d235fd92308900e98a7e642526ba4a51dcd1b65fc7f1d9e448d8a8c5752e53247e24fba96a7b112cb29b6b8a99df46dae9857e71bbce573e3c9114a911e6eb4cf5dd6c8c2fd39e1454b8e6d857182d230a164ecdf158b79353d1eee1b02d86867d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h29a467791295fb24afc147fc6de03fbbd5f65cf457ac3441a8de31363dde68d21d50c620d8f0e09f4db424492cd1282b8733501591f5be8c7ac0faa7b1ddcca704acd77ed3e9393d82789b9b35ee36f515568d0c75243cd2cef801d72798652620a5f32652c45c881c81460aaa224177e9e6ab751aad805d1cac8b496e9405fc08de9c74fe9260888be3375361b0b960a7f8416df8d65af59cd0b57dec5dcbfc76628d90e1f40e7a0b128c1ceae53d078681504e8ee2e843fad269738eef278ae354bfc8238eb158ab9302a0132b01772056f433751fd4931954b13ef73b9e1451bbc3aa5c45e1a8dd5100e4b18c0b2260788d4e48c09841fedeb3df09892f8042c398f49a07a3a472ea9a62d7236387100e348a7a495ec0724ab2e948fb4700924cbeb4d105dad0f86d1b66bbc83121af39ac26b93de60a4d7a0311fdf6296dd351e6b67f3b4e2556f82115b7404e4e578773b10b9b30510634762cd44b04c6b5311cb8020d0e4a9978e9aef79ec2afd19edb6b5f58e6e45aaef5b7a78896ff50a9654552ec628de30ca3bd0048a0a1e6345e79cd85d7da2abbd4aac76e32f66ee2fe3536df97a8bdf2f9a958572d26eaab5b0fe7a3f3a4d4e068ca0b3b904f1f7bec5d6f318adc916e358fa3c9745a1ea50ee040dc4e2724a8bf68f61f1bedfb34d0fd13d357a013c0a43a5be70e934f4e271578f326ffd3726b8d955c32bd220c89531d158dbc13fedac74b23a791b7515e403b296313c2a06db184944fb63c3b60022eb380438bd3f4a0b8fbaafdb0b9e4b3316c239e9e28d7b6f5ef66c76fce5cee2ad63fec4403c4a939e39252e7cc76e6de843e40b54ff4b986d60574e89de0f8d822f1926a2026118115266bc389b042992696918de0a1cead782da5cff36fc0eab6f8e3ccba0ce98b6c93a690196f169a6769d45527d4755ca5c1ff24f09bac4217f70b1482dc21cfc68a9030aff5cdb7d48298f165883ceb70615b6fd7aa10f98bb65ea1f6ddbf344daab6ffc919903286d08cb9b7ab6669f7ce18fc5af735d09c3d7eb21f0d8bd431fbf612f2324290e4e122b6fa11d2c851d19fac51135979f1c62dc105667a48924a19767017e0d87c41c4b4a2eb9824c0561cc49d125b21a635f5d5e5d7e3d990a8393924cb839a1047046472d5cf93ea23363c162e8254b5b0aeaf766d6db214764c98d8733f332f5ed28645c6448e7a456fb073b3134ca4e02e81d8ccb835fab34f9a12a954e361e25f6cef885eda1bfdd5b3214dc647500a2cd2658ca6ae0e5cc967cd2ffcfac1faef55310821575a9daf569087dd7badca5cea00ab6c0c9cf9efd2c6e30994e17729a31d3e4870a23cb4e65b06303b13d65f579fc39cd15e1ec2eb96734f36eb789c2a81df8fe6c2aa8d8eebbbed17cbab1738dd6801190c7d3cca5743ccb45c2c80554ae348a8c4f543;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfd70faced7dea8cd5406b588a8db3b7e223e618638b457af40df530160ff54980470978d9ae5ffe5b34591a91a1024c7b4f300bf6f018bd170b5144797c3fa737dd49db57538b90c08d59aa71fe29987e675eb9faa52690a269055ffd4d30791afa1a46588ff4e9dd41ac8f358001d29b1d7da0a6a2598a5dbb16837d28553cadb7bb04c35c3094896c4d657b35d883f4482d16f0ca17c46cbda028697f47b6271f8b5b01e030d54e4191a59cab90b1959341ba86144565db30087f73d18c422cd0d1fe7242ded5906210889d3d2c5a58ef1396c714fafbdbbdbdc4fd161e38d69191749030968d354edbe0f2865e2fe81758e40ed73ae4abecbf2a4db3c6cef2af43d7de2e2dc547058a1e4209b68af4a8d7f7117cad6f7e18242b3d0ecc449708e367fa5b0a353ec5dbd7086591961d5afa8f6fa1a32f143f4c371c7101ef5452d3392078085327f9389c469f18ac59f5f345c7cd283b025af3c9c178bb623167593673e44465542644c3aa3a1b5977ad1fccca7d16ea9384a565ee1a57705132c11fb96849dd77638442d01e8032e68f54f37463bfc8f320c6c24512cb73d3835cbf43306ef9a35194062d869b393cc8d639689e4480323f77b6a5c053a7921142662d6281c2b649cbce9c5d45c37c7f0f307110f15868e65d9121a84b2705eb7ff656311df460414a016f5c96bbf8c32b742e057ee35ed5d3c03b98a59ceffb428af6032de075c4e6630fb773dcb3b0c0f7864d1a1898b039b05bf20d6fc9ad4186a13ccf12f686af88e2daecb4013c1451208557b618a8fe46aa7a10726402d07a72d1055f07577b87a600ae03004d284c7414458a4a44a507d66723c08eefaf5b401ffa01a663d8afa7c7c989d318356c7abf8eb8d1503d41a55a07b8fd5e50deb121b1002f10be470240329f03e3a69c532cf94e72f5efec78d462e35b144fea69411306926e8a2ff0fcd75fdf24c5fe19604fd8d21eca1e903981834d3dbc63c45b7c9f289e141044a9ba413d52a9a2461363c609de6276e29ef9cbdf023f8c39a2c42b7f41f7ab8fdef74472e8a53d16c1921a506ce641d1a53d76f00fc78007fef813ac9912761dd26fcb78a2135b18ab8c4793d54db924131a44e901d0d566e916f4edaa110844eeb6855dc34a6d3f2eb5eac47f88e005ad28ed8d23f617cfa1d767cbc59f035224348804900212d6db28b17fbaef36df50cd717b2266223897d8327ac2fd1480aeea47abd2da2157dbb86701a4017d9b3fb1ffdde9f6879d10495a5bc24faa0630d4a71012772311ac9547f79c70b4a2f968484dd8f2dcf990d30173840bbbce2a73c370ea49062fdf16edca96b93909c96a6f95c8e90ac3f95261635ea716662924701d39ca5cab01f7f4a67ae4586a3f9b9001c5eb46810c174c4d34f9da25e2b3baac2f3d9768f6f47cf2f9d8ad94407e96a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6881330e942f23012b5f4d01c08ddad113b2a3420b8a1eef476163e92e732b45fbe2287e25b28e99b1fdb4eee4a3f927584a90a59bf6536cbd4cbda6be06ec87cb939ef93732c7e083a4c1cca2286e8af31b1cbeabdb0d5105913ff93d5f40ab10c7188ba956541e62f80126f3b4c343992b48a2bca028a8155ac72cb102853d6a93fc8fbaf24aea93f958606bde05bbe12015926366f6ea486b421eb39b6239d8ba02af01e26307c8a7c8c32a87b75685fffb11006210de7b1f16903e7b96c56e453a26d94fc4f7c13a28b8cf34d34d8b3a0e32f9fa97b1de2a9df94f724bbf4a35ecd7422eb63c6857e7c87c41f07428ec13ee2b66617276b56a864f57929ec4823979ded6702f4249bcde645c32820f2f2fecf4c769cffc48d9078b3876e2e8f95e3748055cbaa06ef68c6014cf91b650f64f8a9638476b53ed8d6aa9d807ec3734419e24d1ee6d1665d94fe3d8393092f3bcd930b30d5bd71aa42436792270300d5ccc2f41fdb706e54a6d3842e613afa233ab82a50d4a035f2ee8a719e96bef22804974007d6cc1040474209f0e3698e57452f3eb965829d43b0cd4c3ce59d9c814ccf9782afab95942ea4f4dea645007926b20a757fcf9bbf6f11f8b7d19787cfd20372846cbb4b00f1c1b6a8512ae95e9df51a083b5a2d0b791f3d77ff461b654e12252c1f5557218bd3ac826c4c18ee7532bbf1954684d4e4963adf27c4ccbf8c40fb8d0f186896ca47ae70595cc78101c98a6e45835c3fe612fb745ba2a45f4c6dfe2204859667deff97d262d99b6c3b1a16ac2d8dd586f9787c0ac65482cde1e12c00239ecffb966a420c1d1851a801922dd90f05ca2d0c2bd3139ed376b2abd485686897c5aa8ef9e91b4297915d32b043ae7a1b57647e0323f5299352bdcef9412fef7f8defd0be2d018faf7d3140daebf414d082745fb4360c1c88edee53811a9b1f3576cdf731ba65de033eff7626fd2079053c57a0c009c4d1064ceabf7f874e9bbdcd903a1159ceb1c58cbc8582ef6b717180fd70f7423ed67cf3469fd17a7af81fee247269bdf58100ed486b46ae5cc5b1cbaad38937b9c7e436d93ae12ffca888c6f27e7d4c454596b258d4f9a48dd82145df916eaa9823f25592f9704c9a3556a74ea5c192fcd1ecc055f2b84a68a2b14ebfca7383deae137a0edba6979acf0ff46631f24bd5fa0a928c938b8699a2cde2d91769765ef2bee7886609026686428f21f0e8c060936a5b60d41773bca8bde78afa6d9dd8a707704799ea4cdfbe650ac8e397c061efba6bfd37e429146b4ea72c9c40e1a256c807ac7be300ea08833f631199a3be8b386e0b50a3211a87b9070ba07a1aebc534e01a78d7d251f9c50cff134002dbc0d9247e923729a8cb0a58b881e002b8d67925d5f7f2b5af25ad28582d7f21ea3bc081b85145bfa4ee9a5e6088e26041f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h500b3ad9658dd286f54161c68728f0d2822c6f03c92c76310abc21542d1d7a98aa31a05f950f11b28d3ec51b7c0891209fcf6c5e5568bc6a3a58fd01f843562e88c303045a9f33e3729e3d0d6d49d7ca0f4c704e011abfb4bfaed52fb09a8b7d29e0a092472884b22883162d98c282247ee719f52610245bf50e02e8189a343b523b09ea160709441e9560fe4c20587892de39cc5963c7b13efd0661a5315f3abfda2e7bf2a6f07fcf68f80b9b381ae7ec3d93052c72456d7976149788f7ddc0391b03d2e215a67390d5530acd4c04654c678921b6aaf0193347cffef5d5679dbd4c81e654c342120b9d9d4af1804341702c3623e6439a2754bebf87149fabcc8e3e37c1727d4b733afd40320dda046c08aa257e59635c27bf2ca8fec626e71ed9cb4f18e4e30a64882390de7e3c9a3ef5a446c0e84339b3dc2bc9e05cc3841fdd426870a5bbf8b56fc858f11b52e539201d162b57de0fdbeec8cd9041ff1d7236087d858d4233d5190fb89a43be0f83b8d41c280a0e827db5aeb056aabee8956922618e087aec5d006d6fcb4ce08040a68cf86a0aeb12959fff4bc13f9d0f6a90378f13ea35e23d3a1a402377f36ec6bff93db85cffe5a8df62d0ead7f33af90d049ec2c425657c49994562d384c73b2ed25971226647ff51656e06de1a7a15487d76e924f5f1474a59bb5b393f7c21251dbcbf9b259b62bd489d9ba88340e01b753f5e612c4d6aeecfe7b166549d5222fa5b9fee38adb8de7ea0abb878ddcf11fce2a6f33db268604d81f95e6136491c5e70ae32596dc5ac02bcfcffbe97493924a33c31608506fcaa6cc23867d213b6b96a278021f5dfaf4fde333475bf058043edfca8c64dcbb0a5c6ff791aa1c38e7df323902396a30c9d5e7f09170dc7cb4aeca68756e5f9c09da69a20855cd580463cc88565dc739a037143698adddb562482b8f336e1626db2003388c6ade1183c643a291130bb0a0c14d167a294a07f498c9a32d3d7563ec03b4aeda9bc9cc2fbeb3d18dfe003583f2db5cdbd936f1b9c8517c27607ebc39c5131d15917ab53af62bcf984f397fa6d561c04221a79cae7b2ea64cb5a9ecf265542be90be7246072c26882ebe3bc1d905f8a24a36afa92cdabbff39df73c90ae0086f4e48684a87287fcde9d9c25570a0cbc859cd7f0c3c81111fb5bd1b2acc95d732eb4eaa85f30da7064922b6601ba7485da00f5f7d01bbc05aa91bb2781b21811c048b6cc1759bc7ec34949600110dca320e66e520371409ab9f036e9d6c3d542343e84dd4e90cbba52ae2c194eec1b2e87000388939ca8cd5d435c64daa7a9479e42ac1959eeff06b2765dcbe1b35029d7b8cbefc5e9588117ddc7cbb6cccce6a076fd5ffb42383c46272ae77a0768c2f123d3929ff5b0257ea79baeaa91ec9af6b7418c466125809605d1b89973b0710ca7b3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h934a065222dd4e4d97bfd4289ab6bcb7c10ed58cabb27446b7712a902dc0967ad0ca3f8985621887e9ff5a88e5092162b69484742ddda2a2c3afe019bc47111656330f8a7e71ed5846ba6c4b8465d1f111ca7cfcdbf925a3a90d53a47ef1b3d7b8c2ddac49fc47d58f70e37c01c7062b7c63b5e318d66e0c2bf3c59e3f347d3827c465abc2e885dfabf3714e18b0ba460df2a08056dc563a64f0e71561a88414b076f62c7394492b0d63ee054bdf232ad359aa32ded789a4e6a9cfd3e8f89ba0ef3a425d02ade606b572050fd7e6bbd20e339e19b95ff1113eb1ff13bb79f5874750188fbc16d72be27b07de009b41975f24b448f86ed62efe70b21d039450ef0d256c3ef01e5dfb91526d1e77e03bd73c02ee7a078d941037e4512eef54d4f447a8b35f6d3b3d7311a8d980a6525e5a78b1397615d751bca999d19fddb6e4a1d7a94c12307dcc5e0b9b2a7ccbacf986dc76549cb0ca9232303de24a2928c44c39d3f872ca2a9abd897e94a22b2c7ef0a1a96b3a07aa74c6197ce34d48a9d6adef103a8cb5e46c56bbb19be7b9c60a0dcd25bdf3ffa3cdc30bb3b8e9887bc75295f1303f994cb319bce6bb7b42d4f3084e6b2636ab7777e3dc756034aef95dd430b43a924d61e30b43223097a131effcd91a44c5cce16264be4a96e16edf13b929cb3bedd3812f91039c12e5440b83f9ac83a17c2ccf79feff9424a348be216042b33151f6fa74c7ab9cac4ae8b4f7428bba47faf0a19fd3fe4066b3a0abcdd69e99c0cf44d08c023d57a3dd0e4d359ed280c3c9c747b22a8e286fe9da256c3e2aa780b9e42427d9ff471ab5329a558475f96f7fd2c5faa76437ab9046f5203ec6c677627c694232cca9138a752ff1858640b99a42d764cf4585e0eab8036faffab8797e288c25254fcec1a104c2b705b500493a8fcd697dd5981f24f03991a91e4c1245d9f218f7fc2607f729ce64971d00e7281648779854f905cee1f9a777b09df0bb2c9861a5c97fdd22f817c22cfb79c5a2d14e74a9ad47a83ba4aa10767643952b7ad02fa11046a8e63f8edaae386849422c2b48f76edb00371e4595cf8d91416e2a456786751eb0751e3997803edb50271aa411426b4ebc19a333706a7e902f85d2f8be4934df06fbfdfdc438c4f7198b1978d58dfafd06592bc87fa2c0915d74c3e8ca193f76d242438c46b2b4e026ee543af243e8937ef2587771e188d0fc3171d7a87725a629746f01f5200519fb851bc163554807f8d98b53bafb285055b2a3218cefd60a87c9b86b5a3ca0d61e54c2aeb92c1608ef3ca15a7d4bf9cdf7f55179a04c47654c263dac214d0164e9661534ab96a8fa19ec0b03fce24918bf07a73ea020c219d30a793d09c2faadf451d685f9cf386e6801e0d875ada61156eadd8f0c1b45d2a2ff4c95154ae787c39ef565b7b506d5020e7a34f0f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfc564552ff2ad6c7f2cb8afdd9de4e93cfc36c9113692bfd2fc9f6acbd2130c72ea664d8e1d74d0e80ccf62daff1fdfd153eff39dbb17b5e34da833e0987c0fcdae1a877044f0ba61472891102e70f3cc38d53db8a71a4f9c71b029fb312983af01d76f24935a95e2839176b3a2f2d5d6d8d43c5b54a553aa4c91a53aad1ce9b6ad72f1bcdb54ac0620a809e931f519751ae020846aa081dcb03d7febd0ef51885b2feb005269b990a15a31169e0f912e728a645665ae77a69aacba729423dcad76b99aa83a2ffe521bb97a1f7e35c9f5280d3180aba68db1932b7e304714e9a64b06f99a23ed5f42f328eabee6fa133c92c0f77653213d6f3aeb610af6c57add38b3aa612faa77d2c1e6b162ecf04d3fac480a03dbcb5ec0268b199233bf001742edb05da3ef60fbaa7604d929a72064ac077bb56cc240f9e2c47efc6208c87e5f70a55b4a31680e7bcd582c3d01b5b797526341412edd8dad2d7cd1961fc2c1c5daf06490ea8b5a4017d9617637cdc8ef15323fae91715f4e9e21904a2c83b173f4090cf8adf8f049bb2e181f6f1016e61a7b40019f995e4d6ebc16924bed9941af53788230ea8d13632cc49d061b41e54eba9a2cff035d290322a850e85067858f0c8f7df01fdef3da1b498cdc278a0cfc7bb485a259e0d78d51f897456eac7ae775a815cf321489a45644474a0d08c6d1fd908938fdc1dde3063016bf4b7b6ad426a377885e0dc9dc124c84390b4bbf88563d8e8873c916fdeb2d14a63e6ee3ae397b48077664e4f2001d30dbc03741a6c0f656a10886074248adac2a7031247aee6f3a7fa2139a402ed553d5b06136ef80bf9d73f9824fab01469b08ea96a116d7cac3bd96730655f3dd9301d0cd5774aca1f51d6150bd842322f22b6cbcf209c4c57b0600aed0acc42ca1e5619093e5374afcbaa7327bd140c8e301566b4d35534d3805a1f65cdf3293e16d687c959d793118e31ea42d12119fc769519814759aae9664f9a5b2a475b7afc03546bbc370d303491ac5b4d75ad30022061e50a191792e16533d5e2a159c5b3b75df0ea00edebee7f0c9ef66593972e538ec8ab4932f512d76b0759f702b35dc6222022dcad8d238ff08c9dbbb05bc6e1e09705cdbd5a97191e4d99d442f712d734f8bab74e4aa76b1e03d41044408fe05064974033ae821b2bd5b086eb102d762b50efb4305469c06075c526da1180d31e314f730c3e7dfc0f2b92ed78bd1490f8b46321a39929a043b4430b553aef7f143d9f1cf8dd644df5f26fefde77634e5d82f023e1123e814bd389974e484b0f4003bcc54a18d0234e8e6ed17f154e1411f6bd1572f0a05d7698aa7fd044320bc7d89efe337a94301a558aa44a14aed8b8e17cae87c199390ba13ffbcbfa8cca023de4679d87ef9448c0e7c517476c1db5ad38438ef88edba7185297a73ec74ccd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he4dfd6c70d943fb608743fdd0496be8778ec2096b8d84aeb4175a42adf4c21ea16ae66746a42339b5abcbf1044965e10dc9775a99149a21acaa93d810dfe85cdeb83ff68cda9cdc852d1ec4cab348e8d72d2a264510b816c2489083fcd0bf3ec99daac444dd5e16ec0bcdb6f1b4db0aa66d14057a6eb94182761c9d959dd29c7033bfef5c78057f51e392d3dbe0314e6c1e5f64f4b9c1393beaef182972bc9f16bd92e63816f2a5463bbefd0ddb1983ee8f452a18d7c8cdb67b540c5910562710d52fcad4a7da51fb87da430619e1ca34389a0f12196147b68c9269d82e1b516c22b7c61ad3ed871964d376f15110247c4d215d08735e41d5004fa94940d349a5ee16368f15ffd7f2bff66115de3c5812caa0edcc481b4cca413208c1ca53d47fc56827c3f34a0db2d6d08335db5211c68d7b632e1a644484e9a7179cc1d4eef1c136475e12c94acff58f188552aceba18c8b19fee87bb776ec5a4830ee5154a5e00c1d21910ff09195ebeb86cfdf4bcd19de627642f44d2f7816a8e82e9efeba069a06beb5d450d37a308185475987ff4c6e983095fd197f4733133d5ae50c9d98caf2892a130aad65e9e62ef10917343b87f4260f94536d57dc90749e21138aaf2e80a645df3d452b01c5bcbce4935bfa4e00ac9037498742ed3c00cfd9ab9cd0ab79e122825513dd93027cadb4b13bca6fbca98671c35ff3db14a9cc0074b27d02cd7337fb0ca0c859dd583a7ff9ab41d378dddb6d6729cad3d9c3a33fbd1df981b99e7a4a8ed9a46a8a0ff03d438a74e3ba8b2b844a7eadcbbd757fbe90be0038b448154dc4a4df2b68e0913044e8f0ca366a936370152fe0c8c31fcf3856aae0a2dbabea1df7f5f6e28bc604fcf291f39b31a487447618f118876810f4662c10225d9d18c48621e5a58a816229c531ce6fddf8ca3f511127141e8bd776ccd43a905a65e822eab4617baa644d267c841b63b9472a213849524149ff46376e4c972d90ec5db9eac9c55ab4090f8cedcf38cedc08fe68dad884ebe4da24df03e43fb80f28e721e19e15dc95f9c609d0d0bd7495cb6f9c5558a8b4e543656bf6ee9ed766b3eb06002e0b12f58273536ca87cc88616ddc4ad2f49ae272f4f11090500f523a0a20d03213611688d1578016706e2b48588e4ac91518612cac2938d0a1ade45f8f435a987176aad126b31414937dfdb71dd3506b479c821b5fd518313adec55f5adc51b6deeaf3c928193610c1a22b6a45753366f85b04b900caf7ea2e6c829f0bd16f48fd016fd6b3394387aedeeca2cf638f02a1a9955a38e4cae00bac794b7efc393f312074235443edfa06e2baba1802bec50976311a41b5e455cf9aba7568c7ccab87a93453caac1562bf6f67e8c07fe67bc8770c99be150ad0c4eb092fb01586b4439a3494c6223e2d2868498dfb9289dfbedf2b33de560f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h38ff68a923d789f164cd792b0406610479e7e21a85dbed0dfa6a2d74242e4f9a7ca6596347a3124e84d60d739773b27594cdf8657536f67b9cd4f19baf57a4db4990401400ff91677e75087ced28beb408582da17dc0d5bcd559ef1e0ec13839ac1160a688ef0641c67e35a049544c10f0d83006a1d567a6ff9ca72f54d3b9e4dd15a8e7694edb87beb860b5f3478cd5f44a5bc58b1ae3e7fdfce8a87d8908fe22993b538d51f367aca18b43f2151e309ea0c17d46d0c1f39f1570cf619f74e02fd95e724d449543b9d613a078e4b422c9f135d052aa6ad260e6187bfc8f175187fa037438061127c97b12af892312a42bea08f66a6018faf65a7044cb9b7c1a3616c03fc652536aefac7e7dddbbfb201ba4e2cc5089bc4e9063cdad67f6cb75aa5f24a7b4842b7b93fc34a5674081f898e18c0e6023fd390664f3b51903aceee768f63f9d7117ef60cf1704654b281a5c6cd671d0bb9f63f517aada708f7e767bb477fa7782abe4f6203de9d72eaff5b601fc13d94df4e4501bb3eb7e9a5804997eef45acdf8325e2e7b9780a493fc796bee1131e9ee602498dd5235cbdfc6ed8295f24ebac92a56ec31aba7201516549d6f39e3ba6552930e4b19381b72eba52df7197a1da1570187e19fc484097d9c98e64a49853bed9476fb38504b304aeb66dfe290e7843e70b1b9a25419e88d8eb0d9cd1bd91dc69ea781bbecf5f72a28a03f9931addb52929284ab48959979ff834aff623fdc386ba940b0a6155e59c1167c90a5145eb607b715470839abd15260c6fd9a7e4485830d1962049d1efeedd7ef4de6ff9124599159c5d7e965723ebe008cbe643a1f5fddb8bd5426442bebe8225708e907ef505a9665f843bb5630a4c4c72699cf7a74422ca11a11e3e18525dbd3b838e8d39e606bd7c5695849da8a992866883f9547e9cfbab454120eeaa34caad89b65d2c7f5f987a8b3cf56758a1a65a7d0f48a900e639b7cdc9a8c60260635f2af864b1534f0aa89dfefad33a96d00dd17ca99ff2b2bc9da1f3b8a43d103af050c8b44929c272f73bff3e46101b433966638dbc9bd60d639c5185b15bd9d68278e0079293ac5e306a5f58e59dfa73c286e47e0f6256154430dad2535dffefebf3f76732fa68b22348a9bf804ddede7981159cc334fa8f4bb853d516860198c355f60dc6dac480db7558e2e56eff5c425d31dfa86d2f874bf04d36bbb619326e646765f2bcc18a8b7064b83fd4a61b9c300c3bd16dcee4e5902ed48a87db93bc05f6d5faa9e9db0da891a2368a5749bd0223e47985ba0db05d9b0ea40f730355d1f1beb8ab398627e91c3e2888f183769c6c7357d6f4003368bd8354625bcd01460232bcf8dcc3885828d06c53f596ee2549324ec490ce8bf1c73dc5659521d36a6c53aa41b5862146b09a08e8414bb8145d5b8fa0c75d8ba02b2db8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he58ccd612138178215c8b6bec11d1f6614138a8df1bee0876281a25baced05c2ff770c466f8654a74b7b7538683bab81a400cb2b3c4f1f20015c2dc1125a7edb1323e12330e232fc8ae6c3d037144d9afd90e87a1895d1e7764a7a9ad9a3154b04c406035b13b454b82e438600765e70a67ceb6f007d33586a57f71944540d428e6f9029992379d914fa5844f219c35979c93c023a141fc8aa24e73da9e086b82705510f83e365f61c5b6c710bf795e20f18829dda503f09f981ec02cce58ebde13f27f467fe01c5f1e1eb02e2cd7da830b66087bbb64d0d18ed183fe0a7c8004187ffa50a9395da350617d58feb42dc5a9e44c11eac46f45271805f12932ed8923c2141e70fa788d6872317c738e1769d34fe1d629117fa1e1646a131cc42f8320c01331dd713a00b5b0b2cb000291b90eaa8e3e92d4415a0f2ca6ba9634e184adb0cfc35f8f73388fece00fa16392b3c6335acf4a1b94847480e427f7c7dcf7a0df1190c5d65ba8a6ea22a982562d3e8babd31a5bb85f17285cff6cbaec82b5f2bcd63271f337bedeb04aa7bc35fc7ea9c1dbd1989ad2bf0a29417d33dcf0fc985a68095e520b7667a1805295744dbcf429230fb6741e230de415ccff57c2c9a5edeb6003c2dce5ff358f2bc09ca5bf7bed00aa5583b20a68e327861efeaf04a169f639549dd0be454ff0cc4127f6f0c84b7ac719010adf09b852d5afbfd798e6f3e4a2f897b06edb0cc98525cc3fc143f80745058bf40f92c4b3c4e78d66caf81fbed9b1baf2602caca6c3a770a38099c2b221dc9d4359ce84c842c7bc3d74c84cc2a2ea661649fc639d7b241638356dbd064c28f49a9381b28fb5f0dafaeab87e0392fb339acbe85f07e9d0995af7d9f1a9f8f182b2dc60ff5ab26fee766e2fb05720ad636c0451f74f944e5fae51b465ac8661424ea21507ae8cccf2aab5bc01614cb44ce5568551a5f9cb7803d27f3cf30517196c06389c5a59a95c303750e47f10003c3600f95c38b342ada47e1342426353c8033c93696062356b77a7ef293f8953ac02bb99b1df4bb3e486af7027d6c3390c5799d1e82a889a513ba7ea37c44724b99c65b1ae35d79826b250bd5f45b5f74ed94ca490217e6b8daf51c7326db3ccc9352082e58dce3051d98dda05b0449e8c67d55ef793d49c984f443372085969e8454b5d2b573578564734c8940f96781865704b14c9895b46c5e858468342626720d06ba09a471ce0154518e0063097beebf94deffbb11ad90cbed6748532f2098dd33e004f5d6f59c5f6a87e6713163f876fb7d3e27bd35ffc7d363bf01553e685905d3152efdd5d1c866434730834d703d824114466830e45bd89727eececb8af22ab8a76a4855ba710741b2cd46c42d2207fbc8e89eab4cfb39fb110a2d7933bb9bfd11e100834ba7f830c78b3f96ccccdcb42e609a6fa2fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hab39fe261af932aa0cf0dd479f94c38699c7dbfa0297360972e9674ddc738a64a9ab453e4efbbe972dad09c8216ca309ba85fdd944cc10d4108684c52f4c85ecdb50d57f8184e430ec1f7de29f9ff6ed2b477f76b52901ab31b86e471177e3e2f0e7e05788817244e79295742e74529c49d9b4c62ba68b3506176fcc7d06fd2092254511537c1cf92e33f6101c29850578e64f933cbe4ae20122839d8dca5eca9ad2e1aaa91f5e4ce9f3fe8aa8e3603156cdec003b10d9745601fb4a95c258f3dbccceaf71d0738096348a781180d0532efa5c6429d13f80da334bee25754f1544c1edb1ae55d50242aebdda15eccd3a380400b6d09fc317acbf4bc2e7c49baf9080dcb1a8db145d1323c01ba019b61fed888699d3b0ddd519143cf1e0e213093d6d65ae9cc7c667d5a3efafe0e4535ea1a2cb21040da05467d5f88087bbf0b0d838d3958991a466c52fccbc3c307011d5429ecdaafd37279e85a21a75d1d09b685ad83d2e40bea08f5fe5846b3cf08fb57ab1e312616456763e6f5f91108fb6e303642a088ea04e74a449ba2b592a05f6cd47985f27e83ed0a19577b82ddcfbdfda7c87f7841ab6389ec3795f5158d9232a9157057f68221b6d8efc1c696ccbe1963f69abf04b563b5a10264bfa0ef6d59308652c1975dfc683c21bdce8d66e3c57a82b08452f16a81c708af7363828c76c3141f69718e74c0d7e58015b31045a9e6b05d5ed627f343cc4010c590a3388fb22e3c7d2e0518adf157de993de3b0d55fcc1cd3ed3ade9028b04eeb3b8ef69176d040f54ced1add2bfb07442d8a1d069935d0635d0e5c7ee85f4554acdfd631c95d73b3aa88ecaf3de1f345c314566d2cc15768e5c7c9e40e36a6233334d9210ae2a314cda8e5ccf0d417f2739f089a96eb5eea701900a1cc52b361020d5c3f070b34a349e9a4704c735684579c76d818ba5660b9c086b02cea1b48b23e1ad828d8fc057a328396efe8fbe988e4034a4191758ddaa0df00785b755ef5b50a6cba81e5627b80ec095b9b0372633c2aec2078d56bb7ada86a3cf3278762d71e36e3849623a328e4d4413212af9a2d18852218069e4a846669caebb26bf560ac29589db879eaabfa38c63ad52df4cb72f94e1799be3779d30d70f115367cbb52f84e763d8ca40ce2d8008a3abb49db2337e19fe65c502c49d68bc111a5e119573f3b2ead19a873656d60bf39b8be169d5f788f4a9c654abc6a4c89f16e385615eb7395a19a320165786bfe9d1c1f5308a050f81cba80c3ebe417c61092604d700e60e0e5cf3b5b7605c06c2057e80d3b0f79b96adebaac517eee798deb5b289527a29933ca9c3ae48a0cf59c27104b90a8e36ad56e95dfa910dfd2e46b31003e9f857c71b359f7727e805466a825f87f1ffae62971001718a70853c11076d40fa06cc53dd8f332d555173120784b80f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha5869e0b141bc7fd5924e06a2bc9ee787cf9b418fc65e249e9bc602496bef68aba4f7276d914986f797a069aef8a645fbc3730a457023af003840393a9e7ed4b7ae1459847bc509e9c7373b57bc2cdb25616a21b323f795d6ad62b1980661dc21adb9239fe69b01bba9cf3da5fe0762916f6141393cb9f7dc779fb4d013bf30d26063023c33c74215efbcf426c54d31b42bf4801320a7422c91b4a1994ccde98a8d64580cebaf64b375154ff7933b4aef7b5d16ff271b4223e295ccd0a75ff9a1efd98e50d65619ef710e56847a63e0e944bb936850adbe572ef712b59771c2ba977aa72888f41d7e2d0e624957a78a9357ef0e0eb9aec29554511a1141826c407feac8edc8543a2cb1c4465db448aa5dc5a9cdf9f86adfa1e0d76f01c388bb47f776b99725b98de959e136692a72be7e088244cb6f711947b4b0434586b09cd29aedca9db41e9ef9cde5ada051e88247582e07627589839feb0c7905d4b0e7ba269774a987d3fdf2adc42f5b736da0e56a2324ac879f58585968e018f0e686e9dba3ea0ec7f2e2af4a3fc6b3a5ee8485334dce6d88e9cf160a58c6010012b2ea4c4cb3d6c628529b8b7bd598c15e802347811f4d0dd638eed1e61102ee58b4fd65020d8d7489dd4db636cb074b366a0c2f578fd6c7d17ae7858d8cca84d518b1d85dd3e3ad1f7c4b252ce86999f2f87b22ebfe9249084c1fbc53a73a704baf49062b4626bd56910dcbeb2f05ee99f86e53aee9b625a911b3f034b420d59d97721fa0333979c2b4d637a3b7316f1e9603f3e47548bf6952f2009cf055b13687650151b265c675127212e5104ae271091b45bec84b3222d764f7ddbb4502abde6932bf7362203af960578c938e5f252566d3eb5ffa11d7b597e3f1098a7d03fcb644da54f027f839454209ef52d53076983920c92ec4c5ba13049d33142033e20164473ebbd98da89a0d883ee6ddb57f9330aa0d44ba6bb08e19558c7fd9c9db6c92ea842f5dc0ae1fcf1f33f4a777c16507b318cab1ce345f68054e6c3fa5f3fbb0e6f17a695bb8549bd2d1562ad6755a0573c23939fd14632728472243d15d732e5cc59a613b92806045ddd958047ee0903c6a459da037299bcde31a3864f646a9510dbf1d746272bf0f976cc0b8cd1a1da20a5a1c0d452a36d13bbb756183b9d8da0cadd06be67836a2277435a42985a3818788979634f871d4e7d4da3efd5bd1670e56992d2e356703628a1c92da864b93d2c0e3bd436259929fc07c5792984d09f0c6ecc1cec3be78de77a29b557b741d7b162260f02bf8b89ee9261d7eb96e11ed95cc3437fd7ed181e90ea06ba95893e5509a4ea4ef3db281d7ad1231738a0d85707be592f4e2df074e062a119d0f4b721d08579e8b867ab0aa366a08c61cd9def677e10e83329717673347c995ff67319a727e6129bda08a44f3e9fd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1072d3a6f666ede290d89130e11f53240bc0d8e30256a00658fc081737541ec26d88cf00a0f2008eb340012664baecd01a518f5b9be81e74cf0f5d8908daaad38cfc13b3473bd2b3e5eb41d88c6cad7d905876482c1aa2430c58c36c29f3adf1ad2025c07247f4d0a9eceeea30b9e1b1cf36aee39a367157f628f2068cf3f32ba78ce40f3cd97c13ef69aa5f6c18f8117e07dca2bd5693a91411ac24d156aea9d6794552f8d816cc667d2b38b367554c7723ad125276a0794a24727ff391d0894de5dbcefc6bc28328cf6b5e9e3c72a00af863733d5bddbac64d734d29e18b40c692ba42bb3a1aa3341d5004eae7d3a7c2cdfd84508394fdd072057af8a4d6c26e3355a3eb31273bdc55344872a66879de8972ff60fe1692bc5ebd4b4d4fe2027c5adad6234166f75539700ff1c9be71b9f7ff836048a80e73f9f9835ef953cf5b802bd96acdaf7cb7a27aa33f735edc012a80cb84219a11d819defea309827010c79091d7d72240a8da678a695fa677a77e5261596c9534c3d08fc6c02483f60d0be87a2cc1a27c599739def467d22b6b753cfb136ceb837f2940d3983d03335a9c5c97a59ea9d9cf0c1807d561b3a6247ccc76b8c61cbf4bf398d296180b0d5b76c241d1e39545d03c145486045ea8e9a8297fcbbd6bae9b9c6ecac7b13fc02dba06cf43ca24f6549c8bd8814700937ef8d3d7071a7f0c44b172a72c5d8f85bc51c6b2c9a2809bb45c94b6b05a18afa2d33b5a20ca35222f2ac37b42e9e7d3a2f5797ca93f0176ecbf33a43bf88ea61b48fbe21c7a644726024a9d41d829442ab1a280b649709637b63d966ee1aae9ba0ea210e1dcfc607e3a4618949c2361a97f9c094f9e53f6aaf865482939a05e7a451b267754829b69ccfc56987776f2aa2505705a1ccef3b3676a2a1bffc5d2c3d34a0e868650f2c68f0d4f9ad728e6e60523b60bb3a50517202b6509ccfa1f692da7d283111812f156800880c4a133ca6898a236217f23b5147072cc4f82fa86b90f00476b3ee86bb80beede144887c4f023295f6c9db7d1266e825b7ba3d6db77364814f1e90fbf9d0503e369d419fcb8646b0b5b3021a0b881377c049dba37da4a0c886b09f3b78c2391493a6a053816dceaa0cf1f6abf9e5eba75e56d099f70e684f7e8e46b122a02472c8df0027736b99a4271cad43f126c6b85f42d6b5480257b0eaa13cd42fb2e1ccf7159138d783d367a8029ec4ce667700786c4add19e27c9871090195a45b3a72271b2f97b860443b20a8d790a0f116072bff9c0de26ff19caff7a42cba9d7667b0f9153677d0c78080ec0ed9a3481badd90691e459a6e3926d728c6f71710d4a007017672a284e67b7a8c647e2da65f1f20fdbf3fa16e542fcb82c3e52e36d96a147d20be8891c831030524b5f3b45b7a8615af13b1bb2512fdd037a0486422d582879b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had11ce85828b2c1d694cca9abd0200e0bda2fc7fa027b531d1867867b69772e627bca639ec9538297fc1a2806842734e82c078dbc9e86780ff97b73b4938d8de0d64e10ef072d9710448931455de3ef7fa81ce888ffb85054da30367ce92fb0b8dca5e4661bdfa4b60363745b0f960a97ef7c045e2cae3a7c652b98d4d485ef9ec82471efbab7f95edf7dfc3b9737a328ef7ee3bfdeeefe0afe22a74a82c5a157887808c182758a6b9db91833186c79cbd0495a6be7e7238b08dc95ec8501dec22a32c03c5e85597b63d731515ab557cbf179b83c4d3230ab11a9370d51b7119a3e1c10c11ca8c9e0cb474bf31067783cbe64eb78f0ce725e1dc29e581b5e95439ece421e382b3793356c7e7bfc2261d484ee4ee94cc1f8e9d93a367272fadb4cb6e702cd7cd217d66c116f9ba0f3f7fd76e1747ab2b117fec4efab275f165de4f42bf7650a533b656d252c7cc205c074547a05b45e5fb10bc9cfa01ab15bf71d30e880cc3be40d927f55886e2fc388fb964f9b4614b649525f535b3928f212e38b3839ac3f40e5762329d264f7e9ed06951744ec79331261f6366cb9d70b6e23ae5cbb33c943f96c50c0ee8d2efc6191c331e9b72174536231bb71bfe7bd8bd1320aa045d68a4da4c4a5063d523206650bab7527409b2622d50180b8202c0f99b76527379f0a0837dc0fe15ddaed747f367e5be16d435866c50f459c57efe467cb9848b298b120632b5aa88f7f02507332fc56b1faeca62a49201107babad9be4cdbbacc797bbf9a34462b64691865ab9f5919febe89eb640a32bca43cd9f2ee0c86733312402265faaac5dcecd5517ad45d7ed1df4acd7d5796f2204808cd9b70df8bfb248dab83e6ca6d0fd066b8b9b5d96866553704e5f365c1d6082390b1d1f05eaebae51aefef3af3351383c4dfa112c8a454daad4344d95036c6172ca7e41e915b4ac1da8634bf62ea500b7b3d9f9475cf99920301a1806475eef0c5e1d48a72a2a4992803da061bf0fbc0c5f775ea07d55dbf1fad9fd9ae590b9e054805f5eacd6b7e2fe76ea1a313580a6ee047472daf6442aaa20290b84f8cb789b8bd48a0669ea715258d370edfe18e82824b3e522d2cf8727cf6aeb2dd171f7f4fe62b8a129c185ab3dce3230b3856b8b186bac034a7c1f014d3927c94dc8052aba38eb34d831cf4ce138f3e92e81013b65f3b39df1e6a3ec4fa6eb0e3a851a50126ce3ed25e61e4a515da2606482f5394045aaddcc789c74363efa21471bde5f6beed6621177f9bf608966c5cedb5336563cae164905f5e8854bf3a542a5746145ec3e9e186e01bc369076e510f379bdc93ce6d8c3a4664a337e8c0280a15a0d5a04bc74f676c564a13feaa22ca0129fb7dcee08cd7a70efe524ea38aec0b55345afd35fb566df1708b663123adf207616609b44dfc05e7b13efe2a6b0860ece;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9af4847a9f2f45e706e54b94a2fe03f9a87bb9cf6032b81b87272dcf81682165e32146a8ab3dc845022d0cc3423f4d0b3ded31f00ab23abcec627977d8865c8bd42b636cf6ecbf377bbb072ec05c321a05805106173b0b0ed87e08daa77e0b5721480cedd3a72e4f526caa7d0a2c154d895f8be74c011540095a96ab32581e139525838f2b74327c6480aacfa694f729b163eedaed772a5ae7d458764271870150b9f09c812b3b3995c5bdf7eac5e4548a394de969b9d13cc2401680953bc9d4eb785afcbd148564316383c40d3ad27c049975e3a6e8455ad5421f224b469001e4db2b395698c8d0eb375187cdc56ae29f92b5853ee64ab06daead643e9c470012dad5e8e0b3c50136a310855689d0b50844ecb161d01af8e925938daf888d4b970672307b8088f77e67d5bac0d3b38b78b49ac181840ad34130ff3b8d7d5a076d4891f8789161bf62e42f92a1e5a9b78162a4a366eed8fb66b1b22ba41c0eacfc0b1570a5558b691ecb3be9eb020dfb060c5cf6a4c014c5e44982dc8b4c0ef6dba8587a1256d40e215f17d09d298522cdb692fd63a4bce661fedf7e7233693b0f168cf34c1d11478b183e5f6e1bb05cf27c145d7ffe4cff7145ff975c8951589d76c35cc909cdbad6676300b480ccaaed0de13453883c3fe7816ef63bfb7a896e626ea75274ca57882c11c97674f5765fec6826d1206689d0de03269924cc0764d433c183cc16cf3d348efff8b66102305d3b2d434411047bd5e1861914e8785ee14ead035a6831d7f7b9d501962d2f136643c6e1553f17c90e5f217cbf9f6bfd672f4c31aad1cb19d71770804d0314bc7de47178d68e2120c531d418f57715870d92d9cde234816ef8820896597442138dcca840f816002ebeb638d25dfefa2cac9c1192319d9287d0bac648291f6c9139d37b5ae5714b202227b4be6fce5aea72f0bcfa7d7af78ce3f87e4ca4b15a2ced25f44d0b5bc575d8dbb000ceaadda73f403c207649308b60f1bb97eebc79ef9c410fcd7f63722832ea3e72de58d5d9ab91ce2158d901df8e55dc6435ded3ab8472c2f2b59c66383ac50cfbf826fb4e71865da3b0f472ff96bdfd163b8aa6b08593b2ca60c922dd00cef9ffb2916a1f7a7ef3214cdcc0e39fbd17edc4e06520ba2886ce1cc52866e708452e8a4c60c78269dcc1634e3d5c3037fe4687f45e752cd3d0a39641ee54bc22f6a86292852a562c2217d9ba0ecea36d088b2255fa927694e30ec2c859b9efeb4107d083d5baf0fa7dd1184fd6daa4ec017f96887206b23c679138f5323f7d42ffaed781a4ac9bd6c90877cd0c8a902f258690053d00c89ed7e817af7817654b8a03527ce0927b157c9a041df8f7491742401d72b81e7856bdc23dffcaf39c6f31e459290b3bc72f2a29e82402de6399c03792fa9636fedb4af592f333069807a697a4991e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h829305fe707b309cc375ac6937a6a29fffd9bf153cefcc84056e6e3512c82e12410882a749c3fcea3b5820f1339ec8e9723de7ce75f1c90b731c9aa642740a2f1e161c9bdc06b3b51d0d7ca71d5683956748e2a8d5fc513497738dd8b2a8b344b80c39139c24cecc5de31723e3c613c6f91e58a446043453432ad865214b294f137968953e86772c6abca62848941492254c658423a8d783e005fd94205de3e11ded75a0fbb019e4b70c857b4e30d558457c27bfe295bc252295b77471c8181fd745f526b26037f64665586e12613bd0ca4216e20eefc5340a8e25e0f49e141a305587f5a5911027ec633abce5f7ba811fc256a23844f814c079090976d6adf4251227891a2509a56d382a9bbf86fe7b5c34cb58f0c51b9cfcc930df32e289201b66da7db8ef21d88b02271b3b43e6d6f54d8ba562256fa724eec57493d371eca4dd57d13d8e35dafb2398ce04ed9187ddc0d278e98bb23cc5f83529f22c5c07355220655bd4eae1f28d79338d5898143465ed713cdd43d7b4caad6ecc1282fb0aa3a8926f3ab183985fbb421d431302087fec70677121b431727cf74032642e8ede3594bb887715e0e5678ba6b16dac999e1283c1b53facd6ec6d42257224dc539bfed9d23e2a42f594576c9162f7071e15cdd6a02ae7032f71c28d3ebbf350a014a1d4304678a0805de541130894dea3c451a7bf47b2dbd4195880145e4a36a3dc0fa8600003b708aea0a1b129836517d131b44a4375af192e295b68db0ed4839a4bbbc3c821ff41051c09158a1616eececcf674f723240a64aa71563185b6bcc6985c3f63e1c7757b3dae6e3a43836cee21d06a7ba95c713e0e1a6296784c39084868739631c8acee6ba62a7ec53ae6124b44632faa6740ba36a537047e70e524ffcc87c6605681404edb769d6c25bb3161bc0786c278d5f228423cdf94cf331b3c1c6a0455450dc36eb94da6337b393be4cfd23ed9e42526a934b38dff48d557903ce0e1b3b1275d811165b49353a946a2f5cb70adb0e86067cfff321734b1030058ee2f55d30453fa7317f1d94a3ede96bcbbadc32ba3eef227a8b5bf764e136a9ea49779299f47ca2fc29cb693c8c3823e0eb0255b7fdc9db95e328038346a9af9dd8cc4cdbd91b4eb5320890568ea22ce863b711f3fd5bf19045a5791229e38825cbfa9d4acbc52792d5df12eadb12e5dc1bf5d78393c5971feb9e37b200266b5c1d36a7b95465be531cc3b63abf772967515142ffdaa1a7c6c67d1f8a5f4c9ef0bab5bf931cc5a576663800bb9908285766d3e9234bdf0193f530ccb7df7a68788f1885efc21c553c27c761d8e5e23066268b1466f6a888bbada5f5bbe0847dd9b74cc099ebd57b37cb63d13cbfdc9837e73d59655946c96403c282204ad9c701eebe9e9a85db7ad081495f67937a1b8484e4816172e327f69405100;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he399f3b556816d0ec39b4f8565e66e67e61912ab5ec61489b780c68b13a9739c53a73831ef2de11d7de86820b4f50938e38563aa93e2b8f8a57d7e6b2e3e2fa3e84fe4b8cb208ca7cf5643f09b17029452d759e59c06c267ffbec4f06b3ec7af428b3b0dad06d3d29a038015f97efd58ecfad78ac0d6e6bdedf9046b9bb360e39184fefa24f28c2211db1f1c4725076ff02ae167f02c62c5ef82677e919588ed5e912493a44d15b4ade5917cfb3c2fd8775489ab05a96dda9354911be3f6bf3d87972a2cf76729768386419ba3e9ed36d3b519893c0eb38e814dc704f9bfee663efd2dc19506f9d9a532e7519ac765345d5c7cee2c19f39318d985fabe1db13fe547ac7dacb4d0e65fd919fdebc1f7089f02bc17863698c757cf38683e2ffe93adeafacd2189bcddf5a00f82fa6ae78d48d95def8825b3e2352dc96dd2191dc577a9914d1d3e52c7059cc2680c9ef0cc20e47249a6bd639a36934e6ea7ff77214486f2da554fef199eaadac9e82d5d3c2c2f828ef7da6970e9f1eca802ce7fe56d83bf9d871ddd64a023b6322df1b6fa2d9e4316794598d97622e45d97ff2f133b404a988cbb81363e51321bf54cf2d96c54ccba8c2bdc4e8addf9668441b6d116c40ad69d0eb5493ea43cf5c4acf7dea6e2a11bc8a6e300a08ed083d9620b1d13e22825cc2ddb2a6eecdaf0d46c65ec44bccdeeb8bc52cda78cccc7a1d55678fc807a506e6379aaeb11ca3168c5f5d60a8dc226df01e1f14ae9509f92cb1384c14a37e9f77088802af865210c2f4655dd4d972e9aa541bb6acb2a56a175a762507f194a3a1e73d62d78246d9188309ed9dd6acca9bd6e871efad77093f2146e8073adab937314425e033c1c0caef37e4e040c7e711757e8575f71e561bccc1a9f321ac3476173b66a29363da9ea5090adeab6d911bc70cb87f5b64075ff2c34df940a1ec5a5957d425ae9f16df01421e3324af2ab111e2ded3c3f987d935e5161dd5516c432fa211f59bf4ac9e95cf3946200e7ff0e4b3afa09789fa3df4b9c249f887b6b1c3c21d61fe20f1d85ee0a183d2b14de4fb55bd302cacf6eb7ac38351fadbfc1a825887e8a929345d50021d689c5446c6ffdb333a24bb5d86d5dc60bbec404b167d772c25cd3afbc09b701069a091c9b2113112f819ee5b27d4f1f9ebb0b51de4fff69adf70c572ad26d02b46f98aa77c8a2dccac9f97c8f911fbe20ec7945a220d478be5f137eb5699b8e43d1bd90ab97043c895543d75fac1eb1039b43279e2098659d349d386f18d59db3bd163d309bb5d63d48ebe461275a800e7313e7f5704578d8664fa7285d01937c81f33c304253c001b24fed7c7d03f017b52f411812bfc7c5514d4be695bea95dc6530759d17365d44695a7ce67a0a2f29ea39232f89d20f8a8658126f9f7cf2051f25001695b9b08c13de70c78fb60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5925b20020049090229496834267f0e1f9ad78a38da2a0f82fd3e94a2ded5f255b8b81d8cf5881166253baeb07810f09af9fb0556cce0e591a8bc5abd8daa8876029ebc92a691e1bf56973d09c81eac54f39646eb1884d8647a36b44ca6d0748ac0242d0f6a787a442160db7cbca578b56c77304555cfd4cc5d9ae9f0447735d5ae107de5d51d9770e6dec2bb0140dcb5c49fbffeba0e1e6f4391c901ab8d9cd2c05d53a3d60c27ed07e47605e3ea01af32d1429966bf1f189e3d24144167343dac7638ba0a21ffce6690152af85ac85f1337b09b3e4c61c6a323c2b7717cba7bf5cacce2148884aa194a0647038b32234d064c3e9e09ad33c9bc1340d62a60fc9262756ab9484740fbc7f97e837ce37fff0e6e676ff919d13b3aa0d48ea9686347ea1acb27346a0587baa1ca93101b98b4ae1793eabd950e5bf2434676df478bc5ac88cd3067c2ad10c72039d4eb69a859f6f363d44816e9c9e4b431419d550720fdc2501dfc61cbe4fb7b9e67b077322c94e60a809edf488437dd327e106005e70b59ff0321082f74159cda27f75ced6c10edf20b1455640fdd5bd6dd2945a6db0facd92a19ba00205613bef044579ed98a6cebc8ac1722ad40cd3bb903ad0aec3e1c3de8e9343cc4db453eb03243c00808ba34297b92016716e6e201a69355f841b4634930c4180534dde906805a8fae325dd68b8ac955fddb0cb3b0923200f9f697a60f098527dd5e3fb760e9ae4d308583482bc974d49d64aa28c7a21b8019ad86c476f6b218351c22d250b4c6bbed9e2c7cfa6d33ced8a233ce98dff9ae09fd2700c116662b954d75e5954965678354ec5e928e0267fae2ee7c58930b07afea066c9a1bf68ad0e2ccc21a2b256c8ccb87ca6652c3414dc110bd6d78a5a7845845f0596972ef86985d5c8e6ad8803f88a4f57756aaf433227ee99ede5f8fa2bc171d7060cbc309c400931dced2e9169bb2b9246b779af7555cd3e34965277d4b9a095a6aaaad5a00a4da58d41182cc407a584eab35b425ac6abb8d3b4c41ff4d0943a436579ee8f2e5d973f15450bec51b260b960644567ab66cab835fd935a55b0d22348ec6bbc428bff7638252d58a31ff9f122da571e12940b44dffd08e3a0508569e1a443daa46b0f190506cfa9edb1da77d1ce742bcdb99af23131085582a9a2ba8e8994c4451aa1856e391fd5a0033b92ae37047ee555021845797c21ed3714f2685c607b3eaf3e914cc9a4e008b4d7485ab47536d04f2b8120efe7121aab5064e36d1e7c62113b42a870924c8c3ea308156db14d14f4738e9144ee62ad4c0a8ffc72bc89aa957d348fb38959d53779c17ff0931aefce16977d46ff0a48ca54229b0fed6fccc1c8604fde6f06d8032553dd473d32a4c636c9ef409598e00e3744c92a6d1a71fca0e69fb6282136c47c83b0e33a882b35423a1ffd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc3acf55f81d2f394a759479891c66a117e325717b89460adadf1fb6e6471dbd1de7e4d4ce50245ca74cb4abab783670ecd0526d1196f652aa17da5c4286ff09822f5b424575d0bfd206e775f40352d0aa951f3f50ad49dbcca8760596832c5300e6f44feff0cc64e8f4c57eb8ba4fabdcd8040379c94c2e93bb84dfb982184f8c44303aab0a03b1f57bfc7766162c74d94b6b20268e4761404619718bfe349a70aaa75f932a0c53d0f6f55ad11b60272efef85a1123fca7014c323fb582364aa19cc723a528e24d037dac591cfe4376b6db6dcab451eb8326e4f57ed460e3e1a277667cbef1ec7fde217c35eb5cababc6bfb28662f1d84f6285067d7bea60812034c08f9f8312037589872169647b8b53c6bb87f35036bcf45ba74d17ff7bef07657cb9eedb8e341f3af661c6ab66726e4d7bf61bdb69eacb93634946b93e53542c49cce13193ff32e42aee28f62eca3169fceb016c259d72879aecb6eab9c295bfceab5cbabefa548bf7d5a1158ba5d7160776627e27903a9ee21d6e655d41d26457a86371a39e874c4afb665ab075031f8cadb2c094487a59bcb09e217726c8d07867f12d1f29d3df27fc02ee436e48a84955e81ecafb35d00d35323aea08e7512aab871963cfd579a20bec12b71ce6fb463e40785c60458123e01ecde4aaaf8a1352fb22a6207c4c66565074b323aab16ed7a92262dde6d58093441d519345d26cf53507a36076ce3c9955c5be672b618b9ad332cba6b74382d31ec5d95e460164a83965c765e7e898d780c1c52241d92a560f9aee0efedd3e41fa2afc645088c9b7eb310045053d1d0164a762a8a954f2771e95cc0028193dfc7822beafa85fd2a5f1594eebbd6425234332b611fe89f0bc31303d6e24b6e42033ee0536229147bf8ea0b85ae88950d1ce234e2339926a2fb6ae329b52acbac92fc724f5e3baac4b71c80e09994cd16552a9b4d37253fdc536d57fe57e247947b9152f0c091ae40446a759fd3478093bc4bcd47c6b5b5ab1dee3b37df7f4faad44a213df6df315568670c5986967ed95e6e69c6b8ce7d938a738b689882b778c8e2cfd02d067141a51295dd8ff676d36b11108f112dc9176781917e20259ca69e2340dcfa1d8d05eb51ba4883374bdc6fabfb02e1a21e2fcb30b78e15401d80f3f5f83b96367c9c15e79c3a066db2c92ae1f632bc11e966b6771166336cfe4d97bd2dcd349702c56764fd98cc30c0b2e5a3a4780e64620b585b95d412ccd05f3732667823407137e04edac787c4b5c56e36c87e67b1663043389c677335d64fa57e72e83e9f0d2fa282cf42dfebe4287cfd210550a1cb48c82095d6bdb4bdbd1b074a38f9d73b4593c735c00f561acebe8fedc8ff78094bff0c98921330d25474b8df7b68d1e2a1ff62e6a57bc2d1e47382f691e0c718f1e08d807f8be50c58db454e36b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc8f6a263032595cc7768b7e0a97d3aa581f324f1e0e572360541b99f2881395360b936ab16ce30b898b5f938c5094cb41d9effab3d0a4c96571e0d7186fc9d7a0fc66ac491572af86200d81c311b76b8319011fa93bcc968bcb7b46129fe2c8bba513fe943b89c2e5df4aa3e59076ad9eedf85ab1eeb5417194c506b0a25f9f48be98680d2acd1235696c9dfaf44356045aabed3ada311bb3f54c7cafc3340a95f1598990c6b79aec4fa6e65ef14b16446efdc1b517800f4a038c60ff413cc60806646276f33878816bd20f36b6eb1acf0f036c3c9ff1de494974a3076d642b0e2729dbee089520a104b82c146cfb1d48ddc67cdad05ec01cac01692cd16af5047f61d6d0f59df1ece4708cd51a668d02e74b985a46a3eceb5d825744a6f425ec70f563bde500f42236cb38ca0c2a894a828ffed126db19b18e50eb6815f4701813726df426934c868b88f5c2e2e63615fcca3d152afc51a8a2f6f9fbd927dffb75e259faccd8f9dfff9624a383bbf504cec453a769b0fb822ebad42f2eff4ddab3dcce9359ef740609adb9d0724c86d88fea7957b8d5f6c3d6d04109190ff2b17f8f65e8d52837ec220a3a35644a61a2dc72e0b231ab96125165eb01d76217a33b5886705b6f83a58e4401df52ebba3d73a322cca6539a97236deff1751eaaf1f701855ec6525a712cac015e3b8b5bd0a7901a0b5d7d82563b07a1ca49a3f509933f6018f55cc78a12dfaedb87a9ab009314b9a4df20e1d9eb5a9652a2e78241ac92282a7607fcbf22f6d7d4223e007b4a2ab9eb38df2ae73368d431893105c0c77cc3bf72d4e79db37397e4f4e50ac4a2f0da3124de84f931fbc1a29327db4cca721500991c10d2132132c341a6eb7e171ad23e26958bbfdfa0b9bb30f44a74ffa600aea6b4c82766add3c1ecff20b607c810143d6e14f325f0c9d49982b5489aab6290e66ce01f6e00bea4163d5bc1c74989e1247163931d6027835716b349f9088559329995959a183fe577192e66a3de156917ef4b70252452543704f2cac7da38d8e17b71e956934b82535cc1e8a0ab1870723720161ee2db9be998e0025798a9622e900f116735572193115e21be3938ca209e363723baffee06b4511aa421e5d617a33fd0ac7cd3ecf24257a0ddd8a516a4d5f428156203ac4dd7fa6ec9fd040caeaea534499a1965e7f3ca541961f64fb7297e37366890809e3b4a009f0d6b081f433ceeeb981c294633e3cd646376d33615c5837ae935309bdc6b67c9c0d8d391e87a674c0fb488a75c2c8427da82bbba6133fee1b0a2e490a83422d0249951eb99027c255cda2a4c656a246449dfffdffe2623eb95ab19602a05724b24c83652058bb2a329761b64078d29bbe018619c7d3c923a77f0065db9724d564bab2f13d43dcb354bcd49f97eb0594107197ef8b059513882a0a727edbf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5217bc1f3ff728f2b6102d843192d4aab6d5f2cea0551079639ee88f140067cb0ee7c8d6e806208ddfa558178495d835a9083cd9bdbdd95321c3cb5bbc323df62a6dcf753ec5e4e68a7483f8b92aada0f6fb301d0c0136d233e6c0846d4c3825efc8d210168fdb1b473e0be59a603a3185c5585da44ef244b64c0e9d6aa459540d43695eecb1bd7f46e751cb7007b63ea9c9afce16a3b7e7f64dfc5ebd4d01004cb175d8cb425436d1f925628d65df380b1397bfd6b0486dddb9408419d25901861ee7be7557478255ba178039496171df7c9a7c222cb54ce09795d6f37feefd7a5f714edfd887b4efb7dcbeb0678a3c4905c08294e63ade11047bcba19975a1dcf45c133c738ff260c9efcad378138dab8fa7a4d124279830e814583e1a6ccd6b959e2c40fc25aa1a9a98ce7f83cc771eb496f64cfad9592818682b552b8e53a83811903804fc79840c958ab906428db9bd1e6172b0ba0bd06a4481a39e18d5ee281087c220b6f3587074b4e58a090ae34726324636fd8cc7a48d4211afac756b0bd9d09d58eaecfac813cbd27a9366e41105b65f5a934b2e883f8ce9136c6646f62f7da4f6bb6d3345c997704fd8314d2143379ad85ec785166636112006332d5f8d6ec58af1f91af2eed9311c386c1b5f5ae61a26a8d7f3101416ca2668084ebf8ba2fd4ea9831214ca58858df98b4a1ff115010dc83f7c2d9242ea6339a5ba77f9760d8a26f50af2442597e7668865ba178f96885fed4ae333f5d7cd08bee4237385265626b29043b6465dc02539b5eb341b9ed5a7cec96e85e2b1efa990ea093a860e5c13ac3c781ea4584c62e258d47d0d1dd9b8a538c041c0ff05a4c74c65a38d2c6fa231f591dc236f152b875ef5947782fc5880ba13edb74d7d8316223717ba9239f0deb6d8f9d8b859fc0d664984bca487f9206a6a1780cffe4317fad76030df72a2bcd950dabc20e9f720eccd48a5da414e9b9de471f4b261879606f8010678efb47170cb418762011c639b1096112760c895efab585adcbcc2c9e5a07646d4c365e6757a8ac795cbfcd2cccd1b48ae865c0658ba1c18a51d717f342c68301a0c1b214827fee3aba1b45918fbede8387304e48f9dc983c0d8272a16e3fd5897d2c123907c505d1b7c702b26a9db50d58d8b1948b7b7ba2362b8d470d79b2b8d4f876044c3b29b4588d9825650375e17f20e5884a845f9fc3662c05d8afb291364eb11dba68e7b288e3986f8137c01a57669eafacac04c8393a1a67e321d48d4095823e613bb01f95b87df82c971072772330fc287dfe380e9f62a77a1d2dfbb0e709639f2c28fdbdb340188e1450d4afc2375a90f9cd726da68bb5e9e5f417d61ee1a34d40699afad95e475a62e0f50f4a3e350859be44e4aa0a765413918e00287aa86bbd3b34e3c59d400c729ed9cd00d89779f4a1f9239526b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd11293293b2c30b670615570f1e9e34e0597b13f07a13ecd5cb1ab27c4c281afe76d60756196b9c382f314b606e3115e0dfba0b09d2b7909f8f361ad113830b22625c901dfa7c458ff226c62fe1be76b67b685615dec6f2e9f0e91b5c2279418b2f10321057005635eddd5e31106af45027afbafa7adbd19066992ff957b943614571033a3087dbe27652fc01729934a1a15d952f938a18103d2b9e0f3241897aa1a6f915360fa055b380cba844d68383c46604874410abb8162eddb05ba8f98ffd395bf0a336c8ba6eee9e3b61e08fe867fd5bd5b05c77cb0ff9cbe7fefc88940e41a0e23b15d55f140e8d82f3a013f1959bdbb2a72f34db88e9eb20d7b6afa77ea09d0ccc155773514b8e7bf832d969b0f4fb2645beba55924af88845910fcfc67b8bb0b68dc547effe2b815be450b418d3f66d874973dfb5ba7883e8177f19f285cd5c828bc809b03849a8bb513ac4291fc997dbcd11782d9e8a6582e39391fc65b164333fce13644cf5f3cdf530002042f50271d7bf719356f9dff44213ee03bf28d7deb0da8ace5f868ef188fa02dac63c066952b9b8a910bb6f76c67539ed9a79f4adb8abe434736a7fea08041247c94cb99481602125f4179f44d253349c0be6a9c1e806a6b74db2ef93c103bdcf9b304fee1e0ee965c9b881d35ed01b6e7671c23b851bada76039be8d7d374064dc922e288a918c76e7400fa92d3b1d15270279b502384aa4517d0d335a68bc4fa9589ffc769807205aec4da255b695756ca3ae3676906b644db0b5f0f9438688be19fb98a3894ee8a3e809310b54247dc59851ef1ae959d09a584e997ecef7119bc72d21a108caf6dea4be5841b4c29d392e6ce23baee8efc0d8ac98eca2fa9cde4715dd46e0dc60a6ca30e69e57601be0b901b58c404deca188851f521101b10ab1a5ccda46868b1c0a67e3cb057fcf4c62440d2c0373a8c5e2d499fbc66eb537893cb21c143c81ec92b2b7180ab54b0de985e1f56a96af983d32fe434d4d4cf613742cc4c38464f06f37debb548575d3a4552b5780ff8a72965abc171148029a4deac78fe44941bb415c92e7e42dbb2b91b139df429ed7ff131ea374b3e1813e0c84d5369d711849d4ae6a551fb2d4fff042df827695c09b65e3936edcda8aab3ff60a8db79f88e3c7b8a796127e0416b78c9bb852d5aa769a4815c8a50b071b8ad398df0a837048a414931a5cf00f31fe02d4bac18816b0ca0ec9720e9670e094031d5a8efa972b24508f476cd366ad2432120d930d5ea5b2b639e217d6265807d4b3f5633cad3dc6dc52fd9695a6de50157bfc783adbecf560eb89059089ab3957d55548e009391a9b2bf05b3e7bd9104bd006b2fa0b9a418a67edf8848478c51f812371aca13f3d236f5efa7bf01bd073739df6c67687bf317dd59270b36ede3e04d348d40cde6ebebf49b90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h51fa1b82520a1e290c36bda95f3662f3b75630256f4e1dd067fcf07837e279d8cf6dc5bb6179a033f2e19c81a79137f9ed0bdb8f0887d96c030eb85137d768cff92f3240fb406494446e448301e3b1277e5461152ddd44d86f085045dde9e0ec34025525392f19e6891f04a941c839c5651854e4a7fbe63beceab53320dc17f3a37f9d4a07451c30cb3fcde974aca30ccfcbab24ff8aeb20e4e893e520e2d0022f51b4f71932981baa85d0257204bf88132ec74f250e6995d2e77c90188d44f70d84945d69619aa5193862a62a209086cc267b57eca53946e9b1d83c843fa22721a9d737d4f5dc34732de78e887518ed6fef4f67d14e1e06ee5d95bc6e0392b73e986033f57d54907b4e55033978bdcdac4f57a27ef6d879857afef84aedb14c25a102fa27ab4850cbc68b928e558f60b7ee7d93e61c6db4fc23c4da859c32d4d85c845c2313f06f3b788fa901c85adb8b8bf4321c361e8afca5234fe49c39bc9f589f6bc258031cf0af1c018a1eca6f1b2504ba3a8a98eeeb71288cec465de26023bb5e20159d78eb88dfdc5042b5e544775605f767406f93a1ff3aa530d627682a5e96d79653282eba8e44e45bded3797c55ac4b8c127bf4c616bc5e3fcc0e62da423e5c88b1d56fb067f0208b237111df12b7bfaec0db8fe9e39988f5fec3201bc36157f93ba13adb1b26ada2d3031a3d7535fe6b5bccfda4bc181596c96d29e3b14cde95a8c095481c3fc5391e8328ce5e49f0aadf3d447c6ff155c1cd4b0f680bc31076f81fbbec87f5407f75225e84651a922a35adb79890114155839fed3be2a3d0c018f157d433fd66535230059f0735a58106dbb09424b4729698d6611617648eae94b5ae1d1da91cc0b00c6c2bfc88c955b5ce87adc931168cb5f3bb734f40c81bae23251865dbb6f49c19b7505361104f483ff24df40809b23ce572f0876504ba963039ebefb40bccbe4646fcb583dea4a2f972dcdd4e5873793bd707738f89de317b5d47644695d5823cbccf809f5d1dad89e89a5b0928d9e2e0298821d50d506f591acd8872dc2efb13da8ac718d650352f9afe4a5e420c847341ba7231d322576e5ed5b549fc8e41ba4e1038c8cfc35ea8cf882f66b2ed14f46a0af7ccc5e76ca510aad375d1825d0a46ad890533f4fae35256d69289b7b26258ded288154decbdf930e27811c7a93062081efbff7c3362f84a7d39da16c40811d968420c480df3e1a26c36e3308b195adec8b41b772aa5747b9b4b44088154a0be2a9d29dcb02f79f5642f2307d20c93d2a46ff7656bc95b258cab104f7d6e5f0389f84fbd1df4405c33263b0e6f458f87bb656bd742854575e206d838a9ab3005702b0eca6f54c583145a9809067e6e64f73980c299765a97c186c4741896018fbd89497f84204c010eef6f0d4f01e9cfcc38e97d261e8dfd7b87f67fdb27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heacdc5fc9d585df84897902faf22c9b7305219d954d1db61b490c3b03b4077edfed8adf8312bf766d0c4048f1c184124524ec4dd294d8293d29455ec58eacbfe0a8f77d74cc96700455f149775f929aebf044b307aafa2c3932d372c058959131de400456954c19defe02dc5e4a0dc07de8b6cfd9da93a9d696dd870b113a665c1ac5d125e9e2412421c0ce750d5d3621fd7ed5f85018db3c7e570ce6a94944b2e430e1056fdb1077a7cf016fe05959ee9928ec3ee70c4b6f18606d93ead0ce5e2f454aa42c11d2583b8ce3a77671539b2ca32d174d0bc35f922170b2f1e788af3c4452054faa75c7da978c1eca747aca509b58cdf73d9c7bb7820d28b7f97a73066f34bfb1be989154c8e536afaf9938d085661d0b68d11aaf63be54c48e2585092f511d43c5fdc0edfe7fd051d063cc2f046d72eb8614b88a4a0486b7a2c45fcb2520e75b7f1847c6da24487cd7cde55062388ad8ff3df1a63635e8a4e570eaa6fa679f8cf1331bcd191527a052fa5a8c96640f70a7be66173e703a182924f56830b02dc17abde878b5ea4d11736163e5d4b15996b70151857a1bdd4bb7aeb4ea402aa45a41eea164dab6d89ac010354de9c8026f394cd1b7285fa6b5c6351670edde5e4ac025cb2c88fe7c64fb69c3c8e6d4bdb46615eaef14417517f9b3eb04d772e5b63f39e885e7e09b69a376a13940c343b0ad636c5103ebe58eb5dc7dbadc2b79f8749b59e4855c723f21611adfa5bdc480d9ef523c406408dfff21a1ebcc1e5967908122ca9f2914e55d9e76deea329a580db3469bf227d4b573e9c4ae6a93858da712876b2ea2a9f566ef5a4ce167c9967179673208a61602ab154ddf0d07a033bfd1dfa3d222ccf9956c6e1789f2d6911773a8a727943a802b3802b1ce97ffc3bc4a56138e6aaafaa386459751907ad5027212e0d8e3370a66eb836a509d8582b121299ef5fd51e1413583ed2c8938f92419278ba35d7485637e18018dba1d1ffbd0ec039b052e85d4153ba6ef3a6e9623e5ef9eeda93899861326680654c4f5b9d4b13e5d73c8df1c49d7c09fc4be5d1a9fe88acd1b81a21c64758fd5db5ee072e7edc68f4820b51f536a8e73b7e577e9322c027f6730f98e64e8617fad1e2c91579a4c140b6e3000a263d43fbf3ab36e68457858c3b16a84f5d70c01b9ad8414dbd3925ee57f1a49221a38499ecd973fb7e80a15ec0bdf33955e88271b5ed54eabebf4845d244984bf0c7fee3f59f74334f98f1639f574f26ac8ea6bde2a43b2f485e3bdc2fa5a02722ca981c8efd85c5a2707a266c085b59604189307041031fbd7a1fdcdae52e45d4babf0d7271662a5171f6c62c577ab236929c42af54a73095470fcc13cff83468a5b0b5efe4b98fa31aafa2e13875dc1e788712f67d0d1f4be7a5826ce3cbfecca29620d339f90dd7cd95234f9c4a02cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hada42a070f0357005e09762ac9d9830472b20ea5cf79902daf6eedeb0e37153902e88fa3449e059ba5388a2da859a567b79c3b9563794d653c394be90e51124b2aad320a06ea0cc6be3042a044454b524d7832bf6f19372c562ebea37305515d15d82a0dae6e519d87a2604e1c7097bdf1b5087ec3518f5eb61ac75d1c85874572436ab03dc02f9b29dbf12f598f2cb274812c6b249af7492da7dc070f5f1c650e89a800de72edcdeb133f56e54cf1411256ae3247baa46d5cf69c70a1fb88aba8b94e49249a75936fb22f4ffb547484eb12110ad31e3ea846f78ad9724171d48ae84302e562c10b9b10780460d5d38d7c20d76dae2caba51323cd92de3ba79c9e2ce36924a4f3ef349de7a7c1cdc5865825e0b44f99cccf77bd50ad576deae893220de8c52abc7d6d89d865560f0f187eb4119540427ee1b91e8344f77964b69d149c00ef2bfb473570c4f82a8be43751358968f395fbac6c539783eb23006d2725f0ba97cfdb85d30f270e3b389fb3378e2540b4b3b4f29540eac6f12c4f6e143633e3f0e84ca0e95d6e5b99a7778eefb75bc1474300aeb60af8ac5ef86ab8eccceae0798caab4b93cd1dfada9609764ef6acb015bf1c16e76393446bd662dcc4c78dc89c7d2840e15ce93c98c6e7ac9d311aa7efcf8825f96dc4d05555bbb15e1bc2ea4631319efdf23115c32c2446d9621865f30989f06363ae5412892f805436f8b3f2a3bac6c135feb0a60b055dd5d5876b239e8d908847e9647c1e5e254da6944fcae35c328bb7657a35b126da1d68a53a32d07ce598818b9febe72afe3a86f2d04928047c04ba5f310a6f7d4d62cf597d607623c6acd37dc0a2590d083d4db5a16e53cb41a313b5e52f42b101f013e4344f36afe7be916fa0c58c70cef5ca8a45c12950ff2ab34c145a5b6cb5c81bf54ff44d2960a278a0fa37da83cf3360f7f69c03e15c78e38fbfd394351223535cda569c7856407dd3e93591ad3e5548082b330d34e7a9693e71ba59c8df38de0890faa7c0478039a5c731e97c7a8981a27c60bdb0a1343e30cbf9622061a3f3f482d6ce830305d33ed979e3ac171b137030257c3b989137403d6a478ff4eea909437847707458eca2ff5c7a0a75eb48ae518807f4358363402692df1a91249b585f591591d8dad542e6964e719e163374a6ef295db6eadec0a3f9ca2bab10a6f690455a766991ede0ac3347610197c6782cb0bc7c177e02dab197dcfa7a90a3898d087edfaf773876e6d22c58d77983b03d7841193333094e264dcdad3b8798181a854ee61a5decf58b01724da911f47e06567b3f5f1c58a28c91cfa83502edccfdaf4050f8057bf2a9ccc10ea47749973e148cc3cf4a7c445003337ded25dce5479536aca66336d065b671fc141704899fb5b6212636053bb3d8e1c8497deb2533c3d1e569abc57d89e105629;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he0fac186d63e4016e8d4caa7491a92591eb81d78dc7cf3055bb1a54617bed96e6e56b6319835bc3fd53b24a5d075b66f4df5216672d36c8e66ca5fcc914767dccf6adf45b49dc2a668e67ac5267969164f4c0c6f0e700ee2b433201adf48e4d50422129d8e0bc766034f7fdaaf876355f28637df9499b64a46f8e969ab1a36af98fc2bbd895fdee57c1c7e2384889f5194494064a130f1f22fd9e87f5dbdb8fd31fdb37284c9ed5759f1d468df67852824e532bedfb275eb3179ce6fc02a120f04785244f98b1c0eeaeb379b2a0ceefc3c76c46904920aca0d6b912f3992a74f328aa33786fdca8f0452080f6f88cf599f834b37d10eb439a56c405544483baabec7f8532debad5eb11f72f6715203614171aa83e26ef2079eb460ad1c7d0bd9f5fcee27c93bb028ea87e4acb0d19ec13fd446b62d8fc65da6ce332dd3291cd21a02dae6d45e424faf53f1bd729506c60f114f9f297962d6ff00dd098ac0238040bdc598583a220be8733de4af0fc60e04250e76cfafa3f3014a310ad84aeb0cbcac93cf1359494ee69922e9d481815ce3ae813fd1823edc944d9e5e044e60ab62ca75a4d275a97231d5a119a923f17a097b4a2167cf759b343faea132b370ed3bbee9826a1ccb4ace4f4ac93f34b761f48f23171f3b45b247282a55401e242c51003f6596cbb5765e74cf0598332b5bb3f9ec9fea11488617c1ddd85d1aa37275f1873d976df81d659a52be101d267dde73c82593f1c3126b45ad4906812ebfd269110c621691dd7fbda5de1d60b02d56f8b713f5fb033700c37029aadc16b0c95ee39ceb06e64d62035c319b58f99340de0825105cec2729e3f216a1ff315d721537a16b0cf45f3d96e3435cfa55fb5476fe6a7d3c609e6952d12c28955afff03d363c143b84e4e3532aa17e82f520ea5a961f1af8d4c61fced06812b0b4f8ccc323370f159e6919d561c23c91874bbb06a8124dac5e499852de393522bc9c7421f2d3e34211f9ca782ba22db7b66e1849153fe4ab5d24870b035926f7d6240f41fa8fe1d39ad5f4651ca5ed5e0fee577dbcc88fd5ea8c889296774f1873eb1b9acef96f8b51142a55349aafa9c90f866ffa8f090d6deee15bec1f7afa9abe06b91e01ffd2056e3307b8a8a265eca7c050a46396d7a040dc147d3c7e2cf129e427672f2ef075b4d9b5de2dae490734793011c112775c6134f0be8f5f531750dee354c97213992c3613971d9a67e5b5b1a60c9af40bd99529b8894f321e5940ad7caa648965bfb61fd41b11f2a2a2a193f18c3f5f8e6f7b2f6ce057c8b14881b525cdb90e6f1276d969c3efcf93210ef53f58687fa164bad3c3a315ba226af9f12367fda13c5257bc3ca9e31f68ba3f2e6b9f663a2496cbd992b9c2a88f42fc075100c0ed6120785355d7037e73f7f2dfc7d80d2a11e47ffaa905bbad1602b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h77697698645709e069ec2027deabc004096ab3960a9f7faf11d8019883a58d9470104586cbad656f7de2c6c9d06c0b8ac38e61de0e5bbf07ce28ebc96ffd1de301317cabf5f22e3d78889a5ee0134423ddda6bfe5d9d6ff0ab5bfc236344e360baa5af9fe196fab4d95e365fbe0d769b6b311bdfc3161235fbc7a2765d9de084359e255e85d30cab1cf7c21148f9889cb2e9a712a63b24120a136ae9fba6db1739cd2a0eb8db4bb87e00d520499db5e16ebae6abe18daf0b450b0659cd414a93968dc12b255ed71ef5c112ed1c7563bbd8fbef15ce672fc1280d11129ea694a2b54eae23643f40dfc1c2345a66e035a3825843f296e9924c01d4dea8b09aa95e8207984a78b7aca467b1913f0e99d23b06206dc7d2a24e2b9d2ec1179d9eb7ed21b939c27ebe794bba0990444bb916f1e5f2ab6ad91578a257cb2e1358fecc15914f0174a9de6eb600645c8a8938e48c48eddec25860d31991f149aba01ffaa356c121d5e611f7015f03e308a5d91c968b30ea2f8a67cda2a1a5948d3bb2e4a86b8ca910596589c3b6d77cf8905a67bac08fd02dfac774432f1cee41c87f7712539411434865d7799aa92c73edf49c5ff90701bac02b3bb4579ac8b8163eca5ce01f25bbcadf7d7601505ae14b799302de3f7760dba7fbf95eea31acc639a13fcc5fcde7fcfc51ea81183880adf3480e50e579218d78e93490818335a997bb0519e45b63da75cdec486626b681b1681a01748c93eb54153de315fbb55a0e751e38f97201ddb4229d97945f746c9b82a775ffb440f7a7ca05bc9e85e302965761b6b1f2866a6ff466b281228a47aa8aebc164b9a1a9c99004318a1ac37b8f17c23703d3f058c638bf52ccb9c8a9d067d47cdd341fdb59c9bc2c11e54276edaece776188ee4c23846ce9e860d180ab570f19b3c8e185541b35e5cca2452bce2e3f9a9d1948de4701c95e84595db6d8a701633a9eba9060adb8f9ab4f0353f2433c971878bc30e7d11b31ab3601e54d72cb115c0046a94faf7068288ac70b804136f1248df0e1293e4a3d7c51b88597dce6b56506c077e39640616882834d10f34356821cd425732024c72389456d65c710d18f13bbeccdfff057699c480342721e50bd3b2a81843d85db980a1951af929f8f854ef914f969240cad5d1f635d7f64b57f7014308e2beb0bee3ecabee0c92f1b339c86826e6d62633bef9dbe1a57fbe5908cce7483ce79eb87d4b20f7897b2f238c3b41e00a4e1d02ffa2f06bb5b027029b1c729238e0615eb51f360cd5090b62a94333b47b23d50a9a85fb2ddd0fbcddb047a4294c525ca58b5c25d7ec4fe8c13b99f09917a6f7be6a0742bc19ac1261f4e4ffc5478dc377ce8bcd050192db08096b42149ff25570fcd62f9765c62f9ac95f95282531e3f38338fbfa8073ea0733527add3b64aedd6186fc88a2f3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3984cf33c8056e52f4b15f7f2d8d4fd8a6305350f5b399a39cdca210e968084100cc3f6f79817d6717f9b004d54b11af28e56e572956290cc8cd7a572778d2cc82ff2fcaeda405f6c15c4a8e8dff977023f0a544c20cecd299bbf0d5bb80c73e7231a54a3462c6bbc9a43739afd2ca4cbe077144ffacdc8dce67eb65abdddef8b9cf747657a6d4ee02b6f24b458ed6aca09e9c89a73ec249d12a6e19fcab5772e3efdeb6fc586af6cbe35b0a607b0e2a5523fa633aee5cd6e490ecb0565e8bc77584547edc982adde93b35404fef6286eaadedb6bae09a824a8bf1519ca4975c0191e937627a60bb03a944d71151f41703370fc575f6ebdeedf1b2e60bcca8341b7e018cbeaa2cecd2b8be120bec3995b964395f2c81c472ac4dc04cc4644dd135bccbb298f6b2717a0f7f8ecaf2a5af8a70cd516d69aefe80368157cc8c0cb360054925de44811291148164668f4573ad6d5edfa633cf95ee64c3546f5d8b423cb6fc5e6a87707a09f333dcdd93f4e3fe01e1f4556dffe253cd059c23f3232fcb470ded020c9544563fe850ded344e5ebc23d7830fa4882ec15c76dceed84076a31d96d3c1667783141c1fe8086f9a0054f3ccc18754019b09a6526590a582a71936503996259f3548f670170ad9d71c2b27086d8ad9b63e57346aa5f6586a46306306f8f98ac6429d33ccc39b88694bc401bb6ff3bdcb5be2d0fc939548add9cb0debcb81ef1069fdb89bd15b5cc526754378dce31898180399bacf242a7fdbf05dcb0d198e5679ae29dec5c2b41a9ad71a666dd0f4e7023a36bccb45c5dacf3e121b75487aa2f2eb40819fe256ba7faa08cd820fa004e1b3fe9065587c728e431e26f1dcac3e65ae702d3ef6d939693655fa859ac82facbdffd8f1285d747d4d0c4322b279fc467b0761d9359385e4d3c8f29690fa66d31f135dadad5eba4bf72587f7ea83766eb733a8c2890bb2dcc89b03363a1ee43cae3ca81900a0b4a36144e20054b7ad52235f594664b182d5406b20c3d2d6f52bf7f3591729acd90fe71ff1be1168394c5f6d6b6a3a805a7b46f229f5506a9390664f5ee80d4ce9d9881de24b2754ebc8d7a6dce8f77a9623479a3a9112341017d7512fd76f2a37ff8f21545faff02a3a2c0430b1aa800fc0003dbf41f2cff3322a773d81d758016e5feed6499233551893a124c4f2c1f8892810c8ecc21664d880139a8ceb08622fc8f7047c6d33be6efb7aca711635264e486bb647f02aa5ef8c7a8bb8f0380d96b76b831d556d41edaba0cf6f9791a58af83569d084378cd47341003b9fe5c8c236f9b1f1e8af9d3766f364baf244d24e6ca502366dd4e883677cba0ea75b9e52e144fd95ebc55c2141336a0c34951246dc53aac8260e441c807326737ef9932a28c8f802c344c19633ed980425499b5ef2c0b5a5f8d2f60522fcf9d628f99ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6ba585f04b04e744c0da7d63c19a14645358acf1663b9fec4ceb458c391b852f1936212aad9bea29b848ed3ec585223e3621111092e1b241f85cb9e8ea2b3881a933702ed1ef2e0a4dbb9b09a406d87a68c20994973373034574a734710eaaea54eb8041fef2b83423513c7c797c59b00468cdaf4097b3ee00dc98ac73922ca1557c20b36551398d324df9e46006ce92ba7c418608fd6af806a31334cebabd1c967250dd9b2e012675b895d05ffe02f797ca8e18c7f715dbdfa2a304aec0c8bbce82ee4c741b9ae32dbb022cf546b352170341c9d906fa0a327ab2c346bfe943db0c36a36d5bfaf5ad5156f7fb1ecedfcf5fb14e4db0fd1da1ec3ae52c969418d70b3ebd344cdf6137cfe2bd6e73576eadabd72822a4c5041af0f47461ea6bd2eebcf80c8d6e6c4980194e0f3c7049ed520c4217529bbc45e3021a97ad04e73648cb61a9755d3506aadb792186b91967ecbc10609f219ff2469ef3d9c09e7aa7100867d725248c0ad57732b277b31d8d9100da280cf87f0f52ab38ca7ce13bbb509a2c17e73a75f30d293e1ca16bec24782543fbe792a23d4a0e779c211a94e6c48e2a92b31ce1f405faefcd586644a1fd44d6ae2fa9f793060fd6d861b948b986bb783660b47fa66893ebf612bbb058771c36ad8a8fcd7b5caa48c8b38b83ecaf5c2848f4f01dc1225c39c5749ef851eb18f420006de82ba8f7e1d82a54839608bd6335e8ab177d6c1ef8d733ca4ee3d0906ea1b03b91c340907c50b9413e6701804bb55304fc1975393c0e5cfd607202a9d2bc078c61eb3f7857d3411a58f9b089dd1f4615109b40283b6faac3b59550d6634c3459708e9c997711ff0ee6c0cf8f23d587ff6041bb7e537191e8388f0cf9cf528bcc81b5c087d30aaae5561eb6d93637bdfd61025174e55472404548f9b5755745b26e6d5c10174e298abb6888e0a3b4573b949c311ff23c7cc78b4a4ff410d45c001a456e75dc3bc069bd4eeb8c096afa2f5387e5b190ccefd39ea969ba8fe91cb9c72cb7bedf8791225f88915f8068c7a6206b78d254eda9a3210447a0a95b6f645a00232aa6dde3d8f274cda3ff3b3f4c8a3cd83adfb23559aef3cadd6f9bc81495f699c2ecf90655ac7440ec345dac2c5e86f5d95cc322198b4aaf453c0cbdeab9f77ebf40ad6feefe3cc6e91040920d8effe3b0d2a889a685f2e50a1b58e723bdcabd135e7ff65901489c53b7fc15b2db1ebdf04fcf886170644130d5146adf21ad6a36c6dfb7842f47e0d2e3d4c2778ddbbad8e0807d476817a0a133cb9d848c540422c6d4c88d7da4b1a48a11044ae24adaf504637ccc4f9560bc1aa24f5014e00dbb0600586028aa4b1eb9ddb4ee92b46947ead6a7f50e2a4d056ab3f0d824e149a2891e59495147c17ea04e666cc300c2782499bce400ff764427a1a2e3689ed7d8348f2f1964c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h902591243dfc8f6c391daeb2d9a2fdf4e824be39bf2e05d3fa332bada643f5f32110d83ffe0fd4c136ed6ec97a0f1d8352477b5c88b0d6cc996eb729f792cb5f27386493e1c7ccd21d9827f80aef537d44938840a4ce8aabecc6aca223c4088f854a25c8355cda4eb914a2a59d0ee8771309aa55b7f4fd1543402c58add254ec569b88aa6ed2c724af9572165b0fba8f73d4010da1eb1a80f67db96f52ef90cc33bbd7fad51754f77cdd0f829d9b24ee6234d838e50f7cb43329668784cc2ff3b269eaf52e5f4150f65e6b09e9b580e8ccc1fbd6dd773f05e7ead78c28980f5462a22ede76607a6db7b3bed8594913c129bbb793e23849aad093ec459db677350ec50553b54efed56a6ce76f70ce1c663dfde1e0e68e2dddfc25521ee30bf8a0cdb5fad69982afcf5e7a996f5201046ca1306041067c14f83d4db5597600a9eeba09b0b57511d4bc32fcc2abb0eac83ae0401f1daf3305215d78dfa17828253226df73b9dd01fcc133e4c1c13fc85d36c71cb8578188c642521a09521fc24578fd57906749ae9f611b6149ff52bf97cf4962d815adbf40468378d59c74f21af0629f7805484ab1377492a5be6ad099acdfa58417303f5b5d7d701f90f430b0765618ac17bc02fc0c7a1e554d680bca4e8cddc12c15d29391cc621607406256a581e98fbb92cf80fca29c263ff0d6f8e68c484c0addf7275fc131224ba9e916cfde0acc8bbafd249f0fac16ec6e85b75687c689d1a93d9374d74fe319d944eb85e541748677acd6e0d4acd3b9ed0029216708a813105890ef11b35164cc0e488061a8a07073c4d545a8b290619e2c527cc4448bd27092f35948a519980afb655d0378186a76dcd30cce858630e4807aeef795ba41143c938781da61f46ab36c7307cb72b5bb61b6c16aee1cdfed5fd5ddffec21757d20769f36e91951face41b8f5e1c73542d30b3bb506dc24cc38629e4347c5c7be4d1204f439197e549229ff69730039246b6e0e6ff6a307f9c7e0d84dc07b1b5f080deeddda599f5e4e66b5bc872a12b64ad2a9db7377c6284d73638e746fc80969adba0ad354651cfd2e485f82f92baca6e145027b71a014609638a7c12eb78c101823dc27640b42600a194517be22867a2fc97decf59a8334c18435e1022f5cd8428a2632e5d9699e90ef3a1b1add44f2121a744ff2ba6f58c5685be0fd7c73f9be3a8756800ae7f785f1ab8967dc359feec3998af8ff4fecefae7258961e23b11d5545f433cd6552ee3d44b16152ad3fe3108692b9382791cb822cbc3af5f395766d94a02bc79c67d43c0ab19925ae09aa8e90cad0c410fb87a881c6dc01276adf5694771bca62d1503897ed66479fecce74a1c3ed1895d6101c79916a66c12272926db95260283e9cabc74ea0e717731b100360038aac61d3c44e1271ccc2115ddb8b37bd48f5724e42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbf5d737a0baff2ca3d676b7dbb7870bf34eaae95833669e09b68578c38271362caa94c5174e04eaf60cdabb9a84b08fbf033caa3c1a4bc37b068166495c31405a6f91aab7a413e2ffc3e1c4786f4fc4b974f9d254dce6673aaac8c71e60cc76a4e476284f9829b10fcf11ee359233c6b3eee2f5093468c04939d424ddbc0c2ec1d83adf706806316d3db7b84bc4ccad4e17b353323719eb79c4e8e3b50cd3286a4e39ee4f5e5546540325526cc0696a8ff725cd8eedee13f2a50144f85de911f24eee111d7d9b2e29f5c445f83eb8561ea44f1d7a87aa5db2d29f04e11269ab48353cf7a2f2ec3b475c7e687350a975e5dd8a4babb6896f95a6c1feb864b48438188838f18c0e2873f4c0019f4f1ec96bf62affb3e5a169c41099ba180acaa05ce3a815d10e55a76521decf0aa5965236bb7a29e5f7a2d0fa1b03d205979cda792a370e639c20a094116f4d370dab66049a432299438ee1524c80ecb11f7298f017fc29ecf562bfae6239c2920cb1a24d271b8cf91dcfc03a7a3d254004c012e7586d4ed6cb33338a93be935336b5fd99dc0c6d016b6d088398569c37e98bc91f6e2508f68a47067b5cd25307b1f1f7dbb75acd6589b66769e014ed8f476455ef20ca271cb8ed50afd9b1c9a9f0f9ed021e0a23a27c3e0dd6b4c7e6d5b87cf52b07b9a17873c45ef892e117eae3d0bc9ee6ad9516cfe84a5672fdf3b038158c5857073efec5a49be974f05bc00acbdfcc30fdb72e705ca1e97700b58ef4b90abf71ecbc8ffddeaaaabec811aa68ea4ce70268866afd654c100fd0b0195014f84812339b015c0b0efa35bc64c24cff17815deebdf803fd074e26c4bda42ce9351b7fe37bfe28b4a0ffd84548bc6f2622f418501ba7c62d63a75d1345f89ab531b5f9d9176a3a285f0d830163f6d4d44d91f4b14ea065806fbacb777ef8101b71ec3d42513835ca16a2b9200d12352fd79c50f8d8587c7c0214bb197a842ab1364cbfe9835d45ab0daa8fc7384b9e10e071fe59b6e896679ee0de082f52e19637b39f8ccb0201280489a23072627745bbb191b11d2905c3ef64b9310c2e95a6c80fe1bd2a8db52e83c9eef78fdb6662ece991b554a6b2eb0b5505d1c7806eefb3a0a9703e45ebed4dceee57cf58131b3a84ef8e53c6d43a360ac4f0c24f3b01d245fd3b9451ee3787a78d560409baab7ddfc2f4a7a130758ad8290958c4d940b58fd7e9afa08be1b1d68fcd0bf65e26c833b4d49b5c327988ae09b36530232140147820eee0ab129abf6af99add89e95a3f82eff4c5186bf31d5eda6db195a8d7fd1d3283cb6dca5c7722dd42df65ec417a90c0e9b2fd643284bb5b7a4abad3fa3c1dc9f656d4082ce3bf94c07e75d5f1a621745b0e1ed8829d15bf4645a3b236815dece7df33e84e7bb458c2877a7dca14ae56c2c12cbebceee73179db65a0838;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf6a9173ca4d2b9694b960f7b3bec827c6c0a22c89ebd7aaed4001fb18ef12f26b22ff07faaf3cabe326ab16e1748d6c793b7f33ce3400f80764ee63ad139200d2cdc4da56df37a7d15f1498b8abe4b6a6d5b023ffe1c224fafb3f87ce6c850179638fe614fd74cb12c6043e9927a2accc81da739c72c9361cd16e3ac5021a0c94f567da47f429d656dc4dcd480aeb68e12105ac38a45ab12bb761f5bc8dcf1f278fa03d7fecfcfe3c7e8a3f5d913d1a87e9dae2a66acba3b50863d4a955f21fc5a2ae4ddf9ad456ecf3796d022e3c14d581bb09171152ca54fc3733564b0bca0b591d47b0727a517a11df483746c85c4488f70cd33d942cc2fb10e301185f76b7049dca9cf26589e5493aafd53c6238939a478a389f633fbd282e0e8f2265048cb0aa315c3df1259440bfc014d5a74d088188312e69522e22b5c1f020b11686b18490b04ac12d12d1519fb253102235d96761ce7f283345234626609a3b5a3404682fee020f48660c42251bce058388d3884ff73777cb490d34138ef2d24ccfb569bd40c893b4f5d4527ce994302a4584829ccd8d79c9df77b84d7fc570ba74db965a7ec9023f1025263306d78580aa6ca486c565376bf5d39f6a45cc2a3396ef46ace004ebb88933307621adcb0b3fb05d6aa75fdac4bac6ea535962447b93fdccabdbedda0edc856deab72a03500288999f97c2ea007eda78f9b50f5ad320d524d64973b05fa0e2004d173e09ce8a67a850252b2591e183c3bdfc6829d0309abfbcda379ef8724d4c3b11dd6573a607ae4bbed2706f038f2988a2730dae65f5c8cbb5de76b0df9b7297ac3be4976ffb1f02e5d140db8793bf875cdc96a56b43c10722902bbe4ad8974f70f0caa9f08925c63d3b0eb0477c3c55a32b6d59e9d8bdfe43e3e6b257488c308f15310908634e360527ce79398da302005434b1cec5a91fdbe5c75afbc9d1e696818eeb1f907a42c1a2d8b6e6a47b37664576f5f978d07ca19e73d91f0c4db349314e77bc717152c4b5ab60a4eb4dd120736386d4c55cfd92c17f3f39271a7f3ca4ae0246165244da1b05b54771e49d150e048a187ac3f6626b4378dbc54d4826b709bf96278e2980d4cdd30caae1630acd31abc30282e088492674118f50deb3e79c7a19878259df63331b4f1368223f0e60daf0fb63922c2f2ec6d56aa0e62641b21615301fa3a02457f71e1425e04ea01e0bd5e998af54358f653e4594ed28cb921cc18f28043d22dcf85fb5ea0a1be15fcbfa85e744d9d4a0962a69ed7893cd14fdd9a882ec8bf5060766593de47bcf6ec5981e3d40d7f3e94c73eba1ba1bb87c61d1476fb860e06bd50ae23178ce81d2e60ebaf45756c035eeaf0aa9d243c4d464e79c4dd1f06b436e67cad1295fb48499290fe7174338abf8a80a016900b54e7cf9c26a34a455aae3af4a5154e86326af758;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcf5b41f97f7a38886a638f63e54e58e8db4894f173993bc719ff643ef12db06f17e770aee26be5f44ab0ffc43cae284872e899a4b78fd11effdfe4defb7bde3ceda737d8af01e46925768d7ce12b8d49272c5d2ef5a1c3947cccb598ea1985ffcde0e766c5204cb48e858af473d32347595240d457a49a87bfdbad9bff10449608e65335aa1135453256bb85af9d4adff261aebf6e54629956b1c809a977088d4814932664d254833ba54c8c1d87b1f0c7daecc3037fa5c95b7b9a85734118ea863884d2ebc0ad9ae7077550570dfeb6a6c1b4f8bad7faed997f90c8e99bee3f7fd0e37a3c381758412ee257981d86ceee65fae935eb354e5b4552b405feda97cafc7d931074af6da91e7e96b6a75252a7dc15703b5a7a127b05e537b58742d3902e0953465de87faf51b5c3d10e6bd37151d5789dcbf00612f1be3f30be8bcb02a5594897b224cd7d7002835b86580068fc07c463f19c0b5ca1868d6607e7689f2c352d3d26bb44e2704959c281acbc93ed8b9c152a6b2b44c2d5c9c908ab7a658c935470a7f367674a24bde25498a2488706c85619c6a7934021c99407161ce9636a7dd8a3f2218b209cdfddd2cb58520ea0cbb3e7ce99c39f65e27162eb4e59b99c1f2f410fe58cc68962ae3c5d206e6a27fcb4d2a66836cfe825751eb57cfe5f2c07ceba19580e2825b26febb55a14d415f1cfa0a9a0bedc47445e48aa204712cf2ac23cc40e0d2643b0b641b47cef6ed384cc6c54c0edbdd28727d512f6cf78aa6cf9ed6c31572e758f9eb9311f6f7f586a430d4d5e4e98ed363630605da8463b82baec5e26ce0974f8a86cd4ad675eb40a39754133df65edd7459f7215b727e958b30f567e8777cdb865b8e57a301c72d0c38c1797954d72e8d76daa93c03fc6eede360a729b97134153202bc88f0421d15d7d495953f9684f2b3ce19d1adc5afb4b8333ac0ec19a682f11a80a79a7801def93146b3f5fdbd42bc750fe9202292b1ee94774ca95178ff4bda355d43bd6312190d3cf9c41ddf1b834b1ca25feb8ec220a2b745d767ab370af7ddde352a56685d64f921f9008e31c655c183a35b7b98677a91ec801e9dfc0c56892f584247a457acd282f4904211fab54eee877608bfec7887c3ad498727a18e8a8e5cb02f401183fd29e00e1c670a7f55ac7de741598837dc7c8be10d5315cc51898450330220e72d5e66ffa3b47ab84dc23ab8e8f73b4d63307df08f79ccc15c563a916051bc7f68578082727e6093101afebf5d38e8833e857bb8a7270ed8e9d07a48ea6f6c95d2a8e18aa7918a204d55773441969ea2f900b6c9b7f684844e6586671a8fee5d60faac7bcdd193ac600dc6b85c525d66f0e375e917133e4372aa10a3272897cad043b8bd7aafcff807d614a03de0d92c1cf73a2e4619db54bb4ec2a4bdb0d2587020783b8bde0c50297;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf8bb0a1cf62936c328dd120ed248517dd5c0c300aa542d18f42a824a7fb13bc2dc9f21b2cd6b925015f0d3d319a8e4f179e061771b7e88627fce10ae9ef32281a2fae0c1c6f303d1df0fe76e21570a6e48acff2af320a4d309078c3a3ce67e55ddf09b3b185ea80cf714f5629f5b0d0fbac2835bc051ed5c95e59154b6d3425c8c4ef2f1433068617f6ac0a274dae165836791beaad62e33b63ca12a52da9183235652e342ee59e641fa6575b70aa5d39306827e657b7d2a98226278273bf7133a6c16a88bfddb520387e3f0e34ae56ed5952f0d07a078676c00b390baec7ab754c02f0a73292577c7d8b8a5e49fe1db94553f58f7afa9ea9d23df3356dc34f0f680931589bd8a5257958c3750a0f99e2321e2778c622303c40925978354958afca9b07cecbf0bfcd812773a45df30eea979813de72cb2e23b4ea96b6713f212c91a6343ccff7d20eb3cdba390b3ecd29a4110025bd53c8d9fc8da04916a87d81552f70cdc2860fe3f94d8e7f88f2ba0fd884fac529f3efd1b515a6b402a93db66de0c8434e4272e02c0adeafdd9a58598907014a8b0a7a857aa161bb5c01bed4f3b079f3f4bf7705beeab120a4f9510f66b499133eadfb0eb453061676de7f2d9b5b997a4ce5d3a4d1cfd2e6ea13b2cbed286014f51f283feba4af7662576ae97f31ed1fb8f7563e4f6c51f3ae03fa53ebf0ac9f775e8bc737c48236ad4ca14ef0fb6ef299a7ea9ff58f27e34a39e2aa15f100890f89ba76d172f2a3090b194767e76918caccf8348236ecc46df58605cab7a65141271cf56844ad5c7b420ab61da3df0b7407558939b07bfea4e6d5810ec51663ec2dae5ee6b4345150768348cdf696a10b7644ddd6debce7439f0c2af449058f956a62fc1271814abbdd2a4ad69d40b4d721051afdbf63d92372cfe2ab7e48cb9a4e5aad8f71434e09eda8621864998d8855e74e2bd239b095a2259d5402abe7f408ca3e74810796a1779b1ce62f3fda93578678d45feb8836da59586df25884424eb284c4b285824d93199153cf7c980d85823c2563701e264fa06c79230eb5129b263f2baa288eba158a898d88a1467fdc67e04956f40a9ad2bb15296f1b6afe11c68e96d0490a36db02dfa0171d3bc34f9fa3460e7071e4dce93ddf87a32841e49ae8e87f168ab90338510a47cbdeb070f268641e008132a66644da6d05c6d68c4f6c1aedf1d47faa0fd3d5bbc1457a51d5c51a3f3fec2e8ad3480d03218f173df8a63da37831a33dc4c6420d75d99dc82b7b598be9ef01e89af1622c970d5083312319991014cd9d6354229c6701aa7487eeeeb84bd9d5e411cf26c0834c1757e0957f5980c53549ef6e58037b3c70e08a29b257d7e6f4fbb9556758b213af849c169be07e2353e6c94e88de8cac1bb87d929440570ed831393c4b58192dde895fc38e88a6072982ab4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc9c6ed12b60b29dd1f05580f70616b0d304ba029a8ddb9f45d405d990b1ad383bbc839908097dcf7ca1dc602b7ea1b989b8e1fbfc79c7095c9605c94d6e18826c06e8f586ed56e93526f4ed99b195b006828a87035ee7ca86cc35231457c76775f16bb3832f460cb0b519e15ee4005396ce90991e9291cdbe3c38bda88b410b754fb33c0fa0200271371454de104a68c49fe457867e1c2eb6a718b9bdb4394742211201c71611244acf3b90ac379586b11696e50217c1759758e7b5f2215c50a59c488662112382b1a38742bd0af4f00af6433d4b60b7a7565f53ff398d08d2799f9405aeb99a227a5bd70e44024f26715a570e2a33a2a835000b0cc4bdb6d288ad7fe83ea950c37afd8c31feba2a532e22925c85dd048546af9467ced813b2bcfffb6a8ac30462d4fc07e2566d7b481814ddd1100fc64dcdb4136d1a3152678d797f84749d9a9894732132dce0a0ede2bf166ed882c1b6120d0969f2cb55add2892f0ccdc5d34d22b11f80b2de4c2fa3a56a9013e60a13554f5c91f683c9b382c26e811c3d9afe3ab944823526d4ef11b2c3324cb687f31b1f363045b8ddce0a15594890368a893aa4106e804dfa52549d3e523567e3ac94609647cdfdf32169bfdf7e007a4bcc5c0b857743415356051ccf12088202b44aa75381672817d33dddc74397b5bc723e87456ed7d0019f1085c3cdd9d18540cb14afe529ff4a73bff6ade920a8c9f2fcffc14687bdf8a95018d0c6f5223908ff6a760d110d728c658b14de195a7db07b8fed51599634c9d6e5478b0eeb96ccaeecec32c10675c387d69d69f8ddfaa1df854f63a8cec2939ba66e26b8acb550d0e5ea3cf19822a894762932ce43e8675d8d3cbe0a97dd9f7311d27ff6ba92f8b491b4181ce3aea52d5d1eddca0936f0cc434694cfea76fc27ad0e5da79fbf32f413aed399e7b17da8fc94a105e9ffcfc65bdee92b3842c9697368522b7b0edd581a86c6a1a0c032274cf426bd48d01ee35515ff0b87578f9da8938ff8541ca69e719c54f2ceab5adbf299ee4156fbd51fee6329ce69131117119a7726681b1d1ede39b79e1f9670215ea65e79bb71acca0015881be2173dd229cf61431675ad4af76da4898f3c640e90d9e1d897d3a4340b662bb29c67a8ad333a5a4952557ad711f68a3c072de9a3b0c0ffcc4987ee590e3189948ef5e78e3840604b7aff6073aa739db8ee37bb3592cdda6b496ca5618470fdccf72dcd8175de7fbd6c3a6a13e0639de5b8398534efc3d11e289f52bb58b5fae291ae95c1cda1de235d6b9f9538b9a8fb3fe2f9e82d707d6c02f48552be4dc0fdf0e300fe63552147f6c9383eb71e1766f240a6ecb8c6c8d899066b117ba8112d30b03ece3cd656cae8296f2f05b17274426d973fbc1731fe16f11e50db3f0e273c302692120e8ca1076a0d4923def36a2d056f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he0a46d73b78a819fc9266db16a565e99ca7cdabe2e02645ffb1220c6bf8c2683d8eef3c9ed2931b16796873fcf6faf90c005a445a9701b56739d221a14704bbf5f008b092f854336e731a7f04a7e319309fdb370d195740154782782d00ecc45a8b88b3402f3c10f3fb3a48a12f724dfcf8fd728fb9e896d525e3adf2a95c99d12fc71d45fabc70c78d0eb2c36c1ed306e5d8853dddcd69788889b2ca6ec8a87fdd9d41952208b45218afac472eb18ef16a3c354aa407c04dc710fb9927d4c3db12226b7b815f2ada89454ba3ee320ca7beb373dee4be29f5adb02b2b9059d67c54e4dfa5eab9847d5365ef611565e781986342167723e954f8704d802469d0892a550417ecadd6ac5609ac5ca79b0ff6eb32b3e24fb1d2e2751672260d3b9f7d2cbf3d4119ea1f78966ddc458348481007aaa216483b265803c0fde19958204050b5dfa1086ecd00ea4ba84670d10a5661990888c9106454bcc55f383a17b29da7190dfb5f840b5f2db6d8fa57cf87b4547c326611be21e27c37146ea727ba8defa360aa6714f621efb6e0c9dad61012e9b94571da583eeb514658c05d9b5c4f1e082320a6050de9a48e39154262d821a235ada9b966b5aec2f0ca7262f672b0d4685db72e79e566962ab29a11b4346eb2ec600f1f28d39949a38531bca5f4bc991d7831a5b7866fa521b41aca78730a9ce91b3dc2ddd362041e8edce196a4dc531e1a01591c5b61e6b8aeddc59bc1df4ee16b3caf7cdecff8497d715da9a285c70651b7b3c2012b7b8be942820d46a9a19c56383f89f86c24dbc7cffbb575d64150e9c0b9ab96766c4e36b6640b747421192d88366d228bdb62f57499762c419a8134bd24b1cbac72b8e601f3a6edfdb742bb6c03207fd129f1e128b9c0153f97acb8f9b1084d1a35f74463b5642236a4518b89fd271da5dba26f3335d9db16051d00ca5bc81d41d7839eeff8bcb7a77dc5fae54d80ee91c1c6f281fd05d87865de2f8f2c2fdcc3c323b88fe82f47f9223381f8d37054d5d7a5f6b09e4419ff19a2161b144a27f45c94811b8a6be20b4f683e249a4a0ae69958ff6f7dca5d73ce981e83c6a1d337504c18beb888c67a703d3196c64ed21806b3eb90336636c48f77b649cc40c23aed38099264ec28f9e94e12b75c8d4314ee530ef8a8bd64b11c03f25bb07e93f782a8b2586ab0a2e27749bc250fea310a41aa600535d9aa925631bfeef9d38306edc20f814a476017ee5285d8b4a2c1329aa5575d59e428e7a92c3b3a2e6171fa4a60a1b2a3eb3b9fc81ef4c4f254e2cbbdad187d093c6419da607c22ee471b04d6a03a0992366d1db67a787aec76b3882929d709b68775ed3f9736517f046cf26ee9c2b0d920d5d8a1e7d2efdd41410a6cd506098c1bc9860a483d0ecc980af69e19e980acab8240e36b480dcedae85c21364e104d3bbab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd6c4e8c248031417decb3a9a18190a86634ad9c98c77327d15e3ccd2c5966a40cf8ab210473fedc612d05cad13a5cfc444b9844237d9e733876c744056a0f4ff78d6a9978ad0ca56830249a9157be08cd18333c8e5cd65dec61edb9cf99b145be17ad1fd236bcb50a9ee85d68e7b848bf2ac897b5ea4109537066f35bcb32056ee5b8425a17f4bdf8b79b4561128e70dee6f7481b95fe0489d24335e42eb53e4bb7da8ed0d114f2d1ae120e5401bc51ac8c7eaf1e862e81e97557bd23a62ce93f53dea72f451d4148c50652fe192d8a031ac1f0bca961e297d9196fab5cf76663fc948aa69a41c88d6b220e928bfbb55d65a219ed794897fb19b5a4232d3fa7753e8d76136deee06c0632ab74631de609e2d5af8909f03c8f39a9cd19fcca63a6dbc08e42fdcbb1458a6c1671919caf96541f8ed9b4aff6fd58f4b19ba9dc2a1e48af9746e173e75ca40ec450d6d4450fa26e3e88bc76946cc807620f5d13438a334b8e4ee5af94c9e5ffbb4b9e34b132783665f612ec2ffde74987f9fc90d93edca3d54971cb759b58caebe317d43cc58926b186aec048211f31b73da5622b14fc86ade174342b3a6b85632473e3a51a0ac22441aee7b5a98b37c8862588a5ecd76da24c35c7b99569fd41df59b2de0a486a1cb879bce0467af55ea3872919af59e795d33b90b8113e3a14de138d361f18e9d83b6488cb2616d470d8f7e00a58635533cf843a8c30f47bc32b72a808a2e33a8778ee1c5d319e4ce0ada6a67569027188214c9621d0cbed57461844dba2b0b2d93094198b788ab8d92fbedcaaedf3796a0778f3bd5c4933348e375585426811a800375f82c969ea8ae180ac14646ad7c9d5ca26879914be6e8d9c25c0aea657b52b1df6d76ff1f60d6b770b8263449de2d4ae34adde1bae45acfd0713c96e50302443b6ba3fc48e1bc01965139a7bb98431ae537cd03474d173f892ac54844658d6291f0527e32c239528a59f87af76b5248f74c9ac4a9bb1d2761d2e9c605cc9415f99b67ed4d29daa0cc03a53573a3170e1dd990845b393ca4bd4b82525816e8b6414ec748ab52c11d48f531acc841d6fac1c1022938a2daed52d5d22ca243f50842291bbbdf9e7c3ff97702471aa6f11efffb18f1681faa4bb66530af7a7ecfa87ddfa680fc5a88e1ef0f347f642210a04234813e02a341ef61a35b6879e28e4191c4c122bf3893291a90bd21b8a41e2f6757a238151b200cb5d65dab1f1e8147a6ee4f055155547db9c2a6c04b4965ba2868148e344bef9b078b9156acc98c621e2e063334d221f49371b43a8187303720a85d459aa926b6461f712514b49fb7a8f5562474b21f594e2dd44cd27d7768329d198dd455a31ebf8705df918f9a2dbe74511d0861b3f426805735c91338b07c010f596a9d6ce9b9571c1b9c48b68192247d24625e40ec3d8a1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9f0803b77f98736bffe3f26eb160cb020f4ffebc4ae475633ea58b5991be198d316511b9b71e8e6240b090ddf48a63802884f40fe5275d8611ef0579b28b1552a48bb80c4261ab53f9ff7c65b53ae6eb7194f45dd1470aa1651bdb298f41ce88de56501ea9a6729b46c3040c8fc9060861c1493a237b3e07da4c8188453c5514d1407ea037534629eb4ed86c82ae73b180bac317109e020caad14effb460c88d8792100415fa193f8a19efb2413b7dddbf53c15ee273d6b516d52d059bd9c04709db5b09e71241df7f0b18730d1b1edcdc8f6b1291ad923a1e706665ec983e3874a4c14752070804ed28a820474e54c75320e860233fa7649786774a38c79f33d1f9b291c25428803f46e8295be883b8ad488c68c28a4d1e6144f9e96ed8fd401c3113fecb98c459b0b16225b33960063e099baa99020cd5718a22741e621f0f65eb84c8345f6ca1ae8622d9ca92a3bf9c820c135eee32f443597173100227cf0ce12a052bb73b9d70f247e740606d3f2d3ae46d8212c09c1b8a5056365c0a9f7c29ef016d07bd2271572259f6ce1c6d43730a898cfb5a8660cac45af507a7ce4b781e81d58d1136f6de2d2b1dffe68350834b63c1bc4ffed09734ae902420dda877a5e84e93797db9600b19efbd1d27ed1100fd6a69e1d5807f26241c81ce45556171fe6a81276d20792b02792b36d1a70c0106e5ceca7265b004f1c119cc1a56cde9ae71b9458a1b492c5be9149f57ce71dfe267295bcf9394546950f3280e18f5373041f545b504c1ef8d1008339a633301f24069d995eaa21bf2f8b0a89d41618634c4bdd1c03a335a1ee2a2102a431c067bf04bc25a9b886ee8b6a5e4b29236e406feca7707c628b8f022a49fc84d91687fd65f9a6c280b0578c5a6b0d2a5bb7020743414c2ae9be118f010ee0f5dd6c8314c1d8d2b993a352ed1e5ba862ff801f20d4e35ff0460c85b920dab33e1152bae6d4e81e6e0aab0ecebe6f68eba5c8ea7a2cabdb9aae6239a2c7da0bd45b36711e181a89c9f44c4a669055ecddb872494748c599eb2a3f2b25cfe882f2f324741058804e4fd50171ced277d2da250ee55947838788306a54e1c4fa60aa2c125bf0384be6c57b1318163a6ff18efeb07f8b6197af7a40d82ec297e8abd63673e24bbfcd3d2112e3a21088ad9d40aeded46931b093552a90ebe07e0bda9a70c3d4e0d7407a8b5f7e59c073e9a253bbdb1dfbcbdb747b68778451ed4f735c17011e02b503351e8332cdd6920129a6dfa3215455db1d7d2eb02a25f232ec10bd59cebaee98749fe6f3a9dabae7ad71821371408850cb27c5eadf8889d51f693322280a4d03e5c82cda03bfb4b12732228bd34ead4633c67b95a2dc61ca1fcb9d212415de760acb500a2c1d28244c2a179779b97c42ff1ca8b48334c389b92401378a75038824ecfc335a4cf706360;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had8c3c39a29c82e73cc44f226a58c467137ea64fcd21c5ebed33f13f5f1ae5d39b0df231cba5649e2f6cc8977ff0c2a601865253ba27b51b9b54c21f0d4544892197d58eb084d275126d3eb6c04661543ce9dbe045219800a1649586d8d3980f8a18b8e0aaa1bd1ea6df35a622b2bb820a7a738d60d2d9239e5e704f9b6522d994232f540f7ae963d2510957fba8010229ae939bd086a9c6c4d6c365b4e4392c3082e45dea2a4deb667033fd72af099a3aa06daeae944e80f5304489888aa3770580d8f1839696cf5a9f2f8e86b3e021ff65fc411a818bb2ddd8bab9a74fbae31f94b7dabf5c0eb63272edf1a68689df9901f81e440ecb13d36bd278d7e2459cc022ddb3cfc19d9f22577b83d1b7c434f6dd6b143c0b19deee64154fde78022a83416451dde3424ed6c8abd5f13584d2bcec00effc9ef2c41271792108335b9a099b8c9d275a06283c58e2d9aaef28dc9f0bc7fbccdcf76bff24f52d78ecad2d46f73ed6a5bf066f402ab55ec542c7ab51c4be199b7dad48bcad38478509fa83b4e6680e744830e8d442996f08c80acfefaf9a8e3e85c84aa4cfd5175063215126498944fb04a255196cb0e559e7446a47f441a9472cdfe01b19b63c90b684123e1c91c52a849c0763b5740deb58023cae956cb1974dddc915d19a617240b4d6e4b08d6a4aa6b7100d8c9717d831f88c7bb62f7b3c9b8e5cc0a3ea8ad5473299a0933a68e624c94b7312c6ca3ef1cea4fd30c0ef008eced3bd7e12f38321192cb8aabf035a16a81bd2fa866e8c2bca76fca000a91ed21679943f3120fb9201022f4fa6be19635a2ccfd46800dd54d1f79c7e541fd7dbe9100c41d95d9be936d719b76264ad97ad71308dfce9a12b4dbc3c474f82e03f5094277f2bba004c7386c3e9938dcfc8283f139800d4259e6a44e03844e83a690d7513365459f624182c064d790225b3b26a8549029bf88a1b938cc8ea6a07535e318df360621e56c492b07074383a17bdaf7c7ba1ff7ec509dc58f56023f7ab5db6313c83dcf38b4461c8edaa8f429c9ad306796ea2d520ea360580f3805016d2d310a06dd9dce198d3799f7e8f32100ca52a6462bb081930389f4f24c08aa3f55e4f03339e4171c83478d2313a84e7d06295aefdf895a6b765f8a5c9cf70511cdfc42ac92ff810a19aee1566b31a1ea05c6427a7094371de7c12a5b3aceaacd31f5e37ee193aba5b5abf9ba35a3fd104d85d0dcc4ef03aae9014d90f3ff0b32e016c473f772a85edb29ac008dfdcac83012d1a70c3eaf601f668a7783da748cbf9e1938d3ee5fb9db507a559425a26fe207c896069670adfd4a51ec2e579d7c21072e8bcd1dec60b76c046f7fe3591f5e0be6baef0956424b1760ecfadd02ce8536d27ea7d4316db3c7d4bc65d1f869aa8ac2ebec23abe847f3d6e9819dda7c2e9448efe6be755a68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8aec06f8ecea2f0b71890ef02a3efcaa851ac7e1d59fd97a999cb8416202e26f32fdf3ef91f9f7ab2886d21ec2415d7f5dc17ea68f47e7637da377623c5b9e38acffe7cba40530eb9d6b1c063bdd55273e2dedc988c437829a25a5dd5d69bc7ef836b3f5382cce9b740760ae5d0442e639a68d2da48daac89879c53b8a2fc857d57a1eaa2f0f55e1f76b066e125a289f9bc9d5c4a88b9aa8f34654c9be72743733f474cc4b1de09d1080557ccc0bbc24178367e4b9a7784d8ddae5b93798634ddb73246e5030ca7d88378e18898c59d255d7b8bbf67501690774c1c19bd4a6bc5ccf688defc7da72565bbd0baea58ad9620136947e28ff9754835305ce21c671f8059aded2467f57e0e75503e13c180db2edcb876d5e9d3788e086d7767404ce08a120cdc5cf95825f140f138ac82c7d73a929c54e89c88edf4232bacece861db82c6c36c16952d602fc32b4fbbb2771b2e775721cc1e99b0df696c9a417da1078da0100d4227c2a0beeb77a825848091fd65a4afa7ef4ef079065f6f20ac0b79d944acfe84c017331f6528445c3e801c624c36383616fb4670b175862b806b09e0d7c8b4820867776966d4a8f1d2f8dbe510c5680777421aa61d95a8901988dd6481a361384f1790d5db95bf6c78eadd91d1f8da3a9ed28bd8794e6c305380dd2630ef6f3b287344d6dfc27e50f149b1bfd9c93bf8d054abc7deb293237db8defc2bc16fb5b32afc65d635079243cd58d7d943339f28c5aae2d7ef72e53344b3c4c6bf843e8a839804b65b1b54803689a753671f3c4c9dc86241603179124ff64d295a2c5490cdad8fab87030817761486eeb0a9996478e939b57c4101bcfd98e2f33262372262db18ab3e51c81339607dc016b2e0deb6711796454dd2c648327546302615d802e77fc9f2e0e64f4b4efb8d13470510a2dfc2517dcd119428c62950ee01a29c4220de3411181e3be44c7239d137fb575748d562557d6975ef0c86091ea94a1fddc6b709807b6a24b67cb0b17ddecc0199fb4335c1c8bad35ac206d5232450f5e46a31dcdca2021acd5ac7ef639e577ebff3d644b91bc9cba4cb65cd9d8ef77e55e64f9ddc2574a74e4258407175bf949ee01b0a0267070e55ec3ab955beb25c0d7c46137c724bb9b08567f276f33fce41a4b4335d66514d6edb9b46fa68a4508c5f9caad65e7403206c3f4a321bcecd7f21efb70415b9f66f55ca724d2a6db92a4d4f682d87b756b131f7d82c3521000d1c9b96f57fb2699136dda112625857cf62dc5813be98887994a49aae4c4ceae6041c77fa66c8b5ef9246171e2b208ddaa017a74c9485dc0c73d791e33b72fd3b6b77a4dda68c7b3439adf222f22450da6969dac0c676e3ae4f2fa4b0144d61b57d4d0ad76558f81a79ff30fd6504e290f6ae197a84f63ef976c968d9198e931dae5b0b18bc04658e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7348ea1a195a894c034d99e6b86d2b8a37278db032500edebc517d84f9d9464fbdd1f543a37a8f5cc82995a3272331f4e08e746ae746e89ff1c37266161db1c4216fbb49e44c7bb21c1192f341337bd9f29a809db55aa340cd3be77f16ecc18989bb1fc7281d4e51a20f17be849b5b80ea0349ca47eb129a52c1b0ba7e5c66e7c25a94195f50e9e58a450ffe5eb7a18b26b2636dc66013a97db37eaf5a145631f3f282669c7aec9bb240b0998afc57f18fd4a97d2f74aee797eb5cf4af5181f7472733626feca1a574f45e51ce62ea945f2de78de739ee7aae961b960ba6645f167ce8e47b504a181c43128460a592fe1e1cb5715f7667a2e7d7add949ddb4528a63b426224a6e1fcb1109e6079089c7303ecfd0cd8262fc14344489857dabc6c9f720ff8df5a8104c30fff708afccca40b2250ba26b1c47b1f67523f4890d5ce556460158462ad2a7d9250fd754c7867722df4af06fd4fded4365502e5e6802faa5f9f66a82ded1f991f487e9f28a1af9026b91428c21ea1f899205a5246f617ac7853fdfa29431f3ee2636b0302e31d0b3cfde6298cac61933264f88b4089f6f3cab5515e20a051240a8d11f6cfd648281f3d7eed82228aed2880b1e496d000e4a78a04288e7183cdc4f0657c243d98ceb46f76f4d3bffdedd0ffb0418c6a7da1f6a2841931370f641c62e0d91e63503229570c47fb7b8093b24781ba2074290b97237380dc88d404f6d0232cbe5c62fa91a83753732eb1fcc28196f278dfcf872c8c08152ba383bd5d699dd107ab8fd5f2bcb24da30f8ac1737d7ddd767d435786eb2d448fdda77ea246ef7b6d20392c682cc4712c75a9118c7211ea1274793c1cd91963194283ee2c10ef145b728e553314cb8347d372b9b2f53d59631ff491b16d08f4177d045b606273e085193c94ebe40f9e663148d889991f3622ad86080bf2c0c49d12b8a5e979cd06a488678ba4fbe3a1a5fe0effe03c9d890deb5a61f14019d99f46f0f24a66f4f488150a1048d3879a20222e98ad021207814904d12b9cc95f793ed5afbc4f0aa2a908e5f09ac02189041d7cc0b324f08b359755338584e384e52978fac2fff7d226a3b19bab77ed6c87900fd0faa4f8507b0acbf01b8bcac867a7c59d84fc3ea7e871637eac8b9c912a99ab4361074a841316ea191e30d8e05b297117860f4e7298c2f704ba3e6deaa121ead79b8afd99474eb164c8fe236f880954abeebbf14eda9bd14e39a9d41afe86923bbddd2dedbdbf8ee89876033ebb0237ff3c6a7ee1cb81b8ebd52522998f1d2bfc1bd66b183b5edcf7c8788fdfc6c3bd66f1ebce09dc31afe918659fd28ecd3b19fc68f8436792e10ba58a35a923a27d87355b221d9dd61fd059d1e697222e1d26613c179412f8c51e1105f374382e8331b92bb70839f96ed2fdc7dc85b3c217cfb021b4c55eb1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3bf3308f47e9fb78f168c99fd56ffb8bd09e620f6b025e6482d9cacfeb8a4ddc24a06c51681babdb45a0d1bef79a4d4e1ece53502f3a415ac5ce15f41a822e5bea26b8c0370d26eebd55cb917765d89046d524fb29306baf14bca2ffc4337302f4cc7c7deb8e263c6dbb1821ea8ab79c35376f70a4e6ff89b7a2c0bd18513878928eae407f90b4792924ab343971ba948c505a094f473d4f9293337393744ede221ac71a543edc227ec3369f72f84ce625d44c5b45847e688fc5f271e7975e0ab089a5eeb848204b4abb2238b087829c5e34e6895a8152f366a836d59b87235a093b9a2f92390a4bb97803b8472f7d806442a107b72dcdcf140c63921490ecf1843e6825f3435c3efb7e94f482042fc9bcec9f821a7fc6cfad52b7696eb5f22eb5de7ca0287983d899cc83d1c2dfc59043e7af35ba61c2344032f5899f20ba85d38fb65e08f0c954158c12193876924e4ff7cc4f22d7b17d2d934e4ddb42adee12a9fab6651dd335055e9f80c427dfee71a5a583de1fd2449ad7709848c1d1c582fc76afa067a770a5b6e566f9281ff30711c06a8f65850b2fb7bc4dc01287874754910ac8b0cfbb76a194067edcee57d975f60ac1e4d7fc6a85ae92194a6856b853c8ce0386306e42f2201a1f04fe0fd6fc94b465d6af4584b831055ec1127a5f9733263fe65db4e2bb9b52b8454aecf9b59b1ec5fb9d9441e5569f3a075caebdd6f7c6df83d196543666c6ab4b5efefd44f009882f51e5e256f450eff597d6eae18b482a6eac858f40de8cbfebaaf17972e66d5c17ff1fd18f55ff5dc153d99e98946700c6dee2c6f18940d1f3a2233a9ac21001fc8de39b460a2715a81b12c99f6818d5c758d1cb971fba027aaf1e9c46f6f8b35bf4a58058126d70cfbfd44b8a6e542056ba4f8f10973a47256413521ef49950e5adbb81a6570a23aff6db78d44dfd380c8a2ecc38bbd34d25338459501fa932fdd26d59011db5391f31087fb4b705948ba452d70d8f58ee63c08e5927ca83d02fcab99d3dc2537ea434424d6e3351740f55bb688bf7c564c6a489c3a550fb3caba58cef54033493869c8e2ad7de1231aabd333eb9cde351f7491a1ef1eb8ae75fd7e62b3d3ba617ebdce63ae1c1646f281e77dda49a712334e87ae822df457a4d5ce496aec300b85f5c0301a52cca5f25209c0e23d20ba76f6e0fac23658a6de00ade2ae73bca7226de002fc1a4dcff5f8d36713f84258da8077a7e1ea7743f641c37c82e2024ee6319c1c494a51582dfe9dea6567a6547c25dd4e0915bc79974caf7ede75e320bcf9f5ef08fa481ff809c5ef47eae44a5ab0b3bf284c43679196bf60e68f785178978ed6eb3fb8686f7e7d6485feeda9255ee81d0d125cb17fe4abb6a5de5ad5b794ca5e9f036750c8445f64e3b067f444bcd860485ea401a7dcfffda4b4450d5891bfe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8ce4ec05a0edc183039c18b8abb08dce3f5b0d46ca062e601985bd0a902bb7ac0a667b0c5e2dd8d777976979e4b36ead7930e9c1331a88081962998c65c6d3c14dc1a9194b7f2b356cd1031f593eecc0a9f80e13797f08ef0e8f134ad26fd26c883fadf667c72a1b24432ac56342eb521bbbd90f12220d5ea968e97f160aa1bbcbc11aee37c18a77ef559f67590b428741d277abd9e7f6368b489b963fe36db5a6613fc374e5723f3c7f0b3ab4cf4a4630436ac4bb31463d401bafa9093b160e1e60380d1833e5e483668d7db0ee3cb7a689c25ab57ca16a4be13ba7ed54de040d97d9911d1e6a965b78ee3c0b9d1ca49bf4fd6fbb7fef748bd2ee391f152a422cf526ecefaf3a4ab13ca97c2d97bcacdc51c0a23f92dc8307b5e2b6d6b146db662617044dccb7d07effc7dfa84358b5e88c5c83b82bff5134716b50a68b87f8c7fb0be7d457224427abb484360d2272b9389ded9ba288987cfb9cf48590c331670faba6b09eddac59e897fdfc667c971e320cf6609dedfed2379958ed6648a563fa5859e33c9287bec50da8f507f280b5f6b0837bd6846cdc55033cc62ca3f3198dd890d938c87af1297386504fc084501800f82b34a888245f50b0d2da2b54d5206dd7a8669d9470164c1d03a795092dab49861ccf60865f9fca838b312c303727aff451b3a0b3e639502e67d6756ba089969ac6957e47cbfed09a700bdd743cb46c3afcc43d5a7cb2d15d97c82e31f9d037e4bee03eeb7daef0507b62ab7874bf01cfc9b6c1edcec6699c20238b8960028e9c3cbb946c1c0327b16c7ead22c765b57c3904d089c01b0d4da292f24ac781751f3a35224c7393e67a9c1f36ea4cc0db20502b5aceb9ab58e4abc7850b2885d97da8dac2e92522735b03eca861ba0dfd98dad186479abdf04c632b48b660115fd0535924be38f201b7ea4d7c55b5537230340f03de4d243ff7baed09118eb0bfb987b718d23307b12b65db46f07d74aaf4d945d8b81c093204e7107aee5bcbcc7f11de57302409ea532d9f6e47a5f3efbc719a3c2ae08c354ce0c1dbefb5ca1a9a317e219c82abfc4e229c0c3c9db739f48e3dcf6b331f3336b6c05d76eba0da2317a8e7fa29d2bb7623f0332121aa8d52a28e0fb83602b7700ce51d03613856e5e9b49ccb191f41d3ab7720553e4bea446c125309f10ebb5917b5931fa7eeb0c808e46bdb66c455e4b5cac3afdab9e364656b3cbbf89f5dc6c08dbf651dd4afac5e7197234099ab2e7835e3bc47aaf00051c31d49dfcf9c662f902313204cc23b84a20f75a05d48d8a0793309678634d37144aa5d412db3a899b6dda9e5b603ad71879a981e98d286a84ac5f94b4defaaefeade5946ffa03fd571b48934ecae221f8c4a56d50baf54d2c4fe67b59452f0ea244c3f07fbd4a554568fd20e7f4757b65c25def4266a73a8f6761a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfbace3f67893f78f6e632cea8227b04e641be2436dc066acb22429ee67b239e8a1072719f3d3606eff2a4f1e66fbf5bdea9c85b42a92c16a724c5d1ff43a8341abbef487a2c256bc171ac18648da5b8404823db9ce6b2c0617396506c8ef234ed956b9bea7f3fdb192b746a1403e47807e7d5988bfbf73fcf71c78f7c8ebdcb3fff12b8082e45d7d176d62d1b534b3f5b66bd6bda8e166e0cb7e7a550235c1a534accb953e508e60e8a3907f214952e7dc94d88038bfd6a7ae31ec57415a1d42ae7a461e071dba0211c53fae14b57da974f29a240c579cd00861bb3bd7153a0b7343c54fa2f7c35d3719c62e4370c28c202a33fabbb97fd78ac89305f87a18dba8ad6ee7a990af232696ec6764f3c20176357e24d948dea16db8a6e7475fb4b18a9fe72b2cae9f7a6ce7e96453dc9e33afca0e7e20d83cc594ef75d9e3f5b430364cce76e882905639af8d7cd6e12a096da0243b2ab726040ec045601e7c7d97771fbaf8a41f2bee3252b8f231af14433cb64a3a105a4210754738aa12d7f2eae3465e74abefedd1016a162606d157a084a0bd052652d87de06ed5979d7ff3cc473c2035a08401b59d6f6f95ca8b1535015ef241a6a980c7b18fa0416a7e5bfa5add84506298e320fac5ebdb5eb32570415b5e519ac71e37b3b95b13aded28ede9b26eeea13da9fa450ba33b7f62581bbbad76ae26034ae8a8722f0ee712e61e7ccd14142e2a70912cb9cbc1558df14093c5bdeaccede788edaa66c9391454aea297a5d3d04ae2daba5f51903367cb36e7c6a239759858f3800c0088c92f7d31b00f05bb9c47edfc9469ce16719d922b643521a257e780109aae256ce69ba6e4f2c4d3c154aaf2df0599ad5031b1286e552946020a6d27c051f947af88d3611ac29cef9c78e836e1134b0422aafc844d25d0f9a3b85a9bafe44eb8189cbcaab323057678d91206c88f77976e66c50c84cce5f506505fa6cd6589617ad4bd4b31977b40a986492475932f29d0ad4cf6c107d7a316f5cb4c9962df3ffb5873e3797e77ddba9fb9be8dc8a5eab7bd33c485cd9d297a7f033fb63d729d7f8ad0c9eb97e71ae435a2b772d70fb4ab09d476d34915596b56db38327b0889641cb81d6eaa1373fc6f35445d281faa5ba281a55daac0b7c36c0de6faf5625f776e5769b85d34641cecde6edd67f625a008a61f44f062a05190db26ff617fcc3106c87460b88b52788682baf2c2ea2e09f570f0153544c2bc40fa5a7d6f0544ac2ebbb070e614d1f56aafc5b4c7988a0851987c505c4f1bab566b80d0d25f5896603e2c85855f7087f0f05ee2c6595cadae4a0f191830386d6685d30b4b4ad7c61388745eb0ac3b35e4dfbe3d7860530ba69628bc429426db55e26c03135acc6624b00c40a99c6e83b3b719046daebf9f3e72fc1ea2c2e7a0039e503b24d3e8cb0fb98970;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbd4ff2326cb87bf6577618646686e0b1029171ef7e3fb3c109626d883cffa1abd562d8bd7db0673f801be35b1cbf76214e76257e9493812b4964fa1f50d694ead7c47647195660306eca811e2706c78404e05d85b2c9658bd280c0e0b14e321df2f68c64d97199ae2cd4d861f17a4c12425338977dacb90f96cc0d635427f8cd7b2d9e91ccdb97874f5c448bcbc193a853edf09bc9ee9ee6f3d9f33d5aef33b50e1818823b2bcdd92ae84dd1fd1b0613833ffb523a55bac7a33d3a5b520909083021a12140da94fd31340e327d713f827cbe3dbe8fb78338ec72ea63c448c488a329fc46a2586abbc9a50f8979fb1e1698c4f2a2c9e7346d911a64228a79f0ff3f89e876ecf8ee010b02120df7ed459a29722e029a30965a7e1a7e9a26d162b441858008e0cfb0f8f6aeed15a09abc3978ed05a02c18fe69f53e75af8b1fb11cf0de0ad34097cd090c01b5be38240e0ef1f4bead22b1b05134492815476cd92dfd5e7cb6fd6f1ba55a693517adc4689efb03158c69bc57f7ea513fd28c10a7721449dc7492e2d53a749dd0985c63d02185ddf57e52e5c40b8e3069c5e0ff67b63ac05776a68aab2aa869991e9bb46fe4bc52d725a39dfcdd156d43e08b6ef1a421e49ed9fcf0be3595b1d6300ab375a6b0bfda8a6573d6ac9742ed4e96a8a953d331ba996a04dfe9740583ae000ac6a1c3a2597ec4601e57f6549665b5a26d8ad6d0b66e17aa78ad80576aba97ce5f8e3e4e3907aebe0671a92320427f97d0c406204e1b2e182306710cf91c6ec9a28b097e0ae950b63c419d0a8e8f629b9105ebd59e2ac4d29bcaba5d820654a84667664ba89ee3319ea6f0d03a9dd65f399a76e228ad230c8ffc6858c71ef94be54e4d44a88c0f823669b19eba7719e3e74bb585baa2b1ad64e79b8d1b7e1d1033fda06d2a15fe39fa94a2d5333d3b22f0a776e51577e96f0f5c3316fe3cf1581763ad2e45794fc583839aae468b6540c56e75b41495208d33c9d91e778a09a912072399bbc0486a887c11062764d9c805e997bf55e448bd4f190b14d98e10ee24ee612a05b7d6b869aad3654994e0f7b1a72b976f38f15c5a7169653df142c2c5b0c1128ee4f7a43bd4943aa524ff47f981c3b320e825c0dfe4f7bf9848113587e4057003b8351456456a40518227c144108f317195629f9e8bad0f4ec4de6c481a42eadfad784574d1720cf9fffa53be482d82982bc67bd1ab84c8e4918c8fc43bb165c2c140adf2b63fce754ac1841c3af597cca1f90b97ee16369854a6129a78e598e6473c648dde0d110abeb20499cde26538970c43ba27fd6d0e78055bebe812c2228808191ecc213360af6ad5534ec9a2f0225776316952ad018c793a5fbeddc21b6d8d1d1fa376ff8f5a9e95b9ed6219a7990356573e1c951b5dd479edb7c0bde36009d49a2773f642aa070a1584;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hde1bead32e5473922bb21a75ba419c2a3382d1123f80ba1e04408b3df94d71489184ffc11e92de1606825f7bd1e88ee05e3272ef169bb0bab517f7a52baf423e87401efd65667359b7cca4d63e1cbc0af5ed4394b5abdd33ff4eb57ae17a3d224766c7fad6771bfa3f2448c053169a5990d983841cd3c0cb2788afc69af6f29327aba51ed42168fe8a4aaeecaeb9f1188677bd7a7b7bbad56957b648bc9f6a13223dd4101658f724c53a51e08343f912c10362a359136c60c9a232acdf09c8f666338c6cf96d04fb1c7192d1fd9c242e5ebcf3363b0ed4baa9468019f61cde3bc88a36eb2021c6db4615d416affcc39ae43def24f8b7486a4c4b18d64cb6ddaea1ce6d0b92a0042cdd4999083691a5dc577bf856735377cb6c4ab784dd4f5aa68f5750a392b9d7ce9bb7aa050a35b316c9a1bb0c28ba658d88ccc9d5021fe6894800acc08dc202fc5fa93727b9ff111cb62f6a70f96ea37f3d3a4816297a7b9612b78dd29c094cb1099eb4960d8c43ccbe27c802fdb6ba19a04dbdbc6c1e5a51ece4ff458ab2bdcb99e605c2350d31f8580915c54900a5fae99a3b318a2a11085ed0b7bce86baddcbef3076a51171005576e80eec0ed0056ab0a9b00be3f709f09a5c861dd27e82b7b33f7e62f07b638237d9ce2571383d1293740f74f62ecc4a20a4e68176dfbce05b144c4f03ca39ad4a6571a80cd73f1388494278c4cab79501d648a0d4b4479077a3d2caf31894d6a78019249a8ca1bc7254a8919b2111e51a9f0967ebda3f2b09afcee7068bca31e541ecf79d723de235606c20928429e70ae569ec4b900043166b7d2c74f880d1aad3b78d08869309edc5443e677d146f9daabdbca6391be19300310b38861d1e7287469d1df1b2a042bdb195dbadf9302ce76f7cd3c03ee5ee8c38e1e73ce24a78be1fec8807c41c0c6a28ad3b0f0a13cabffb458dba65e81c385074d67eaedc8919c252a008625348b33000e631a62cee1e4e6700816f7bee30d193e48fe7d85217c587c0d0620d669a10f51d91bbb0a96cde19721240d8d38f0c9c7b064e10c8c2b0ea3ae803474c6bfe368cdccdb2ccbd332a95e3460b36f6fd15a5ecc64dd3432a89c9d839766cfe28a335f144922d609158f8b1cfbb54f77c68950cf0663d3888195202ed4a28c64552aa30ac6db735017567dc61da027a9cd7210376f710c86e074b688b96b7481b6f90a2b6a5d67b739be83da4f3e1736155b8fc5acc9cde20e18ef49c97d02caed98af623b4b11a3fbbf7f8aab02ae3a15dba10d204c0111d386e8255c6babcb007ccae20484653849bac15f982a83b7a9202c9d1a3d6b426ead47faff374f452311085b9583458613b1c29d01e59920f86fb497ee40cd8682d96272c5fa28b86a8ff31270a2737452cfb16c72b5e0164e21c6bd3df8bb4085b245e44889ef1aa71cef94c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4bac9b8d46290b9b785d7cb9db55946be7ed8815f5391ebddf979184351f36656909eef36f168e2b9da20edc4e2fcf3017b4bbae56d35b6d7443eb687ad5454b70b72e0ceb540b364afacc506c5d0bf9d2ddfb0e0cb0be9906c5318f5ea2421fd9f970f0993370380e8303aaf4a0eb9804f5c470647724579b29368894bf1e401f7aaa5f62919e7cc166dd5ec8b6bd4b60eceff021fc67051bdcb936df487840fc33a4be47a989a2e15ceac4136d8df0ab4d1be1a134a56efbbad0e8c3c72b234cdbdb29f583a25828a4430489a345752e1bb9883f9765a3f87f1a117d1fbf0fcec7a443df2972bd936849b704f2d45383a0faeea3c8d5a876d0bdd3447242a249c8f75b79e9d7d0fc410280d02c382c8b62da80b75829cfeb0ad077b4d11a77691a51e8fb0fa135535e210b66e6ace5f99a8fd6cb3ac285ab17cdf4594a039e7d7450d7087021fd5af8fe5b3f9d8848cdf90e47e56eebe7759b47525c6c7a638b5f68b0d7ebfd9992ef792e0336c1010cbb5ba638871ac1ca17fa273550a464e19b3874e755e298b9056de4b70d353248ed44c7fc406d25886521cb5c66ef620b8d47fbbd2f6b70d040cb3ff557d67c39586162125ae6f55008d8f88f742bf5747f61c048d66c9e70e73bc6b4bd103450491f9597144b837f887c6225aed30183cd383bd34ed983394f56db0f1d8b3f6a6f2df19328a46d08e3aa21a6e90050bb3e7001fe8bdff133bca0b70fd18b17573fd7e9178beafcbd3ef5c8fa3fcf039eef2a7cc98aa013701e1cdb37590fad9c5aea4c1eb1561c0c9d42db2000354aa2b8096839bf89fe703944d31cc5200aa7a520ea86850f98681f3671a2073b5549264acd325f81ec1926f2dba8ba5eefe1a68ddde3dab875972214e27fc5a1dd5b3efcc59216a08aceb14d0395917df3d9a20173d69828a61ac053533195e65aa0d5dbe33595b049652c6a31fcbb1c22e436ae7f3e5931723166af0f030acd87f30ae6c1bcb0dcc02f62c32a1e18dd762f26ac903001ef8acaf60cf7e630cb4f8b6918ff1ef01981e09ec2a17cfe362cdcb374f48a54ba687afa338f9426fc42067fa86ceca2e9705bb7a7f2d1f6945976ec31d4468a520316f31c94a1163dc26238a8f1d9310ad2914d9f2db760bf305e81378d5a4e073f5e09262c2fe24c70d94aaf3337a9af46d535516fb319e495df37e0db06c80920d4b6e34fd44a65eef0d33d552462e4b78a1c7f2459dc4b28a2abaf45d36836972dce43e5c07994afa877a01ac5ac3da62b091357e7de006a9d11fe0f58307c4dc51c1371ac5fe08482a90f573090f50103ae63dd564692bf9b0cc6cc92e98b2b67f17af800797ee2c7b2a1c7a7e840dd46fa8d777edbd5998e230dd0cab33fc5bae1f08eb5165776bcd9dce2a1b13ffa56d7d0ac1d2aa73ce59664e262e5e8a4599bea9203a7e159;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he8fe077b041fa2e9a7894b6e41738eed5d832339f0a68f61d5f00101a85921506f4be185b9d9aac340ad204b47e0b2ec71ee2ae0595f9e26468ac2164e50a742c19b749c9928c62ab24bf94d3c6f4848dd294f50333900338b718e11aafd3334026c1d5b138891a52b6c7ca921490d6cdfc8c542317a7cf4820320b3b44d6f2f2d54bfee26be5c93d1c345bd3146d2f1d68b43d6c66617be17e68d6eaeb9a120b827b8fd346c955a73594238772085ce5504ae635d481b025e356ff503258a722915e30cfdaee64c4c0070cef6d17f6a7b7b3ef00f7ce43b18d91d2da0de4a04f1c92308ec907d400a9b41c4cb700710da7333a364ab8d3efdd9d664cfe34260fdf2482067a6d457f7bcef10116e004742686228340e0ec86ad9757a0ab8a527f908088000c39358ad8accf66653775c880b1da621023b9162954e357ad6bcdb562bc841301c0ef3c47d5065ac48ad54c690e238fce7ab3dbb36c886ca9a2c63f8a57855a0a4b9d3e3679e59d513a0ce9f837c4b0c62f8acee1efc8796b5197d44e64c670b05151d11f26593b1865e9431746fa967cc4a1b1ce7d4eb2b5c05f92607c6de54b1404ca29fdb83c8bedf1dd18f70657af7f3b952cd1617a4bbdfb196fec36ae48d9d1ad03aaf3f110cb6e9a31e2800c4cc6c9454b5b2aeab8f772959e2701ea3bcac1f9f214c5b42b3dce4c4f8dc41caab255eac2ed0985a7f26489b67e42b4c9b46e69181ddfef8b28ff822302fa6d8d52701382d2dd2a6da7fdc91d3291c6ecc5ea3d110a2b6e31f900a93bf225a6ec343832caaa91ac4e62d4ef6dbea654d625264f3ea82047cebafd05d290c1b0c8960165a5ce193f824f1953f08a1107b78b34736d85e340ccd1855e946bb586556bdcb998f6ef1383cb4a2c21c1dcf652a42ad738f577f0cb2bb2bac17606e84ba1aa69e7114e98ab237405484a17eb1fe76309114d979b0483a7d81472a87ee85941b455c50f313a6389e50b0010a63be6b71a586eed6a492a729e355f2482b673de48869f8da0f48f2aa1de111012101b5c3f4221182fc4e3e8c012f883c83e04cee315324fc22616a63904fa4a31a2c85d77c4d6f5a4f580635c4b06d048a78e49d8f5627cfcda22e5cf3d9b5282d7b003ddcb089471a87373d1b52fd8ac80a580b24fea74150986a9063ee6b083e61f8feb0cd8fcac48ae45be8d473eb107bd606efafb2d451e56cf3121abfc84007f39414daf646784c7dbb9bddf4245f22c98a8ff45a5e4d28812ed485d3ab340e95583ccbebe35e918b96dbdd6831f09f606aaa04847db1757a7c0d52d9408b6a41522dd2e76cfee8feee68a417410bab0804299277cc4ee02a2006389662f20430f647586d90bc95b2bebd9656cfad07a22bdc58c943be4c9cdc4bede9b644e16cf5ebca6fff3f96425d789fb38949713317b40f320a23a91134;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h92759d0c9232e462e3257d142a445ff05d03f151ad9062db8f62a53765122e34ef422ce8b4074495aa5916ee9418e05d1247baa88cd260064b61d379d1c057a2244f274b117cb942f6ab8c11744e477f1cfa497f989e07e315867e343aacb90dabbf6cc35bee4b1f779cbfde859e047f0b1b4621b1f2714480d84d2cc47c8e82fc720a6afe1dc1c8c26bd8e6707c2c5fdc20439c30a9f36df1f40d8faaa340c840961ea53e6ebdb66ed2e5233a4e248bdade1684f2487c2fbe591505cf34154488a02222d4cf9807d5c401cfdc4310cb365cf1e05f5c4d7b585f7ed8ca39aadf002a1946ea259b78c59c3d926c44829b87a568feefee4cefb7176c2fa744da755f4a03bafe937114f7a7ade7acf40f0ff8d0b238b94760be9803cb7a290a17aa0ce1eade98c6ab2b42cb5dc760749037c023159aca1a06b0dbace6ba1456eba8b147b1d69747e0fd06c7630674f28b31567f6033923493aa6ce671faa21b799d59397fe0fba511ec70bcc81059a3554f2d78475b956b00aafc2a157b49d9359b162a71582b912bbd37034233a4cd9e7d3ff3bf0aff290ddb59f8cf29f00b2f87d552df922950ce40f0cafad12cd004221eb5ff6ed28a1dd106236aace288fd0d8476b7bed10d2f8f5b8120e5c7f23d45e9fdd1b34c449caadbd70bd7bb99941498d5f76f2e40454c108cd5ae753484e0514743bde53feae295fc76b5da439d6f791793c465e5addfe752d682fde0c5df88bffffffc5a2dd6c0947d75a6d16098bc754cbb7067481ba12069a8197f4ec6bb56929e4ce4c03c4cb508ed954bc8c1c7df095f3925440317f7d8b62872e250d3cfe37b3044a8c67a3a25b91d2f72852cd550e0497e3b255d99fb8d6665590a5b2362d053b8618246ee9a064cae73c196587eb44ead46f35fc57e4c78314a302c42b9c801ec9606ac7da571aeee95e54bb2ecaf1156a3686b4763a164d00e7ce11b11ef582ebe42efe4fd03fe85dc605f85cd5196b27570c1c394b825fd7848bda05382e1036b485fe9ac1a249efc23d4cd9f3f1a746c50a902dba392a58227638095af81cfd05a6fa2c58e9e0970c4e244cb9b09c25976a5b80ae2ab7165969c84c654ef33308f1fcc7a60d53a872133769ffb6eebb8949690828bbbb68904ef69cdfd58383f4e46f28aa49a50ee7f6ef0e335880eddc4370f784ea88f729bad06c4f89f42138e14a1ae9886cde7c3f9c2f152c23c5dc7f5d4e672476c15ce0391ad65a08e8897d0e4a1fa3e7e0c24142e4bda267cc868f9df202a87b52ffebe6547253eadb4f9ce31d58e1be6cbfd2433616b672b3bb9ef7c1d0cfb574efe6715e350567cf782c0a70a88e21a2d8e96ab42d84c1df1cb6f4ca637c3383d2513225595a6eec0e220318f99ac806ac83c19b78da7d5aa0344fcfd8c8a4f746c73dc84bf11be40aaf3f5c751a7f6dedb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bde1b6bf332334cc9899eeb810f1890edcbb3a94b828d98fc50caa9e31ff10578a87898a4e2da19bb35b4e3a8141fb3bc6e00653a1d7ea80d6accb0a7506bdf3560efcb7988c863b49e5ef4ceb8b410e9cc29d5e88ae5f6a04930780f575c2819750f3e75c36c1cf80bf80c10ebed7ed98284332c9ebef91e65758c0b51754a92120100e7d830825a68d7b519ba5dddd28b4ce28a02c26000bb579b564550b8f3b158655ddf60f0ac708a7c39ed7f2d1ecb81feb284e98d4cf2e26f15fb0c489c2563a21897be755e9f68ddd1ac4b405a79c56739340c16b09736dac7e5c5a0f67c7e505dd9cf7611c1cdffc2276c558a246bd4a903661a092697bfe0b56265a00f3e799667b6269e156082ef4a3ee7e4cf93f8bcbea1b8a0180bbd03dc1624900d07060e4f416d4762a35e09549951c31a17fc889253be107a420ae024f6fffe0f7973328d08e959ce514dd76c2cfbcdb734df8b4c4cecc16d9af84881e5f9547282461dcfc695cf03c5d8ed249d1bf17ecc92aab1ecf89e20fd853a0808550d8758ff77cacb714a461ae6441409c334d459a16f7c0b75eb1cdf07089981529bbcc0d701453365e9356547c46d9d4bd1587df81eb85b17e096e64df53c8445e8e8a8b51ae828f95c681e0baf8f3d04b1927cf51f6bdcf2535bfd4c6c8d56868d00f6f7c4edf7c53870587d9e548920a8f14a4a8832d07c7901ba982bf6bb7f17fd54108e28b02bf5f78a474ee66a4cfe58f0bbccfa3e59552d9e6da8ee85c07cb445bc0c1b7437cd8649740fc84f587d1354ba961031c03e636983c998992289c8730292c4c7899395d1a585780ac8824df09de69631def758841aa725f634e899990608e44e0885698d630138c72f47a60b6c0fd4eb19c184568dab8967251b92261c4cfc61a5726cd7788ab818f5071be7d36662bd31aad92367e9b9eaa7df4c2e1aec6462f97d5d5c973cdc2ff508bded547a515864ecc47b0b3ff31f112d712e6b8d47891bcbdfd1ec3f020a75d51fa5492d699a8dea1f4136c416cceeea27969d84a14a67cfc7222fff6371b57121cccc4a76dd1ad66693f954c67bea49a34391bdab07cf79808d263cd7abe7c38af253dc45b52e1f9a7d636f569230d8a57cee27736de5ea25ebae51038ec8a2ece49f7ed149ad59444fb60f4779fce83dc5d8f5949c02c4ebf49d4df244e9c773b39aecea7b5af94003ff828b372c93033ae2aa64a8f88b7ed8848988a680c61b8fb206ac7a69de7a9e67fb639004349efe67753a633975ca1858f6fe9ee972cae993cb1265e46cbc3471b30c04a682dde640e342b31237348d60221cd47582120c7ea6d6c9cea5b68d959c27c11a08b9a2d12b4d763983c9d24b2c2b58f7708f8d5066ab9e3c7966b6678addf724c7532b2e2c7073e534b9ec6154e19339ddaeb3ec41f077076ff119976c602486;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha18752ef67cc70dc220a189b189c58c36ae2ca75e212d91e30929b6b3a8b2c2be96002f82150d75e3807acfa36d46446ca08eb6fef06729c54bb017d4363851dc258aef9ee2825f586198dcdc0df442eb8828c58b3b570aec0d41bcfb9ccfe8b457150a0ec1a52690ace9f30c37bd504d5bf71d0f25f71f7bd13e952c1231eac5d79bc0e068486ff5c656aca55e18582a670a342b918c752e4c471d26904dd247eeb91c3def9da16d36f935870d9646466645ae4122029bf073b47f6d6b2c887607697507984b93e2d6fb446686c13afda8a281ccb0690345f30da92d9ac9910b00825fbdc8bfae566aa916ca46d858a118199338a344436d61a720ba320de908182d3f4fd786d0acb33111d53102ec551ee6a8c035e4ab7e14f22df54e207b36e33525fb37d91a88670cc4c3272b2317f830f48a529c62c15449c006ac86004cd272267743c657afba64c6236dd23803ff4a2bd5a3bd0877cbde8d66fdeec28386eaca3f00a2ca912b475e70bb7fed9a33038f98e69e537be923b5eace622d727de89cb3980c72cecb80cfdab9a1073e4d4b93d9f29e454f1cd2213fc96bd309d7014eec97c4f79faa355a8edc554de5c70ba0076d89af73cfe4d6871df81055ea0deed9b09a06821b9fad76f032ec1846ac344edddd2f12c985110238215066782065fefec4b18bd2016d05584c55371105ddda9eb8b59fdd70e8e52f4682a59cf7ee4040b36718e1bad459f51d42d57a644ea50fc46b0eb56241fd089e2261b55d67a86328888196c2455ccedf990a104a3f2522e5acdc4d308d2c18f3a6b21e84f2668721a9a21c2d74919676039b76e6cd65722216a9586e6dc6cbf2c0af9b045f8dbae8f3e7d2d7cd076e6f62068151f75f50e5bd67fdcce3103bb463a5d5b01d419969db9b639197727ce6e8a21ec7c8d97677f063c9fa1d52202172c8d04d6e9388d5452aa2dbadde56f87ce6767ad4ef74cb49bc3119aba415dc919129367301bef04d317185bfd365b3a6c3b3b9fca6f0752c0c7ce7f391fb3fae4748af70933e2773ffbb71114378eaf1c702df9cfffdd11998d0dd094aeba913be1e6578d1928cd49207545a6e5c6a0087c79a633d079260431a6519eb144fa80da9f6c8bb37dc7a84b4efdf4da268c6f6cc39a96e1670f97bba9192165c115a634f33b776933b45e9030c0bb09ca866cfff48a9f45bd4a887c5f26d5be53f555295c1e42ff5d7ff2cedb4f30ab0c611ca37472a2c6ce537db33dcac3676be8bb44cd6c330fad662d40bc3e86309d235cfd0d7008d88b2bcd39c66b27c89d03c204a27441f1d93771b0e0a2b492d2ddd11a297be42d721e8411357a239ad3c0c968e82bc400410576b257cecfbf107cfc87cc6ec7a36191912aad53eea09d21dcae4aa127a1f0f369096b1ade97f4ab4468120f77e108c54fbad902dc19b4824a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7156cd1f3d2b542aea8651415a019111c2b0e60362ebca94597687fb0b3a91883c4fb893d2e1b41637032f8a7b275ba7ac71212e60109b96a490e7838d587d90bed93c9d419148c22e61bbc7031152c9661a775286c41178a1cc3b409df7286c9dadeb43010bbd76b3c0415ab030fb9266f2d6a7cf7a283205107ed4d04af9b62975b045ea88841625c09dd6f24c26b0c150fa16b9088580e63fae0abfb91632a274ab9b661f12f09aad304fc68a1dac6c665633e9f460baf3454f33bccd177bf7d8876644d20d2c08c20ad16830397cbc5aa9d80c4bd0cb7691a60257afe9fea5eb175b4d4915703e560e81a39cb0bc88b2114d313961aea167e1aec137e1b3ded36b08ee3cb8399a3aa6ceb4d20bead69c2caafcab03fe2b8deeef133803c40b98a3e2f4fe2f7b97c3e028adfcf05b4788dc8977ff8d76bf3b26d032eb7e3bc03b378267bde2e7fa346f14f5e7d25075c41262f0fb2330b7d20f41c61aa3a7ab701b7d6c665ed70280398731db518f25d79081967738334eedacde38ef0b550cb6aba432d08c022e4964dfcdc34746a7de3568b89e5878e05bec11899daa39430c5f89669d91c4484d879aa0c37ed002ee45461576e7669a6713d039f35485a0ff8287fa94349fca6e6ad470927c761fe94fce039196f39d5525e464c1423429c92003121ad55568de3148e9f5cd9110c0790caa10d6e8b45c81578c197024f3edf7e931a3ddcf3dd7cbe873f33c17b1c94887cdd886a9aea28afbf571c3a7152dc334b4b0de5602373ad4533cf822c71b6bf4ad59fdf26b76f4813c1a7ef4ad178d8eb1f6ab25c595d7978a36a6917c5f903d117133b0fde4b871065c53e5c022d32d610fb69e7cd9bc0503248904bcc835da558d9144b8de0452d5990925074e4fd26a4fd84c75d70d81e8eef7b6af0c87fdda9262a23c4d661726baf66af364091e472622dd714c0ecaa01a311876c308d817cea9319b1d48ffdc1c120aee7dedde749a8e6d295a1c2ca4ae4f63de662465e980d8f0dd235c7631b4ae053c18aa2d008770594bfd2bb4d046169d4bdaed8311ab4d9df578d75246aff3e1ecca83a23bd5db445040d8d56a25880a342461e4b264fe31ddb5d8b5038bde2e18847adb2e7f58e40ccbc83a681963776b42860aaff27b181dd1789092044eedeadf09f915c1da524404a8876b66306327b17f78dff95203e5fc3880b63359ca2fb009c70e4fea76b80e2f9e530a514a77c128e8b85e9bbe08777d52da7d69e386d55bbf9c2d62ae4ae597c5300aeea86a91552fee8fc27a487a806d20fbe00d7f2b38f87ef0a193f6651f390e7df415eb654fa51f3952f78096f21df268c35002b6fbf3d9269c7792ec1ef156d4becf230941109b6cad0f3301ef46fa5c6273a49c1b06a7ef4a3d7b738cc5db35072b41c547e98fbda447575cf69772d71365;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bec7c72e87fdc6f8b6156704b601d2927beb45ff59b0b904e41ad611f7ff7a076b02bc34401e92ac5be2cea1b2cc377419b894bad84dabe6271942a8ef56b8c9216f295975ff4ea40186fadfda9b0c9adaaa1b224915deaea96051fbee14a0194e42f35e9d0822b0674935dffe07f944bfec2f8ce87dbad9f2c66b394d1c0e74c9f161229e6645dbf8919d5f5ed5aa1f3d953e77c7ae2340db9dc76b2055566da731d69867c70c06a48fc2f56dd6f1c3b61268e7fa8fd9285e1bc80c7f1670e471acf92252c9e5ae8b5d8a10038a333178d532c9d5ed42597e8206ac01010cd7453687c5c5d3adde5d468afef84f6ac92a7fe51c92c40065fce74a5b943faf0f48ad6180f3454e3ed75f3e15d948a38bd2665fed4a84e181ef1663a112fbdc01f40f1a18f01976fc41e81af532f1aee5e23b87862deae5e4d012beceb9a6790fd04233818f1aab975d4bf81321e19c8a1e15d4db4ddf120cef19f676a1fff89f48abdb2387ddf99922a94092808dcec8e80aa60f08a30560080df149f1ed5b2204340d55c0e774d088b913c5f8203c1d22f88a058166dd84c9427dced1b7d0355932ca8abfe8526c66f84543ed03bca92240555155bcf8b54569384835960052d56bae184c60ff31837819dd8ebdfed6d9f7e33e73633709e582ca11211da167fbcc6ea2bf373f1c898f1b2b3c2cf2a3fe57ad6fbffd80348f8db4113b89cb188565950385b0245bc5338993ef502f3cc039732e5b67d7c6c511590d067cc6887830a962642cbdd3097d4392518a4bdda8bcd43cabfb43094c3bfc546882d24ff184168a78e91aa4eb52e0dac2943ab9a506841a06b4850d289dc8140b85f25c3a40275f63f8798005e5cb74eacbb0a6b4ba5156c4ec87962abec0721407cab8520ccae0a98b2e0a646a34fddf884baf89fc0edc5826bbc5d609e030572e737989c6d5cde387cae9d25dcfd954d9cee15092788b6654ef66b06b0a9984bf41beb25cc21c1b177a148856ebb77094558b354ad693883d9848e7972b5161e8a22b7bde78fd2290efa3727e3038df1683969e2c2637891914edf746bf724b0acc0641c56115f6602808443a315928f047a737e366736cda2200f2bc6158513efdbded70e4b665e355bb021fd9cc506495c177e4a038bfcdbd63aa5956e277fae7307ea5e791b1c73c857367e75a3ee8ff2b7415cdb31ff9ca5fde1cf70b83b562e122987f40218fd46e56bb10bb27fb140194c2518c5acdd711f1a6c35bb00fb1743a90cd65ae0c8862abed4e32feb4559e45851a1c0206998e35bbdf8351c0c8672845de35fcaae70b7556fcc51be20d5ad7c2a195b36a3d828898ef3a3bb7c1fc00f54bab460c8484e6de1674b8168a98978bd71fe715e4007afe92a89f930192f4a3ce2a320a41b2b2f2f289143f99a50391439e00ada40d87556e616a95595;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3be63764c6f3fee5b08d361e93da2ba61b26ee1283ebf0f80482b3f60c2fdd9ec56bf0c8b108018212a42b23207a302f48db54ccf18a3512d3fbcd72f94dae5e56c7588ac276293e7aca622947875e15db61e9dff8a8526d7e0af027a5f56c1423027e01350b0f6f4ed9961581ea0657410879302d004d98512f8ca4b720c8c73f82249f34b64bd71e67c5f76e17e0c941d64bc313cb88b23fd45623f75802d55305bd4d69f50ad06eaeadf9a4dcfd94721397a50744c64006e4e9283a977dbc8fdd05c94aa4efe2110a5152914109568f1ae76dff43aa28f1720b6473815805c8066bff96e9aacad222f38052a0c9930ccd3f51a5ce0d6c9b2329a9360a0085f0472e4dc992c755039ee04e50a878cba363bd695f36827ec772cf5f1792e873e5ad94c047d83dd33856e2a76039772be252ce82ac5af3f1c507ecc0002ddf71ac2212698e4c098a2ef3b18b7f99a2929323a8baba106a603f2cb2936d1ed3082463247e89ab0cbbbd1b1850d2c30fe5be3c3c77ece444b8de9673549702b2827b739ef193f3ab678c3bd349a6b69f97ac3c28ef5e8a7be5d5aa793c08bcd2aa6a1c68bdf765f104274954a8cfb9f479668ec15cbad4605c950c3a89baba7d3b43d91794d9db46d4a60b8a673ffc81f38cac9f97239a127622868b85829873cf6c829e1ae876434a650181b03d575b600ee4788bebd4e9e84fcbc21faa01d2081f78a7998cd1141b2ad380b039c9a5ac01be5f9823ddc3a1aefe4b6365cdc0d1ac2775e98dd7088c4236f8390ec70ead7365ba39cb615893e7e0e6fa20618d11d29351b2398e77e501035fea88ff7a62c6931693c63585d9664fbd0fc174ea36f4540c05e2dc6f93e7a9652001c2ba0889c2fe385a44c8f839ba02597a6360090bda8c4c8fcc1c64f1201631173e06e592906d8112702831fa224a82f8ba49589ea31c0f0637b102e18b9e172210e143fe0875bf9131746be6988dbd91b383a0b2911cccde4f17549f180672c540dd333b660db9670b6e8e03dd990e7f130f5947a3e1f04ab4d3ba5671869ffdba21ee17a30b57e06e260b8068cbefa071f878814128592cad84840edeb6a7c0a1f38c8879cc4af426342fbc605558f4b75118ff65b4dfb2fb526348e680be0dc44a1ba5a83976a5cd92c877b1ff96a249d6f344e4f676ad4b3aabc08f6cb11b4895b339a612524e4978a6a87e4874d547f07d7478729e06c5a234cde57f1989d48bb11d19890263bc1b42e089629d3a1b303f05e828bb8eab01ffd3cacb992ffb0a2347b56a6e8f6603a8087c52f2b36af4ea2f7dd378310b5e84978ab40284386e79344a3d4e853e7715181ded561fccf0c1ec8f6fdf4d74283ca1320f31897b17a4f9550435f25ed012cef9d387b2f7c55cf9425de8176d8e94050ac8e073929adb572208a36eaa104eb9ce424dc3915d24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd5c7b19acf9b072b933ae69537941586cdb31547204a5c882e280b17f61ad0b313a71a3ee21fede8ce6eae32fa4e904398e991401fd34f2360935ef741450f8da954c5e5bee92a7a6dfbe8c8979053868ce4dee8fe528e7528506f23fb7c03e26d064d6312c43d165b463f388dd0b181cb2be16c35c86c26acd45f3648e1d9d1fa8bc447eade28c99d3c110a36681f2fcfb9a2fb6f2aff039e121110f35cf70af761fcc831eff7dd6e033c026ecbe97ff8c90112704cf30157131d788b9253952f7e1ebe95f530c25e0d7845a6a5c0130ae3b3333899130671b155843f2209f0631dcc5481d7acb5d87bc36e6526a522787650509ca88caeb77acb89b0cced69bb6bbf2b0b614ed33c07d8357d04d33ee916d52b6ab94a084c5abc33cb60fd2be3bd657cb1298f618065ccc06a41a35fa8500bba5348e46ce72dbf9a4b78b6e91f3b9b8a8fa5dddb4d5e42f5428d3ceb35a75deee2894bc6fed4022721fee1481cab2845271dbc4905655b4c6004b15b428b1b0671c747d762031f90e47e92bda4a50bd45f6a10274d3c35e4127717ec0102d70a90a037f1c81bd328e30d034877f930c9445bd594e368c9dfc41761085b4a77b48efee1b08a50e709c4f795e0a676be5fb9da9f1694727044b23980c02bf4476a245a54490e0f5f83c08188200461cae5a311a4c88d55138013ef8eb22cd928a5efbaaaa5e41dce13f396da043d5230098082ff94b610d32b1a25aa9286138f4716a9da0e3b4c4c65153b82dbc8f5ac1022085124ec51911765bafe5cc29a4089fc39f2a260a0095834f434c759f2c8a194184f8b9ef3e60f30a778095599180e7c9f1bdebd7aa8dc073ea631bdf107cecef7be62cdbbcc74b4c8855ef8f7c13b91a7bf65f4265a86a62db7c02fae06cb380e758e893c4416543cb39efb0ed7f5c61fb2ce5f65cd196d1f5939baa40a72ffa39f8cfc81179bab0fb71a3e5682d0cbb5388315a3959baf0038ba798cba340c12250972f67af9f18ad7571ba3831dc8a6c62e0b8e5e9d46761460ea83c17353b1153d6c430335b81fae224af8277731bee2b5c7986e41f90f76ef837a0c2b8c45983a9c05c75f0b6fb0437c896e3c135aa615487165f43d375ad82dad8a89562b1107a9f6e0e020fc079b8330ca97030980fd10958248f1a733cecbb0b3df4ebe4af428713f2bbe05463d71796401ff872ff78cc8188706b3aeb805f319ec6239d6cbd3921349e05fd00a66eb2687e6815ba1f4bdfb16e53a10aa23954ce868867ca2af425e7d897d6f598d8882410d6b6cf60a1848dcf49b0fc6678560978775f190cf47b58e4996206b62ff4422bfc93c37a7374d72c93a02382b8a3799cac5cefb1f4bc7fbca4bd5a5802d0d1e288ff56455665f5948d80e2706e01eb5f3b3517f933c5ea0ee21fb17fdd42cfdec29088b64fe37c904d7146c;
        #1
        $finish();
    end
endmodule
