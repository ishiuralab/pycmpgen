module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [31:0] src31;
    reg [30:0] src32;
    reg [29:0] src33;
    reg [28:0] src34;
    reg [27:0] src35;
    reg [26:0] src36;
    reg [25:0] src37;
    reg [24:0] src38;
    reg [23:0] src39;
    reg [22:0] src40;
    reg [21:0] src41;
    reg [20:0] src42;
    reg [19:0] src43;
    reg [18:0] src44;
    reg [17:0] src45;
    reg [16:0] src46;
    reg [15:0] src47;
    reg [14:0] src48;
    reg [13:0] src49;
    reg [12:0] src50;
    reg [11:0] src51;
    reg [10:0] src52;
    reg [9:0] src53;
    reg [8:0] src54;
    reg [7:0] src55;
    reg [6:0] src56;
    reg [5:0] src57;
    reg [4:0] src58;
    reg [3:0] src59;
    reg [2:0] src60;
    reg [1:0] src61;
    reg [0:0] src62;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [63:0] srcsum;
    wire [63:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3])<<59) + ((src60[0] + src60[1] + src60[2])<<60) + ((src61[0] + src61[1])<<61) + ((src62[0])<<62);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd105046a80d30125e485ce59d0cf7eca296b09045860dbc8e13c8db95c5fbc5d34663bcaa9f2a75435e5718359faab2122168d20b1c82d832e6ccf0b98237401b53d3ec3849e4066e6ba6efa647516d32b8947f6b5c4789ad6386595453896945b415ee7cb2e8640f20c25dbe172324d990865ad1e00d0bda0b6a1eecc81f769;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he911d817198427b8ba17d69c5e19c9a758ff60b3fe8b4eeb260f62271407c333d597032c84bb425478fd89060edd8f2148abbdf433b342a711a81f8f91828c12d65c498b6c7c3d655c1f0a61b33a38c453deaae13b5b5d475576fef0a0277c7e05a2244157c32c27e7fcbc0fd2f0d9202b37bb8ca2424f0c20dcd38f5b2c51c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b5190cf015869b3f2d89b459e4abb29c6b37e1950196b5693fa8bcdc05cd37aa01f9de0712a62a6349ee1ded24634e61bba2062f372193d70f9bbad7d1c8ed0ccec2884aef1c194b9f311a2300ef68c16bd51b183e63096116194faa589dc5e7685ab132bb68b6ab426f7234276f3cff4dcd16a2b86b2eafbee44325ad412bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64c9773595138897ea5806dc868a204661ac2c56c73ccec5032e1349dbba68b5f0df6d5de6894fe5d473dee597a8c59c943f9e1bdc048db5db78cfd276719c86e6afa8cae1633da650ea0edd52cfeb637a218634ccb9f5b4efdd6623ac8fa4c5de6cffe5fab5715ef2aeb1caf8fcf46b991040f075fa733ac8cacdb8902b010f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h132b171fdd9197927624191aa461bbc6d690bc7404c1cf446b66892e0cfbb58456fa8d10e0a5b23f5f7f6cba444a2b70787586c466ea14c589963fdc5865b1d5e31019e3eea83a7ab1670fa78263b88147e6e2cac5d5ef2dbe19bdee0fd56a3e39cd6ca0d69a930b780e9f5195882899ea9be719b9201bb24b17377915aeb212;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb95685bd2f353ae956b42b38333e906a34520ffb2d3496ef5dfd18c0811277fbd20a32b58ae3bb2c0414fcaa2837bda08366eae932fda77c099e7728c38e4611cdf7fffce94542c50dab7c9e1486a6d3ab377d5758e42878c9dab93252daa8cd48cb4937540e1010710bf68cd3c8206582064fb69b4f3392ee77945055fa254a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf998d1787146e86ea0e18406a9a2375b5cb63d9fe4fc212af238655b5a7bb0ab39b832b1286c794eff0f179579c0a30922483bfaf58f915ae7f31a7f855c194cd4ab075ff6f6b1c5918a03546f14fb83a9908c754ef5842fbca82cf5718a9a23bf554e5e38023e18b60baf4a959d466016bd0f861d558824f863ffd98bb3485;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5c5073a3646cc4c666f01aebf2563ba889fde9b24e1672ae0d38271553b5364124c9bbe32e5d5d97aa13b78cb5ee4a58247d1ed557abc62978f9aa26d8ebcdd7d09cef635e5157da7cada1931f35587981be4c5b663876bb4a38544439001b1bf31691cc363746a96a4ac3491f964bf64658109746d24dc6d62a44f470a86a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66daa4c1761e46bbc92982a18bdc503c95acb3fb28925462b37a5ce1b30f3d721d2bb4e0f37a23cb75c9a5d3eb20429f48ea2ffc274932eb528483dcb48611ccbf2fc8c124c5477aa3f25e2ad1807d079ce377185d51394d9772c835ab3a787eb939ac788a8097230d1e5f66957313ae2a7433fb10384b3ffd5f0fffb0cd4963;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55a427539177b8cc711d16d5af3d0721122b579762e89e911fa86dbe4f7c812643f7fa415d1532e7c6b44157eb21b63032cf65e3cca27c3c18c5e461e38fe6803d50dd8078025f51736cda2259452d16c53b42427e9d6b3e0f17d7ab0382304ba0e2ff46ea1fbb6a92afcf6247d2bef9f065b6ff0c6c4e2d3ca89ec3105c9851;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9b66c4c4ee7a81f73b82028353b898e3aac8026a8ce157d8e57904c5148d775f2ebcca47e60d68ad2700752e5607ed1f4598e02db53ac13dae27ae9ebb88c817269da13bbd1f8703ff63cfb9840af9d930d841dda5e6c69e01fa8018a5855ee0548c92434432e473fd66b21afc8131bd65d070ff55e97da31eb2c8db7a28ff8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ff06f243e372f6cb4c247fcfb348937498770e17d33a22c21ab21575c3558f36e5f29e6436c200e9f237bda390281d6c79d7c1c7309db6e889a39ba85808ebee9537ab3a103724b0b0b942b2638f82cc3c60b751bf19b3f7848428efdcd70c88c23a42234284ca9b9105f62bd0be8702ddf0a00cd47d8e66565ecbb2189a6a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc74b2e5ece46e4e86c2d4d5ca2451bf8a9ed3f2ffb04bca6e2640e283cd66a93e2a37b7ee4d8a91f9595944b85705baee6d434c167da61e55c68a4248e37ed845900075deb8ab8acf13f470afdfdc91ea61dc9e53b0e7326004d8c732fd2d9b9d2bb05c8e1ecc514f495d942488e591e61fa6ca64f4816132de25e5e81d7935;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bdadab5ee1ccfe5a824eb9dd858183d6e1124ebed3249ac51c79834fdd653ab92d9f9e53ce68110b6bc41c3dd618fdf816822bf809708119e938c5062e89fdc9447b1ea5e76940a8e17b0c8e7b3154695a894ac6f92c8d3beecd744aa622090c11ca80406a636809d1d07029efbf6f58ed4800978199d1c4757c541a9fa4ca2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d780e0973d56fb1ed6655cb2dfff8649550ffb7517e9405c157037beb20d97714b4a950e29b2b16bf32d3b55285a5c62d1a59275cf3e115a7c25adbbae7ee481899600d444c558679edd9f2569eebd8b5af603181c7cec45802d371a1ea8783b4a8f6cca1c37c2ffec44f8874b179731b2852a9e34f0c97e6bd8e991a8e9b92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37fcfd51e40dd61677a8df4d16eef5f31e5e97f240ace158bd288ac54abf370ee2d897c8dbf3adcd2c3ae82cff411631bf18e6251d154b134aedacf7d1902964c2981445cc357180c603b432df3c4aa19f3a8129f7112bccec796f0d2338015c882e038b1b0e6129270641ffbac1d6bf735a8277816cd2f8835e9516ec1526f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91f7628808d2e7e5fd35ff042178ed6f6b604d7ef53529c8f11389c39f849333a7d1c5c57014dd6cc88a874c829be7ed96530b5889a618f0034f5f1e8bad389cdc694508d485048b71e6186d506d786bf051f87c928f2a3610b5631c05b4ddfa537554ba316d16d51c81e7a05d28b5e16a37c0eff3f3850c1fd7f37772a0a88a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f25095dae16ec2032142179ba444ef253da778a77ed7c4023fae957b55b0711d6ff8392f357ae97170d295ccd4ea10b2d819a2cf65b4901c5c1866d4771b28eead75edd208947665b411dcaf6a3dcbeeff698243ee3a0b61b95fcf362c13021d41b384c4e5b413decc218df8551fad44a96fca6518299fa6d43499c901e1497;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h585d698b16aa02c81d63a9886b98a34672fef1082eadfcc0690d1b96b3fda0f04db08d2b5a23e93aa8863ce9dba35fee6036f8f614652a7b042d60d3c8e85563f475561c1c31b1aa5590009a11642fbb7df7973a345536ecb5c6116480d1077b62494518ae6edd17b4db41e15b2d6ed2847b8dce65276e1c0ab06ef7440f6833;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha505b0f9e6029cf5f8507c47c0bdf5b6c175d73843dad665deba998906fe0e48b2054c63247b62ae552733b8870306e75f66dfb8122ea8b88ed40bdc7252a418120becc949d6c0c99a2ab6168b983068f9feeb5125f30f4538f9c75c811d834bc1d90875cbe6ba49e129d38f0a4c7d7b2e511ce99ac368eeaac15cd978f4dd9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he888801af02e74b79690970449c9f5c7876c4c02469eae029e69fab71a1ba86e9912cae1d77e3e3e8d531c55099370e613b74cec75f517e28c894a01f8657ccf0b29ffc48bb685563067ee86757adecab01f5d8cfe0e300fe3c729efefd06e99f09ea54840e13621c217748ea5ee569581a3824a342aab31c54c01d0baadb062;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h719e0b17c36006983fa621566c62c3cb3f14a57c5e1998d4ad3654b29ac16d24250aa0fc8f018752534fecd8b0807a502b0b31fd862f065a88564b1d30fd4772d611fa0b36777d6032d705a3bc7f6a2920ba0fd5da7a0dfd8f95e52f16afeb510c3022c016e7a061615afa444941de0203b8d671d402ab9d540a08c63754dad5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf833ce320f9d93039cf723a8523c89485b705b64de23069be1efa25b83ce0885c439324aa49ed803159f44228798a8ffc2ccf671d3fe144429aea0f8be6157cf96314a9e46c5e9cbc945a83da54535b63c91259b442d3bdca809c980d79e41c3442795aacf9421db51175a3dfee97efaa8ca08b2d7373b54c00be38d198c8701;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b2fa94d64a394c6d9af21b9d9258ef8c343f34b11f62f6d01a03be421f1571b4ec1fdd9595026942665541f186b16a15eadc8812dae4eebf5b99343c27d7d45f87ba3c13ee25ec07c1f2445d1c1ba1a3ed8d9da1234feae0cd9c95297afb3de6ada75348cfc2965c901649b00da575436a9cc24209323838a9b6c694778c563;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadb230751b310a02bf3d6dab44e0272474295badcd4197da402356249d3242f2af8af029f1bc620d8ce34fc0063e908be2099b032fd1dbf7bda2ee726c0281c0234ada956c655a2a7803b92e01a8d0eee73dfcf19454f5ee5b9564e39a2dd1c33fe642b1a2f298db3fe547fab24da22009008605011f3ba3599908a2a0ddeceb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33cf77db10200d4668bcc9dc9796565e2153ad1044c69ee3ea2fc5d1a096570a32a2fb21f5e6cbfc14185a8c8a1a24e64266b03f5c162ed67d0f03c7308be9c0db0f735ff019ffbf161144bdc6e1dce7841097e1949ab228eea9964d4a5095d813e019132d478351da895366a44bec1d9e02bcbb5ce75b9a8e621c31fdea3cc2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4ec54d8b34662e7f039b7d7919ae664fb3eaff6c6ee1c2fe4b08e9ea8583b93112f46c3bf64f55cd4a159e7aab23cc78ab1d6db64439bcedd03f9675fa225d05e92ce39eaeda391b6c7715133f355b7c610ce2d5d500d74d18f0018bad383f276597239d542b0049cf71249cfe3205be8fae8c1154d21f29eaf76c6cd64f572;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42ff943cc25926fb3d6da64770a667a250ef8ea2e391007ac9040250eb0efc3bbc2117df668078a1c93ae144dfd7350d5206157820edf3d6a7275d40f166949766c3d3819c5dcde8cd8a428678bf32c941464a1f270370f41b2b564f84a4552e5e2ec0c69e58f38fa228e84505850f0f66bb46c392939b28150ae105e2a334c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e39512bd55ece15a0c6307611c74a0a3e989a2d577f8c23bf0e109742c27abd1746ca36adf1cbad641cec2ed5769bd956f97a874bb279f7a746313e1f15bdbe93fa5f383b957f0c20598196d6ff85c0ef7e0d66f58626fe2a6f1d1487beeeb108aa851fcfa47539a72c7f0178a14c1277753e57a6c7bfee0621f808e964055;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe33b1b90ffe9f5a37a7c1afe13128ebd5568b4163e893d48c05b058e7bf973e97551c1856e6b7a409483906978f5947b4afe82f183de87166386ace57cb1ab1131f0561cee4053eec6e05564add2fbf2f0e80a990a041b4e30e8769284f787c66121b1f492ad6485305cde37a779050a49ff772d9cf36cbb6e84f5a4f805204;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7be0c2e1d50c19ea02fc17fd97393bea7619f03088fe655799fe09bf35f4a4ac8dbed0fa65bdf720b330c9e175c7e3806caaf3f9fc71b829530d5285de0c6d60d7e045cf9dde2526a60d3bf5fcfd99ec59e2a5ab53fa92c90abe7f897dc342f132ef0b1715ec799dae3e07b2603ae6be65ed43a36a262891d3ab5612d468b587;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h777aa2cb8d1c3d77cedc1cfb2457fdd2de9f89d5f0dac36d6ff0334e98aba4aa691322f044baba6546f9712bb8a7af07a872592fd597f5f12ef120d7b636769e37578bfdd89daa91c9ebcce681d4501ad4ad934c07a57d9d11c3d5e837151b47c384c674ab4cfe2051fc9de1f1b44bed6ebf4d4f22238851bfdd287901264a2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ee1e15e5cbd9bcff5f92ee7e5507ab5240f69761f15e04a2d4d2c944ed6b53804e03ff52c2def94d9ad1c8ee3040bda5d619f04432127575998e99f4ead618feb41dbc2ed3fc82a48faeb7001193f4327eeb00727a59e4a3f8c734d77a6695d7247b22c23b624b6667594ed7c2dd0ec65597fb4dd754baf11f88b6778712ad6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd77453ebc0371603080649708272955c17756a2dcf33b77bb4fb43288a2193b12aee96dfce8401d4a487d99e565b08045311b9a58bc9ebf8f8033e12ab1a1b3b3e073328535d14dc5b73a4e7afcaa6157d3f9af0bd4fa522fdf81941fb125dfb12779a6c8a330823a480a475e958db7ea2159107bf482a694e87b76756b5d71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90ac8d3e9e072ec98af44e548d4e8d77cac7dbb8dc1797b1e37dd96420379e7db7b1163e5f174fe34756f37d8fc0444062191eaa425244d4c9f2a1f14010afcf3e82098c455b1c655e38288912f8ca6ecd799328b3cc9f1ffccf42c2dab6a51e09752bc4af1b2e4db0baaca4bc16e8a078d12e0d8399e40a6119bc4ee124325d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb2bc2a9f0813f88585f6ebe6a706cd80eb3c518ff72302df232727486e0ae46020d4e4af3cd267b5bdd63b1a465cc3fa063460abd834032889635e13fbf3b2f05302e2ba0f4bb95eec5eed096717f5c2b4609389a878ae506a3b7e57b3151bcf5a6a04692740c98761cb02cae3ffc1ce8906e3a27648d5e096ac033eb5ed724;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74778811b43f1827c9ce44ac48f8ee7ff91b1c0602897a6cf1cbfa475917f973fa1ca15eae4986fee4d23d0da7ae2174cbea0dd5a0feb7f2d7e3850f252b77ce36d48d9a4b2d5bebc49218939cfa26e8d597807b9def99ad10124cea926d4ea1ac35bd1c39f3a4876338274578eccc3ffc70100d1903dc566369c1119f57c8f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha39c13950008e9a9a6749a03c07b7548bd31ff02d75ffbaa2961f0d4137db3fb2553460774c8f043cfa3c2b313ea34b6999fb29c7633fcfa607460c1ec9b7f79020681ec5a6e45381abe689d86c95fe6ab727911fff06658ae76ac49859d21727113ec77e14d4d4f5d7559b0497c649073cac2bd73e2425885be5ec109a94251;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f1248d4bc400e37f56071cce9e0c46f1df09087f2a4f1cc0fc56ce38fdbdfae2dd90837b5b9aaf2a58c86d70335105525e819d0d3f3e6ee577577edd596073c5083154eedb0012fde36f79256e3509b98fbdb6dec8c6f5fdfaeae4fbe2ebadc04918c7c154671e93bafae61ebc8bf41a4b855c5f6518687764fba42a271b36a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d7401d9eb3c7bcfb4d6329a7cf2bcbb0c043cabe426e37a3ed0e7de95c21f969541c02aa9b0ac706abe44d756656b47d7ef9c180aff29b40913114954826af2a2b9ac403fdbdec32509efa242ebc2eb256297249c24524ae68d907fa3aaccf0258012aaa8a91e1a3d8a1396c92dade1e933b1510d2cd12356ccc69bd2419155;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd742481c7716480572548a32a2dd2ae9376da1b353af05f5a85f6a1add598a48ba54c20a736f7f1796ae0d8830b3af27f7905bd93eaea370cfab1f758a41f1109dc8583440ab8e4101356236c75fe785d5d5c94601812db0f98de60dd9714f01aaebde9d00169816315f2cec70076b94aae7003204b3aab6aeb18548872dc58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf41ad1a5741a4c525939275dd7c20398ecac58aa27c3e375e649abd7fbd1ef563b30f4871c34159f8b9d1bca65cdf57ab811bb349f575979e11bbcf7414cfd2aa5c468a001f3746a936bb2109ba85b4bbdf70422e56164f7335511791f025981c67be0bffc6a926a0cec436f908e1fc9c66065576cb011b6df8cbb14fae44bcb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33986153e79d07e0e10b09e3afe783a5a47197820e5c26977424da067589bc78c1f5abff1537249edc1887f69a767378c0c40aee3468ca2f0437155f6132daaf826f1b45d914f5b407fc793c4663a95422a7ca9561e8a9e5b716d0aaa3c603ea0225def0bdd7642e6662d8cd3038a11d0fd22e62f69c3a02abfe6e2b5a17a4bc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f722f93c7fe4e2a13fbc6f699c9337fa85c0a86f2e8906aae95a2ed14fe279b93ce1e1c4f78b46fc6a8fe0c87416d41b97ff46283f5edab5d9f9bf378c7e3483dc92e60d9b37dbabf6838c53ea380220abb2cb5745cc5b2417ae61099fab82266962ff7a3255fe81d203c49fb2aa34e2023fa3156e7d7632732fff078ba00a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6838e8480bb97b87ce62aee5a3f347ca4cdbc48c91350cebd6f8b0f14906c98c680bfee6908267277b6f45f2ff9334744a412cfe629ceb901a06f24aeab4a9884a6353e9e4d6d00643a23c6adbee25591642c5eb797e0f38c65163a5e6558a14c116e983654c77f8f78860a79045d4454d9cff1ca4eeb4f4e58026f76d7ca50;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79cf42c34c32a1e0473abd2b108f29501d1434c330caad65fb324e39e86f1b40bbd4b4b5d3e9ddb9aa596ca8b436e346bd3823fb29cbd6a3db25dce9e181f8f5610941d3d938ce46ad0441e0c87b475a4661477176d684505b81e62bc13ccb17efeda300d0caa4f7fcab6084c0355f321f2f126cca534e7d9d885c1ecfc4bf39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2608fec84ad6498fa9a45e1c0b9d01b9018e85b529254e9cffee6d554b76c921c035b39fad0ba85ebf0f99339822e7c453205fa3c3a0b6fe3314b3b1f6081748e7bb1c65917ed78761443f343d253e745e52e69daf85657cb0b407a170dfc361eaf50c203ac429aa07d8a86bc2b62196aa9330359426ca9d4e4fdc93ee9490f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha956ee5eac699ef52805b1b21f4bcab6bd20471bf791237bb0cb9de9b090dc10b20bbfa410ba3fd6e456a733b718d360ad6a1bdfaa1dbee3678cd228058d1450428d088b7ee7c3d9db3cbeb1068fdc01143912ec54efc674b8018c45498b575e9da01c96c7558f89236cd9b5d7322b555e1bab4524cd393dd41088fc9f7a714e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52f2865a1eaaa6d11676e45f3eb9ffe89299b42af624bafd7c382069d5bce6f27c7982ae26626596644b79a0e64ec7dd659112e48438665678648e2be2c275a640521d8c858dde1277c2eda73a781502f3fa30728f86c125609f570fc993f1e703f601bb0bc9fe489e9d8cab6d991c9fca931d90859a2d747d6104054640f3a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1664f644feaa141bca39b9be4ee19917f2726b2b101ac70d6fe430083d39b21720077ee156fb33c00e49aefd807105b04c252fe5c7d01d05b968df031840b8eaadb99b3e5f8569ebcb30820879b0e4a90c1cc2ed18b22d4a5a6a9542674072ba7f5f4d45ba639722bb44021cab8a703dd7da474db51acff7d3e0bc1c71a8d9f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91aff6c9261cc9170177a9d95e6824321734654af17f95ce0791d75793c624cb789d66ea0d32207194d131dc4ff9c85bbd3491dd187796f73a2f50771c948ff01a2b07f7ff25d48b45b05a65c3c53246b96df4c707d2e9f7b81db10576174e8da0f84b77aac83c527ca6570b90d6f92d0df894f739e53457b6aec75b1494fe12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb15126d4344dc2c95aea5f6f5876b7149d912e17ebe27be37ee3a0c5771c7cae51e7828fd2ef40912b1360d87aff9bb4aa0358d7e5d4d5dac85e912bd4efb29febaa13112c5d94cd473003dfbd1ac6093586bc7118bba84f23d9d67dd633680c819f5240b087625541b12c5af5120c00cdd86e4d286eb5389ece76bee3844dfc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7436bbbcb79212610c2f00c16b1b3002565ce5ba808a0928fdf6833525eea1ba5b6e4d70158939ebb58d58930ec67af42dab0dfd2e437f8edc94b7d5787e8363c0446ca9bc2359e7db2c2a243569970408c247e29ea21a0f3afd6756b67b10b43a698bf2fd48a69cbd48077f863df4abd62dba4e57d3532e52f538e0c4ac5dbf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaa0290daceba64bfe5caa7dc70443e2167365d152d35f71d5c645d29c5d9cefaed34df7f484ca0fb2d719f7966b83a20582c92ca57201e0435b1e4907cf734f203fea0db50f4844e464d6c0127a1a16f20c85061a2950d481cd860484491bd7336d5cbafb32445ce7e76d1ccbdf798e92e2fb27a2065c0edf7d64787087dd5b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bb593329678fcf45024e9b8b820de237c2c8dace3a4f0bad899f80b1b0d96bc035e7e07f26db56889b081fa6225814d723d7e29f9659dee6aea7c9bff7fd73d075e0a6849efabddc829589fb3fd15b647626e4d89f545e180ed77150768c8e364634c60fcc0011dd6bbb532ac6ff06c2c4c891677aa2e729a8107d2a139f8b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae47ba8b2ecd0a49d427f1c8db5f8435fb45c3c120d842740c0b9789db37565d5b0e3af8b88410302933cc33e725eef70c7b0055410865d77079ec3169a4c2764ea1c36753189a831b1f133b26db50999820e2524fdf06d4ea5ab254669abf222af73f1d5123f652c2294508ee5f559ff741092fcfc4a1b007915d903b33b568;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8565a789de8da6596bef8d16532d8a2919ef22521acceda32d40f1e6036db6ab096e00712b5331de4b1e317e92dbe047adb328c0e6308965944ff78781209e66a59f9c1954b26e04d5d02772ac8f4c53844e52c0ec3f6a76428480ef4f51ae489139599a67f8113c1b76359326290b378cc1f315a7588c763b2710e0fd5096d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d502d08c740b9e9909cae83b65e2b9a3c0ea3023b6b61f6437c5144419368793077f2fbe3468c79c3e81ec26eb4d8dd5f269ee89f2f1028fbfce6854aa09233e3b387d53b78a71dc34520af9df3d5cc1d49d82a1b822cf65c31850c689d96cbc9a3538dc5e1dbbc7db84376e61dda2b455ef202b4312b48e07679089679aca3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf21b9b89835048de151cc5e79e96d42c21bc5fa5333a359f01d23952318ea1a19087c74cfe82c0d8c494634dac4b86e7ee118206aef9a3a992df4f4a44402e8842a5c305b2e9ba41714f52900f3671d529a25f9d54c606d0309f90b2eee4786b7a7d1ff865766f99051786ad111566ff54357db0d4de40c88b92dcaa5842a243;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2463ed440f900b37a1212bf217ecf0caec0195c35fdb7c5df108f51971f3605b1ae3451e2814419f33324e12c9ec303f10850efc9b3c1dfc3bf8cb6813353327f4c4bb633abdf6bf1b616c31e487b3828be4128c262d11703c7330ab9ea30701c0ab1050517c9e5914319a286c9c0230aaf8d272d6d18d032acaef7eef8f1653;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde8256b74daac49b80fd3d18209741c94abb9217b99017062c74004b09574eb0370876aee8a997135b2183da1effff00bc5cfc6d2b89426158cf0228ec168cdba4cfa24e54b5a0a2704b913c90b81a5187a526f1e286605c98a3fdc98d2d8bbb71f523becd3c93850927f76b918dc408bbffcfbfc528ccb5bed4c4aa8a54089e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c8b8b80bc15dbf3f78271462cca7dc0531842113f8c26c7565214b3ddaa26854937fb31d5da3bddcadaf11a1685fcfda0bfcf6d108a86ed99d10238450e3ba589bdbc1675454a2002c1dce984c54d36e9a76feff1c935b8f8e997df1d33864a9681c5a26346e22bc7f23045015dc864d081f3a6716b3c448f21fb48206ece28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3fecffa42ca79ff50bae5f700ccc5013416ddc64bf51428440c7cd834b5ac75984e75504f0f0fdb612186949ea6c036e083bffee34394bd1afdd3a1b768612b1402445f69edc697773fd07173511689dd01261a60e9f7ef3b547c859aa9abebbe41ffce0f3c308a9521cd3671c63d20f17abb23b7687798ca5ef05cd3add3b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h537fafedd1aa3b75a25a4bfd6b26b886ec541dc906e5ead47d10044067dbfe155f90a862513e5e1a5c836150183570dc2eab4f9b68a554174b97a41de191c23a021d62b738c571728f7c668e82cbfdd5141209d32b2aec326283436060e8e45320652ad1a12c99e0394ae7e8ad10b2258ecee27c28d71fce9bf0b202b274f6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1aa0256e05cad8f1e00a4546ca4f08f1e299e5e261933767fbdb53fcb0d880f42273dffec467d2d57cf888828cfd6e6b9197ce219232a72aaec28ca96f5fa4f431c6d18a3706e1460c6f5e0ff68b3049cfc3d2d9d1c9d6fadf8e2feea59c123e235a09cde45a1103aeccedc3ffa9c1d6385764d4575cba8d4b4d00e7601662f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14621696d4159e1a0b75366e8e811f8bf84a6ff85934ce7b36dd1048aa104a5bea019a8eb607fde1606068be722f8739b6aab90b6a78ae82b06ff70950556c02b9b6cd47bc729a8b6a01fff0deda16eec9335457f7624e4d8b2f3ccf24fb2f6a4bd6d32d7b530534302be773fd9dcd92cfb78d5c643d510a2c5afb12bc8a8e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6400c2ceb744581d2aa33b8be053099453a1375ecf3e68bd3aad29377721f007ec22868af0392b5e83b2d115a2804c447f535cc97f2cecdbae8ce7213a0621a2243d8dc982cf4f90793bb911312d1f22d99a86963001ef07355012942cae10efc80aae53922e19820c2141470128726ae053751aac5e197df3f96924fed75da0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha28319f270677774dad06932f1e087f181f1e2f0a14c32777821051bb4ed025a50417885b8779b88c6018fd832f4609c02cda60528d880e206be85791cdc0ffa5c593c95b5bf8a70a662630aecfb4f68542165368dbaacae8b50473e1e7d9090d8679b6e51d19dbedc686feabe124b95e2bfd2328ac544d7867451f9f469229c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed57d0ce8cef99dee5329a944ec8ad37ceb12bf7866d71e3c17bab9e0a7effe103fc8bc3750edaa67f5fa56ac0a8c87cfdbfda4adf2230b93b2452142da712d7d4eb22f9bceb7259435d15ed1188edac5885e91eda875d28bf446f34a176bc5bce130ceca9f3d5a018261d92faa05d0945ac05c72498db24eb40a96cafebd152;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d109714c307fb241520028b74656c401943d3c51947448009de134ea7f42e529fe6a1d94f5b60d8bab9bd2f3c702d5e7c3b86137ca5aa7fc089daf7af0ccd942e0999ec90483c26b86d9d612dbf7361965f342682a8f6a211183e599b68a2b12e72333dd56104ff67b389adc3f0463c1fd7c8bd9269ebd59371c1cbb9b81615;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78a55103ed54d32bfacf429e931b8572147edbd91bbee2e91f74d7ec9e206014d5bf58218b9f278104e1bfab31c11b407d131d026ac71f2ea7bf59f0266fbc026e5b2760b69dd0db1d32193fb0dbe9256ba1201d2466db0fcd2bed4f485ea55536de213e5b0fe4e682e2e4088973102ec6d0acff412ffe5effcc7edf8c00a5fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11aa159b78f00948a2b5c0d29ba4f5a377bbac6c2161c504e6a239e9a71fad71937e8b2af3c0d2f0672a9e64b88603cb151485a274b0750d65e0600d0a6f0f4db7f3993abf1900784e440c17d55bd9e91d16bc165608ea73471f86787c224a1c87e831ec0547115566f659f39ccff7ab7378a7205a777a22be78d8eaf1abdc07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h823d5358c0b2ed61ed876be7bd79896336db406dfa7665d79ae90dd569e890738c908e10090f03f13039aa539f82a4e37a01c1c151c5383ad23e5d605df603300938f875e120b721d115a4d6ab8ef68ca5523b1c01221a43e4350128f49f200e919be9fac7cb45507339deb0b9061ccac6b021eb09798e5247cbbd450c871109;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ae1edbd31179331af69d5495b7be8b8553e1799b51452d80a23a6aed66f0437383b66369ea2994e08874b2490d9b00be9e6661e559b035152f12de444ecaee4c005e2e24eeff1002d007f97c0f6821143bf9fc973b7e6ca73e3147bdc2c509b1ea7abb01001055d756364f3fde2d8596469e570e2b69e7496f0685a8a76e93f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf98a204dd469bb2e65ecbedbd52ef38e3e43edb3310df0926f83c457a1ce5998213044bcfa41168397a98b7c6fd0d98c92259b41137f4c6b47d8eee77222a6600342e46be75fc1e6e09cbb6deafaa050db16118145ee44eabad6c20119e22edb59915dbd373409639eddf1be8e2ada531d3d902ece92ac45e67864a0c8281640;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60a02d0a973b706c35af6987bb223ea7406cbba85f649710b957bf7bac88a104e824f6dc982452a71b800ff48d01b54ed31937c2fdc2e37c11bd04afc0f3b37b16b56d8e203c7c99226832f44eabc2a152b74aa1808bc8db829cf0ecd27f2e6ae7eb947f8e9617f5c1ec7398ab17c9c43fd7a797f4baddd207222b85656a0ae1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1603180a5f8f6111a8d45ead82d4bfa0f7b882102595cd97cd1bf8caef838059e32ab5577cd3406c83a7e2cf7d1baff6ff8f21dd46265af8a988925a326d4481b0320d96322985e2722bd7c7dcb336474c7e3c25a99dc6082b5d4ec4a1b98ee3501fb3d03c6d22f092fd56ef0fd8b498b7c09e5e3dee1af5bab429e2861cd00d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10ac167575fe050e251b18e323761a442ea4cc83f6a1f486bc97138e17bdb7b22937ad607371e8df5430ff83835c93b8a4caa75bee8480c20194e544427be8d5a55b6f1a4dc252230acc1ae5253d3a60473f67a8397e9793a85aab186986a2a9da7df571a6070f2b16e43c7235821a417ca2201d60d1ac7987e5fd27dc26441f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f8ea60e8448988fb539db5935c820a793ec66e3c1cb092d602982d1f9aee6b1d8ee179f4d8972ed708fd7d1f1e50037321fe04b98c29616bc5b2a18547d854c3224b770f92f3025e77cabeb9dc8dc174831bda4ecd4e4b130c3234c355416069658c445e439cdf77cf7d6fbc32a7f42d77a011cd9482a9230a386b098f42d2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf43cb3d0d19736075dc296fed2deabc1440a8c703cbd86f0689c20ec930fb1523961e99bb1b913e7bf9ec68c9bcf29c6df9c41084bf54e4b7fb74caa83ab369f4be94b949ff589285274ed8cf5d0262405d0afb5a3460f4d177eafd8ae4577e3560c0b457261513e075d1fe4cf9fa189a4a6a1699491813ef6234fcb397f6d9e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha047df1d2e30bedd5a047ff4882ca896356bbb36628b5999e16c8af007a4ac5501766d54983f77cee295b025cf6ad547ad442ab9e4e7cd005e0f6a941dfb306b0511850c9e9c1f15f98553e94a713c927c9ad1bec4d887840e12c22e6acf92b8370bd4efc58dc3dce84244babdaf7bb8bf1a44a295783b8441ea175c8603d600;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h334eefe5f8a7c650b41196dd33606021d6cda3f079d34cdcfd0b7d108d25b9bb6f978ac2b45d6c6b44ef1fc83d4563dfd3372b6e3b00d778aa92ec713622ecf88ccaee5eabe000b484af19c18d845ae1d741cec77c5f73c473b7e5c7f6a37aba796e6aa23b54569c0eacdce3a6ed76aa2ae1c6ab29ea1b5662ae0c9000d879b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha277ba1de6f66cc6abd88f19a83764a449650e44dd2472d855206f4fbc9056e189f75eadb5970b7d276ce883568171e705758bcbef3b62b48b5e0e7ec29ed8ccdd3383191b7a29faa2c9b359c69a2dfc66bbb1711cc181314489c798739d82e8fe7bca050676f2d26b65345fd7e8eb0992e1c8322beb67fbc51edb619bceaf4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc047a9df6a86061a89ef4b6698b1c3b266f7596d5f96bdfee60adaf26cf4fe70476dff30339fdd09f1a47335a0923a5c9102d6e1e57e7be45ffd9a1f0b6180b70ebac560ee4fc526675fc6ece28e9345637da7d14cad89efa91d0529c4c8fc4c728cd7d87d20d39476da7d2af4b2909fb932178142514fa401b25d594c03967c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc17d0964ce529c72ac82440afb760d2158a4f3c9fb6eda2e2438e730accbb041923270f02a5434822e0e2a37e42c917be07f5b40d010f196f2d8fde0e317b062a9501ec0c40a4d6ad9e6a26c6c569d6f1b84138cb25c1057d6279214d13e631c2b8f0a1cc78f2002a38289e20ad24b48e19adfcc73c1a51b8e61df5b6ad48bf9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7ec4f906932a9591509b1cbcb86681709e8710d12b3f9d2f46d887fd1081d43e61bf8eed9dd5702b6ef4871f2f5fcde7f7745d050145b03e0518c75b753e8af0bedacdbd6b5f13cd6ff8147108e37ed312b920aff3c9aa278734f47625b851bb9e7e2d52d04b57f550808f74e7047ec8a6253cac13213426daf8a991e68b3b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48ba9449e13cdccf8c00d6b55bbf9373cabd3fdca81380cd7857bb8078a28d52594ea26f58ca4f2afd0df9d73ef5d19ad41a72e6e6aa837ad6c5d3d125cb44ed57a05d9d2495896508e741b9ea4a7b6f95b04904a4494aa30311acc8b6927918ceb093a63dfaac5a63556736b97ebb4be4a4cbfb8008b67e7a59b9bfecf7b352;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d58a34f8b759ea4f636f8fa7e1253fb20648636be089fc88bfc468207bf970328473d192e90366bec1e02dc4fec5319894a311dc647cd487bb85e78255e4d67f13d1ce4380b7209ce23d0b85ddee6b0fa98ed9cd3574f98b9e0ac3880c21974ac7ad47b977a4b7099da2482d4c4c75aaf04462d351a90958775437e572e7da1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6824dc1461760833cedbd89782e1ab9dfb01bcb886a5249c33816e7fe7729fe85182a4f5f733abf136c7e2259be59b5906a39691be220f61232ddeee8f23be178b8617260f69c5bb088e998d3a2b700c5a3904b5e18c8d28bf5361bcb5d65728fd773f87b25b6dd945f3f4ac5cab7674336336c3ce28196acafd1209338de694;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf905abf4255e897f6c06c7f7668ef44d031533177cd8d0b45622c75e50dc1b2f25ad4849e82f89e3e3c71fb15a18f60c7ba0a695b167452480159ae2e7c83fa7a74711d795f6ae0918601364d59f724cc226064702a7a3c8fdfc408aeb4f4b4b1c92d393e505ddf8d8a84327a75ab462b06635411c29e4c121eb6928109f9bed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h402d64961923d7f0ad989fc16b3973f4a22ef05ce39192a1e3192429a066e4cfc948b224f35aad52bd6677d6f03bc49f06c8b1b83b44b5598c24f8f7712e23492c85c081d1e1ed3ded48efe408cb66b004a5b051f480169ed74422417686fbcf6c1e4d0c02ae3a917a0f5393b2f21ff0a92f0eb59c8b256f86f553ea75ead10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1be5c6b2ce85ae0b3f3dc544068384f56a8f0e0797e184713a636a34a0b79fc6afa77187b5132443c611dcdfce06b279e495387cd046471d6ce75fb18f3d392caa02c43c8b1be0c5912b733e04078f57f5001e914310df6793a4c88ca50b3b962de2a2f5653a2431b705a2030722c565f89b58b847a6ded35d131fdf27dcf1a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66f70e376926a7e7e8aadfb3a263200a334cfdb888bb430283a55a372131563f23a8c70dc66f9dff8c240229f89d154e411d7446ddcf0be32df34757470060067bffe29835722a1db9fa37eb4c833f06228e17ed51f2d5a590fb8d5475a854ea647d3a935e6bcb4c9855ad0b8b7518aaa4cfd795b3a8d3c35d7f630d6e0bf2b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb17bdc11fceb84f88189cdca5c22c8886e4805d6b76c3278965c5830d4a8c56ff09159e2b2d5c72e682ba0e1db7f549929107c96f52a1d3f0c4bf5d45f0935cebabd80ad747def41a2a3b6249dca0d31fb2578dfb80eb811eb5b34d22cd4be53b3c39e1d28108d82ef0f4d71a603786c8f75ed4ec2b9cc5a701bcec8c13ff7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h953c8722d46356af016bc3f73bc7f34153dcb247a56dd48c7ab295c24888e3df4869ad7d84784688bd582c0a29344c63a4686f37806fa1f0483fe6e5a14cdfa031dc71d6a03ab8d0fe90a41f26ff2bb51f6c849d9f37f8775dbb45e8efebfd857c0dd3ef0e87626ffbe3b7e84eb0add9613b349e6b0ec13bec73fa4e9b1a26d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45903dc6aa4d61d2ac784cf1c4047ccf56a92ba3b8255d6f40e3450cff85d72fc518b2cc07974dc9abe2a3f5d9e2c65e125eefb15f7239c862c384dd6a9deb84ce16b1077260525414cf729807bfb2ea8673630569205d4e25fa250053987d4a194749a0c118d5bdf4e356d5abddae568cb7910965f0c2b850f6876609855eec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e02609c4d1d89b4dfd71221e8457c09ea8a92c7d2b77ed3ecd2f5389b09e1914658915af3d4ecb17fda56e2f6e489b4dd43828bbc8a621b7f4b556e55c381b4608c686a8a9aa97ed19c1b5691f4c66918096f10e4ab0933b9f52f1d819b824379dda3a1fd550c9418fef124ed1012afafca9b0251ad7a7a15c59ffdfe223475;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55e87ed73399669e8a389d3ecb6f14d211e6d32040ab7acbe7462e786d4135ec81ba7ef3639af4bb8b18cba25514d43c21e4966b5afa50f448dcfc2b91262d842668afa32237c77ed9011d8ece6024ff601ec5f5809299399f599326816edad247c9c35c4d6151c4c95784b9ef01ef56099382d466fd5b6f0a720785f7cebba0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba2c3a2f72a3e32bc95f9726909ddb854b131ad379855b97dbe479b25292bc2247dbf75e2f00168bf650a373538e55f4997a0bc786bedc5eb2bb3428b8b7003512d73a89b109d057fcaf8f99d2b1026e51604ff823924588ccc349b35b46fd945be39a9adc5b585284fa184a2ab7e26e56b41d67067e117f75fee35ae319d4f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha78b6a837bce39a4b18bef646f1ff069b0007eee465e6de35019b9dbe7ca6fc3eb77bf4a6649225183107a8e1c5cc8e61524880e582bc048949c314e2374e00a6f2a888ba9c7ee49a1ed6494c5393b3caee831ad36afdda20b6ac8e9e21677ea0e4b6416199f58ce9fbd8ff8647a3d10124e98d968d93453f2b36b3bc1dff523;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f40b693ebca908db9b927cbab7a9c38f2aad4b19bf878f36b8777ac609127a75e2662d0ce6f4376fa67441a0a8a4ea2721cc141716fff08a4a927bd299bddf2c339f780b433680103635d7fd00aeea012ae3fc1810e70ebe60032e6c50a4d950ed61a33ce8afc9728ceb4676060671a8d922a5f4bb1f04a088b73d1b690e160;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf73f7288109426d4edf1a766e8cbcce3675480ffc920d253123734ebf73dc9a8fe92944e0f2aca063e5de9ea00d07e32107ce822416a6e74ba5d10828eeb5f44ecb8a15322e53dab4d7b57c9dcba700d8870bccdb40c1fa0bd72c4bba4f5993ea170606630eb0460e7d17fad7d04feaf556e33f0ce7c7d52ea7bac250c92101;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fc0bb05f1b3c0f067efaac7fc1aff93a8da662819b8c8c7ef3e8e4cc88e69cc363f687ffcf8afc3757660fb418dd6bbf5993f38b8c100f701f0aacc2fa85da64ac1d62adc3b5eeb8afe6c55e2dfe0c507aa6a11a4f724f08d036edbedda989d4127991e76ff7a6d7645e0cf8450b522e96fa0bc7b496ea316c8ccfd1b6bde68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d599f9c8280383a46dea3debe25cb3996acb7e85fb9b93a8abcc5699d45012a783af91db31d928eb31c2bdc6a4b70a4557cea2d7f4aee33a78ca1f3b0a2a5781ee8012cf95e60eb8d5150d99176642d0209d30c457b0960584dd595e0b00a2f7dc2c963585a8768746c8445bb71dd8631f32cb244999d529f4a237f542c7288;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ecce5073706a620884653062e68cc6700b1f603b479caa4ef8e2c24a5141682a12f5cba699dbd4fb0333344442258975acaefea8bb9994d97727da4d11a3c9aba4f6051706d1e0238010dab299639e86004fd10850f7fc5b6a0e68e3f61ee2d5dc2739545e68fa756c06dcd4f6487625ac1234858a52431a5c631c818e092e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf273a78654f352488347f04754b01e87fbedbae64bb40f8ab04bf7c47fe8cfe97725bd025ea09419d74f3403601263337448a875052ec1ca7363547b68e85013fb303d07a934e9ad468afd89fdc49174f5177b61cfbefa308af4423a0ca19125dc409799fd790c15732203da9e9a81c259990824e111fbfa322a6dd6eb79878;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55f9a86df670cf3e0381d62bcb0ae7063b4b471969525129856c5545777efd2310873eebd873af361c0eb17b7e2ac97262316108deabf57d7ed35834e2c63dc67632d119327eee0193edf0a63383415fa81fc530c379c72987466dcc6aebde0452c7ec36731d68b09f7454e9c25f9968dd1ad4b37e3ba325402a84e733bf148b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c618d32f0479f8968db68d247b60084cdaa2c5ec8232ba864352700b8fc52ef8a067a42204102b18dd044b94bcadad1db65c2b6e2b4ce8f8a6bc25dabc7396b3ee451a29fc31ffda31776c8ec298f591a0699e970b7710094cd0303c7cfa2923589cb499a83e57fcbf44351cc8b3b8f6a7de282d2bae21fd3c5ab8f4c494514;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bc1f14371413984a58ec7f5e309bfc66ac888ee549f7102ec1c2146bcbfd396d9633e33ade31ff6243309d8ce84b74fec85af1caf062276c6ff276ffdadab1cf39ccfdee81efc185c73c8a9476a232cfd4c7961d9097758d6ab6b4676be9086788c46ab0fb3a811e6eb5e289c76e83ddac7fd4520661b3af46738847516e825;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbac1b1c39444920b13960ac7593a1e7ad37ee4ba76b5b6e5519cda0e250999d863ff5194193a01c7d3f511e99f95ddc54a6c9266c352eda3ebe6d53edeb5dae8fb16fb8efb87974844376b4aa5ab64ae760be7c86be1dbcef2091975396f505d8a16b7d1c1ce0cf6369acd3f3a86b2822dd79428863e916c5a0a8249a11da3a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60dc8fbce740b8a5f655de3313192ff68229890c3db8a310a18b2b02987f584bb4a8cc4e28553f840277f4085027b304ea3c04210e70dbcb1359160d7daeefdf1fae6c5cc3ff01e2e939cfddd64f096eaed2b49124f82d97448e362c7cbd26911432cc02a3521d8cb774f0f6e6d8ee428bc51c75cfe420a6e2e7e6904ef4548a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28e1296bbea4a92f6572c2ee6429dd9415582fbd4b573e92a450f7486d87e2afddc3bf9253af893f80892a5557ecc1d3fd5d38fd2f7d63cdff82bdde967aa1584d7a87f4fb5ce11ee28b483fed8d58ca4509de5b41d1e2df27c4ce79172a74b1c41dde153c37c0a5622d6d169133be60fe6c691462abb2b1364d423713d6815d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9c48c369118eac381df6c0f5bd14d1b2f1b980c987ef76e3daaa14bc37ea4bcbc803afb51059c33f708a54cd660a25acf1e28ee8f7ce977f6b8f0562ba5cb712c85bcbff7b71b3b95272db39958aab81eac2e49554787ad09b2c79c72ee1d8f88b725e59a89fa990ac5bbd637a70d98f79a7a70742453d1713b2d1c29ed7096;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5af6ad8fbde5dcbc677ec91e2776d9a283bccbf57164ffe879883976d81555a129b8eaf0fe915d92bd413946d5cc47db68cd77621b3bd8a3ab078230672a4b41dbdad6e537b4a2aa42097c2b36be6486d82b61a32c60557cf330ce3ebd6f6b171663f08df20c4c7de6e27d0110fe1811a5e7ef26dc9e9436d296d4e0c024626;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha15bcfd4c33f74adbfb6458fa02af6f41b17aa852d3a55314c9495dc769732ccf6fe10caee278893ae7eafe0b3f14e58cce01de28f4125900c8503bbed955b0bf68e12a56f743397fea58daba6409c387428cb08937e5e5a89eb9bf2c3ef0bd430b000b4c7bd4d87b570138ec210390c86da30df2d8c6b6df1d59ddf0e520a6c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h781558183f412e8e72d3f6ce9fa188b1da7cf8961d41032221c8afb7ed32a35b05998be740ef86cc151a42b628d7e1e9cdb43efc7a865c6b18a4d10a50dc911d7d5e0f0a32a23a4756396d2cef8c53de2d5f93b118c45de897a83651b5b425667e17015af95fd20c53a049c996afec2ce7a1e047821d88b1f20d9956372b5cb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f4840b0013dafa0ccbf7ab73d25b5798b59e1d8a23f7331a2915d44dd4ddac1c1af2bfaa2b9f1df3047b875d13266b85308f9dd2c8b6c687216da12b4fd7d500c12b61bca11cb5d64de346b3dab2bf9077397acfa2c61759f9380ed36e8a66af4b888f1f62c889bf3e3d7b30743ddf90572b268b31e110a28f5c4900c344f6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda29570bd27e4c7d4e9ea8f44ad49de34666873c6c1f9f49f89b2d177232d54f5035e945497a3795d079462fdb94354717ab518c74fe38783aca0feac02b3776a10358dadd809d883b9bd131357723418c35a45f70df09f463f9f27f7484202ab5e01f09a3ba11e304616bfb8420430f521e28552f40fbadac6207726968e37;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h401fa6ead62f6f8d760d8aca15861f2b75756ce866a431291d778f7bd4439c8a38e3a646104744ecb539bc86d50669a91a0f4f04ad7926d5802ca165f1095aa241a386c95f00c3343c513c6ca054a50746518c15b127eb6b5d61ad22fafe3ae37019a233d0743425dda92a46748421e92e896e80c9f2ce6452b9a2c1be8dac65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe41e6bdda8c451383f3773521d8646b85086479827f5fce10dced6d4ee46843afaa43b5daec0f527951959c13828ccfd1dea41d9021fcbb9f31970959781df95242544a991099129e4bb706452648457dae96ad156e5ca0a67e0a998a705c20f1267a5653f738d078719bdf565649fe46bac6281b216a51af395e8cbf45566c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h106867695728f0942ce455b3725f6fda3c7e29a18939b8c1afe44da49b1900c4015dff1c0f33571109065dae4bcc62b91b28357c0d6c293fbc85f89deb6ec905768b6312f735cb7734ae4d88ef48488220e234aacb4190cfd1856c1e52e64ba0e54a6a1f5f517ada90eb98de929ecfcd04e8d6c93604380ef5cf7d2980847c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37168267ac32024058f97f8196a1077ceef7e40d4548fb676c872d5c688eeeb776e0af321c294b1bbeb48afebea9bb79122737eac73a6de5a4e1a7f7a1e91807c846401dac84df3ec5d13cc1798fb7e2259725fbf324c05f28b495aa7d5b8b17fcaa56b017bd9b368508971d3654fb1f18b64fb9abdae41fc5b7af187aeb4876;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3628847043ef5c24481d3098fb7df47e1ee06cb43a9e8ced727933fae58c897d85c73b6a59f845d52693c882c736569615f87ba2a66023faa143ba14c59bfc65fd6802f088799dd64d2b3cd730d99f7c590298c570ae583c8a251958bcdbabfa9fc08b898a4a00bf7b928b83240ca004cb303531dc5e2fdaeed0361bfeb32cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadefd8785fd64474fdf6f07dc8cabd097d8727911fd029387f33f41b672e712c0fa17b03b202938a2d14567683086ca52e2209bc0270e5c931f65071feea39073f870675565594e61d319cb126ddbbcdabc909e6eda3fb7d8877298828a4967a08cd53e0d3a12a90ef0b70d9b09514d8f625c3ec368a1de05e167050d060653f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fd142d2dd28624d93baebc0e249cf46c9cb12c7b1b0028e19ef9d218af98223816b7f3241be1455d2799a72579f3b25fd7ea6d05ad168b0bee834653171c32c592d32a215179cd24c7fcf4f0b9f24d045266405de6ee0b986eb2760747c936f919f82851767796e76cd8e4f2e075d676f729a7cb6e6b9dd2ee83232cb2441b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc03da0bb5a462bd7797e8de16c7e7f79658ece0d76b58a226e6293bf144665527a09d733d489f67462b2b61b2c50b67b3acec1dead2e724382d633421399a73abe3f2f520aab9fb1a63e520a680f011ecfb3a1fb176138c65d95322ebf7a7ca1e7f70f4e0d362208f989f46d35b12f6282aa1c2d1ed3048327eade0abebcc8a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0854db2fef929929788d9c3210d4597953e23e6ca1e154f8a42abced469bea9e3f73de5de0e0a3341d8f273f9a09f627d43aeb50a4f2a9e6ee5b5bafa054729ac46cc0346c4bab4b454b8ea70d079ca4f1c14608b0747e00903ac3876cbb1f050ee20441f9a1037d558705997a7bdba76943d46e81f771c929d66d5dc58d958;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h718283e0ba5731f161636043a5cc0a483cefb7d22e9d5e300c6f9005950968ced87a8dcd4aa89ea552b8ade930c3dbb67c4fb884bf33e404b928ad98f5bb4966d74f3a034ba18004454b46642c97ae8b89d80ebbdda8518ea7bedc6217ef394829270673a95c3438e0314b714ffefdd82f3e4c222b46b548e7e4f2f56a2b2a87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a62cb2813654f3de91f909c8b9533cd01ec66d205658c5ead2887ceb021184edef629dee8c1f654cb7759b8d030b209d0c2b82e4f9ed6aa8f7266634b526ad5303ca3a8dab0f80f0663098b4e62e1712b875e2b57950c2ab76997d69141a36dc5baa7067869454af07c9e1f10a05e039ccff7ae5e0548f641f917f7df30df38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d6e1a55d3bc1b6bdba5f9fd782010ed04144a43ed58072354d186f55fc9e50ff117a069b93f9b5c3413e9bd80b947b5b63910cdfb68a7ea9dd5aa00abfdd1e2c5caae7aac9ae13d59e92fd1d5ee2acca69da50add3fb6d4fefae632970d3185d4f38676d655c29939a3090e5741b3ab9ac2fedc51979e6f07f2e17f864e135;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5105cec7da367f8fc432dfda3d7674426928d30b90f82a815b7c892b5247a5e96c99705cd04290335e065896a8ad8ffe061e611221434b1efc3125ef759114997804f8af4bc826aa94d30040b251bc8c6368ffe2de99e9777876fa873644a3c8d50df89e2f2aef14d99d7327972a5291d6842620dbe81af5959471b21913701a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c74524dea4fa725d117abe223bf170efcec3af6bebd7c5b31d976b235b626ea594bd67e904bb5ef3e7dac66b42ff2291ea81a10c4bc137cfa994380c6b8f5160fd3e4f82bcb26f85733277111401cc89e5cf0f167d9f9ed8d0ad7912091a8b3336cba4ca52ebc47a9577d64a1b0d7743da3c6f9a7787e63d425a154af99a6b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h393512d39b05b626ea577ec9383181f9fb061ff2bda44d2ab9bc734e8f92d0fd9889d55c3ade315c6b623e8557d19493e13b4f56207e30885b2a249d187c6ad23f7d8564e2eddcf28d667b0692ef5a7de28c0032fba2aee3612d93b832ef0bbd8aa90e2422ce8b990cf6a8d2909036912931e35c1203afae6f84b6faec0a816c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb353c5370546b6979f4d5499f9fdf7c1e99a017ebcda777daecc77f9e541b785c5cff26e407ca6f91787ec9f3e75958ebde80d1e1086721c13283d30d7c37544fbc1acb179059fdfdff6f4c76f37e031b2e427cdc04a9d3185930f79e971807da471ee97500efd4d3400092b838220f72610eeaab77473508efbd7a7186f2a06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd413112c9a5f3a96954781e6b484650cdd2b95452f1c2c209eebf2cbfacb60e5a2f5c742889a70a93316565a09d7a0465751d3327eeee384adbcd36fddab7d05e5b036933f33c4704da5320c9e0343b951d963ad004fd2c8db381bc374b6ccdb515c0baeaedda7b0be7e254f46801e7ee116040686ded3904f71559fad13bb4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71de133d781409f5e0ec1577e09bc82965f0c2d631683c35d957cb916519eed1d244075c0edb86d7d95c1e886ee6dc430ead4b8462fdd7bb0a3e775f85cf2b5a39cd536220e70a488c65373162787cd1bb2c452562a1b31a510bf5f9c89bd000a7df18f29474300345909da22884a8e1476a8af15f1e1ac1838f591cc1d809b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c0a755d5255197efbf9caf56b3b6c8424143def1023c7fdf73d7bbcefef91c77bdf018de5d8792bd9da99f69eb64756b3506103d8ee00fb14542610f1bb56786251aa104a643a1a37d7aa97e68cc7d46f6923dd9c0008e2e85e8a050f04fef69cf485ec434115b1bb45e384ccc86f8f253d3e2acbd4f8c40eeff4ad1583116e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3e9fa566b869ff3ea2a24e1d9d5a529a60d95062cdf2e35e89ac84ed90320208b6eaa40b8b0a5ab66c22ca31f1066d8eeb2ff1c873891fb19ba53fe38bc8dd40b9f109ff17e090332c251dcf29df8e282f7ee41fb1b322ee7b43cef4f9b7709da088bf5f224fb5782e62658c724dd72f361b43d44eb83836561bae9935190c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he14f1edee36844406ccaade59cfdf7c794700cc0a9c1f6a122a12f41b7f7b3b07f0c4f51475c0b894e1162757513af687ba0010b4d517710440392e68e901a80c18461dc2fadbd19f4fb30fc5dc0e6826791aab438c5da842e670b98e9b38c443b5acce4afe21fcb7d21e26a064a6716ede6a75b1886f65c86defcecc5c418b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79ba634349a0655c7927719e031d1cb425efcceb0296dcfd3ed899dab4b314958adcbf4de5262e145de117db2f1d697e82e69bfc1b5501bdbff6a7138b2ffb43fc598d4dc23e1fc40183dac7aebe669fbea154b1393ae4a9823c4b4b0187a5bc7a96ebe31cb695435c11eb66df2dddb647d304e2dc59ee2bdaf5f7df56ad4d0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h278622b2213f1a9c83ea92f96df4589e400f74e24462ff2b8a7c4202dca2b92a6ae7457b05d1c06151b351ea13b9ddb668b3811a67c19e734d2427d77d047805a4a3c6f68787a50d5341a738803b842913e9c7d8a75bf25960dc5b573ac604e02151282e9e3d47934d465c12e406e3d1abe973d53f3e5d63d7eafeefae9037cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h984c2da940858c519a1f070900dd30ea5d999ef78faf97a9591b1983472d8dc2554eb195b9990bb0458ff7e509e7d836c7595540dc8bd4772d3c3d53fbb1cf5a5e68635875536e59455cc0140332b995a5397a67f8957e92a7d54cea793ca9b4658cdc763fea329d1455fc5451df0f234952a8dc074422c7e2986c09d1f3a2d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71400bac54f6080bd6d758757819f43202111ad347fb213d66ca626619bd19b2a938f2ef6669508d5baf524c467e786d60d2ad735ac8e63d2d8b6f6704d871715ecfca746232597684d66379be2913044db221f1c2f7f0ffa460af71e271773c606d04275df61027237705645952259ff80889538fe66e4bbbbbcec70d400ec1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb75cf656e8c279ca1b3b4b38421d88b9abca548dc074206f889301f381f5177c2a42762676ed4e3f24891748c4b803585117356c1db2968f7c0f3827c17b6fe737959f74f1bb2416f97bfc36aee4b7498dffd8152da179263cbc48274931f2797f5e193a7cccd2fcc6453f01bd490b5a9c434b9791ff9d587e1d9def7ed30993;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha13cefe3bc34a3135cd026b622b7ffaee9c9eadaa075abed5edfeec74e26563bc96dc65e458906e080e2acd87d03c7f233518a022820b84f83e32fb3da0267ca2492b822eada5312040fda61e73a2d334bc7f22958bbc0a081b258a5373952374af01bd4ae8c61a041ea5576f85f9d944ccec2950f57d9298e7f8f97db1b9f25;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42daeac13b9881c3258adf4a05522acc575eb57540823f9aa846eff6c8449637c8d3c0c3c374ec1c1325c8fe930db76ff834cff7ab31982878b35c678703848263ac475a76a78a8a7b486b2f57064c19fb5e8933b02cbc043ba94e19f02937cb57cedad2e2f35813bb4517a54967ba0970146fdc3686611cfd9881e943e275e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f4d4825905e33b52718bc6b7c0d7a7a0211a1d5550d64a02835c32652669c217ed5550ba249071492acc3addc5de82dbd7bb7c46a426047570f6355867a38f3a203c47cfcd3f25a4ab12097e49c5c5f1a48a42e2066513073b4b5a94cfe2044cbc44e8c268af85a66769ad2045c588d1f0fd64c7567652ac28b5222dafefcea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf15fc404aa35594c98b176d7096f36fe3c0bafe7c3cb37edfac0d003ef7cf52b076d106bb1d6f5aae9be6d4f1c38bae196568f1c2dad132895c128bbb94c756769cef1251cf988d632defa85e9e66bd0dc43de23726f0e21deead1ba8eec036c7c2b234815c12e1ca83725ab1ec68c04b3a74847b76245374801750b253bc74;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h312c663b669af8f2c9708c8aeda681c812d189bc60c810ede68e3947279599ba73a8b65a25cdb01fbe1c443872a6825d0a99714cb94267fca64f6159fcac82c68756d612f5067d9a90e148a425bd17470184640b9a9960e31b4ef3233b849304a1b5913d457d4c225870fd9713b62ba6bf225c869b27c9a94868d472ff6549c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc40ae6099eaba3b708724e761c679b76d86ca1529d593e1e82efc86be3333fd1d424246bb20430e676fb8476c6c15c5508641684a5af77f2b84f72f84372994477dd91130e94c5aa1b345efced5cf5fb325b7f2a79f53be88220e75df9d27b3e4bc3b348dfaf80ef9ebb337694a1342c590c7f9861a1f51bde70fd9a0cc8b5f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5397058663fe0ebcd2539eff9933169514d60f04015dde3582a8111834b14d2966c5d7c148edcd439ecd26f21303e011323f930250825d0488594efacb140a418b68fc646ed68623187a05ef99c84138ba1b4efe927480a9880016fc2f53659830c1ed3c1242caa7b4600a2308fd1e2cb0374f52911bfb04ffdbbd386042611e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb717d4f430be4d38b3df0577adb32a690063faf5764e61dd8e167228391a0df6fc02489a5791804b8a8c98d1836511c242850a957406af40b390200e34c1ec380468cc64dcdaf923506ac4723d707182d90e9a7a4c336daf71dd420754b156cc009f3484b1e15b6212cd9db01bb3d86814aa617434cbc60a060c47c33ec8b2cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7bd9a6832815c26103d415de75d81708e82d04284a531fa2e799a3d40d92d28a34cdc43d73a8e8c0584cba174ca7bced3a31db5746700bdc535d1c169d2cce002b20ffd8a3d09fb4f947b7d2b7853a1d957d048edf32ed445773b07c5bb7cfac54b8773dd51c3e68a135c8fc42c054d72b8b250b0336fceb0e1f6de163484bd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h149a42b0137b40e15531784fe49d590aab5821a6de3dec6cba8474b6e2ea1c1072c07c2cbe3c0a8e0177c6a80f0031e6d70272ed3ee6b9971b2d7edef7d44bccb286bb7ee36615daae0670efa3bacb6e802dc264d023caac96f3f75a56d5a0785d7750c41b79c27db3af6cdaa75d0f844b6820ac89241353e15c68e277d9a570;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3ba753db15cf485f140f81e188935788c4cd9d24233b06a38f19ae54a1e9e4ca6cc4b85cab9ad7b9075f084be382efff3c732afff58fbd8cc7af0cdc24f592069daf41ae22e3d002cf646dd0a63b246cbaabeb496d78301579b6fa7db003139eec28534d1e1b7398b9423c5e596ec0aac407a88b2f5e09b6d8c5621fd7d3fd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h282b7869249ace3dad46df185f58efee924a8b406f5325945758ccf48310623cf647c3125f019c43ef28e7ec949a2f73ae1ff32373e2129f95e59ba5af7fba723b142ff0b3c8e84fbd2ef13ab2822bebec56595a20617d2c1f2bbdc6e81ccc45358fc4f271758b5a559314261f6c36a2a2b693bb19e6ebfbfdb9f2869780ecfc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d80b8380cf558c70bfad9239ac113b2d7979410461fd6816d24448a41c3a14cd0331bae40db5496f8ba4b5d6a5d126d393dae741ee00fdd5ad524ee298ffab6cefc0c416b0de894ce9c29478157a02e60692bdde8f67506ab51978a2e3b7ae549277dfbebe13a854b28ae6b45574e866afa3818750728212aa6d4ede17fb537;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5270da93de91a7e0dc10d303076d82e8b82b12e9ee7370a2b0295d1a47c535febb6bf35d80b43fbff004c998cf538811d6943d4706b21616f8547da8f512dd2e0eb3b1bce29b61b31fdfb189df1fecdf45ae02dd2012d0e757e03a743e3bcff55f16d28813f5086e644e4e6b2d796d01b95000275777eccd6be34bc237ce56ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7969d298a90c9907eec0eb985e00f5497d1f39e9d354e304f3c76d30f9977168238732580f68c26c81cfd166417288fcd59599bd7fbab4493ff01eb77e2aee489178c88158f019d7b02c02cd221091a978c0ca4dea8b7c2c5600a59057407c30aa6942cf1b3067e14d29b457d98453749be54eee70ed6ee06b36350132c3967c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9a3366d5e01d79a4bcd3cfee5c21d23d9afe60a49a3e468b4358a574a01855faa3ba89e1a84dd1a699c60c4cbca30e32ee7587db519ccb30d801c227f386b205706caab004ef126d37cb3a02126e3dbc6a56914c61242175af8e9a94c4efb21d5949bc9f0272633c033f6f426a10eb89b1842dbc1f6dfe2a431e996538b01a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5195b8c5fe992a956c81c55d5a7c570adb3f701cb13ede863e638c3a085090f2380329a08bbbd0fee8a365b15438f4520877a0b199cd6c9f209fc8249517a7c09db2424107ba25ac222b1e260c7d60f403e4e8e5a85bd50f14b6544676ecf7fd1c42d923121ac373db2c38a11670e0e5ae22672673522e32677a0a020a108a9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbac05f6bf0aff81d5d7d5d7077aab8bbc5d32b2553add7e7df85cca3ac206948661b9d2d3ebdefc7eb652246c2a7982b251d6264fff81f0731808e1bc833b421a3536f2cafae40a0427565083229e31053ae0a0da750550465d90dda5496bf64efb1ab594db6a92e7c933c32fc9382b07541a2cd46efa82338cf52a7d4b16af0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35d0effb31aaa81c62b664d70f84f4140826af8ad833a623977cae047234b91f9aa79ce9ae4dee351811ab93996f515acaee3f62c6b9c303c439f437d0919499f1482df09a45a5a2ee63c89b094b3e141de1d9e409579c9c7046f3a4bbfb9bdd267e9821407ab9a0f0112efa00c1501429b0d5ccdfa120798377eff0f2cc8350;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h404075f6ca7a96872f7880f05ea4d49caa81f4a0366ceebd52f708524be1391e1c22de534d11097b86cbc8ed6c131baae69e8ad0a527d9f6de220fcb56fceb0384967e8fa8a7fc370972fb1108675d67253e6efd759b14e5bddd9ae18eaad40070f1862ae919e7f5096ba4d4945a2c49f11090c54036aa63fb2a1ebc135e0382;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90d596a91555e1eb47dc0c78e33acb3040d9d23faa7ed882012610f1cc9d35ca09a1e9ed7f0d35671f53b5afa2928cfca961f8798fd5cfbd80ec33355f91fa479467ac9a5aef890b4a5dbb60c688b0c95a64e3c82dfa6dc54ce8941dfc1c4f8a662d95e82f527a84b1fde5c2e7e076a699e13408f251bc2caa4d874e8ef0ed2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf81a89a3f6c2f271f9c79c9ad2f04622b2565af390baf4e26c857a9d20da62430e5203117985d303168ee6ba22b40c70e6b5f2cd74ef02837c4eaacba92eebfc2ad70b22c91c9fd29810caaaa77ee0f176e696a94c86422796d5958e5625f971ba7086a31ab0225ee03dcd51baf0a08dce19dd82f4c0bd3bf42da64f5eae16f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40a8e828b17440188a4a3d35b29781c9eaf7d864bed7645ccaa7aec7277ae0902f7948372c76a869d688c62b54a56dbc045690f0b42c6aea88dc11db896e9a4a878ad55e42f5b79a261912b7f9ddaf06c6dd6860dc58ff551632d167f7eb16e93d4e0c0b02caaa30b669e9c56362ec764d29b13aeacdbf28cc574912fa6924e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed5a795e5f32117ac3ed60ddfb467a9578022f5e534c62ce7b73df96bd369c64f8e51619964749979e291f743dd2eca7b9d308ae2d444126dcb36ca96fc92b3637127be1399a15632b580db25d5dbd340e9ef49edcc95b7b4f4bb9e74269e9c813dc63a2b129071a807c9cc66fd487fe703ff3d8e6da4e468b6254772bf8675d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he606555b3b6ace5e4492a1187eedf9b8ca4f98f218f66640457438b96211f99685149f2c3b55f3d198fd47e1be3b5203f6fe96bba33feb9b29b5358034a9bbc6ca554e169b3a23137bcbee34c9cd31ecd4ea7031cfbaece2940d2452de3c9e6c6bc38c39ed4c37adc1dd8de9e20027cce79f5fdb1293d141170858821536c28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5479fdb64cad1f11758ad78b21fa1d459d2c05091887e6dd05ca48a22c2c933b511bcdbb3bcfe39118e59dab8c18ac74ba31743c1ef68ba38b46e4b471f12f190d1af4472103b7b29b516d7d0923c2a802c5d01e9796be7378416c7711d55aa9bec2d385247a8ae44a1a690657eb06fbf9d09cb4aeb26fddd035fa09a0b0b95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbeefc366e9f40c77c40410337a56d65de7461e3f34308ac55d527de1122f9a035c723f47d30ab9e5659c11fd240f358984346e23361ebe2bac595576f052b557eb77646c25f87e888a931f526b37f7a830f46e4b7e859fad9abc6ffbcfbeac543acca515b0f9877944d369304cb7fb144facba696df59b648b72167870ecc1f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcd6702714831bbd2036f689f112ad2758e3c9915c147896f12376d5a61824478d4495d67a68d01b2778332898212d39ca94abd60cdb84d2295251c6226a4f8355a32e89fc74365d1db0d0265e75b3ec84a0b11c4daeee53112c9d843dc65c05fa6a9c39a4e25fe958956d668712863ae369f4ac3efd8691889919f459f68843;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2dfe4ac2d22e00670a2a7bf5096786b9dd7465705993cc0e8288e2d6ee4425c2801307adbfc20ef343ff0b02448d01274c39dabb33fa631b06ebfe1ac99ffbb3e8624e41dcd0b5ce71cc9657b8096818d8a3599d1b26f4b6450632eb1cd3594e18a6beb0cf8e246523c0d7d03f50de2e8a4aeade97db949ef0c851d5a079566;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c5d8ed30aeb277fce8521b1bef9229389de8adeb4773669ea06f86d05533648fa1822120714178ab6ef998a286054039902981fd3a1a02473044903a399910a687103a01dfa5fa6119e7ce9006818dde4b236983cac8df1f9b46537a9c001dce1f56013ea620b55054a8b4796694dcf5d62ee3622ff151fbfe8045d2315ab04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75562255f50aea5f79e9f7d76da6e0a5b975020be8d92aeae892f5699a33aca9c4131d09e6321a6446fec0f42250b5ec4a79b4f4dc0c96902f54579536ea24da6bd63d83974d629f4313baf5df4c4a2cc711dd9a649b79cbf0264350fbcb8e2bc8fee651874329da22dd5f9e3387bd2f4d61063bcffdc666910c779dddf281ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h433ffa8ce5c40d4f3295eb62f18d93f0f3654084b9aa5764d4bbfd31e9cec8e0d268642225824eb93c89471207d98e482db4225d6607324ff6cd601a9045857081d9ef4895f426836d2d436afa9a94c229352b658160f50d4f33a955a444143241738d37a2c3be577e9090ef4f2ef8fb498b395d27d0c70ec80b503ab326f7f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddc5d26ec4752a9efadb6162714a0e6692d592ccd822a2e5f3c549cdae52cd39154e0cff83eac14c4a373dfe8160568e4de4b256abb19e1445825e7ff3b2965ac28e159d812fec7f42c0bd731c85e29b11db418f9aad1cc7ecdbdb11bd536acafbbdbdba4c49febf9bb22aac448261c0d46fd2e893f8ebfb0c8a028e8ad1903;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3aa4a9c63dd785240b64470af66dac431ffbc72810b0be6ee5865a11df2b51a6d92251c7719e330937846e394c7961dc2162c9c9a2e194c60808a28160b2817f7b8eccb0f9cbb220af36d1654d7609e88786ea8ddfcc5ed1ce800f35159960c3f1709b1d49d02d2295ffc79e97dd10fed80185fdfc495d428f3902331cf53d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha60bde66d6cc73337a551b1a9a1880780c51b522037f682b638e1fb16b2ea3ec343351526f9af79c9975afbf54a6a247ce9cbd5056b3fb3740f5aeb198be68e7f9e8b189f6f0bf7d1ad7ed45bd954905b63d03ecc908cf76b2e3a1fa37514ced2eef5590cee26c22d88f3d99196fb89c32a0f45690afcf9c938dbd14411766c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf817d5939b0b85468f0f20e05167133735ea6e38171d9a632f180a7d8486220ed7810171b73e5f3a58812d7f0295991a134d8c58d7bdca5b652c602ba15fa88ee531cc57404a6ba56bf6d466f53f66ecbebe373bb0ef9d32c301c25cd3e4e2fcbd80d717981f74b603c50f240f76eb9701d02cf3406fe28330e57fea365ddf6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99ca539574904ef50b759c01b5e7a2612329d6ba0f2bd7f85e6d5f3a41434f203e8852a2630b603cae87b1b6a65f87a04c24f9ae2504c9c739192140d9e5daad3ffbb7df144fe1d89fe3dae89a083b6534c1c0c4a58cc42824a6277aa1b2968d43faf456d94e8791920e5456ed79a64561f9f99b870a8d2e6ee98ff7c7367794;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf873dfd04420c55bf76bd735f42be59f790dc9a99bc05d2f281df92719edeffb7931db9c08672883fcf5ddb6c618e8a207d5a462199ca331e5a75537f9cd726a84064466e2c5ed2c6d1d57c1f47e6d3e0605a819222fb3e955dbb8f2da7ad526f9ccaeb488ac3a5a622b8d83dabca951077834cb99bdc31f19440bf2d8c858f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc53f4cd2c897d40473971d9eaad5af79e62a91eee17ba559beb297b58f4089c806ac3436f82eeb91ab6c3b6fa58c7c169aa9cdb2d5ac65ac96e2b43f73a0a93a0457911e01f9faec1d4d87ffb2492eea43510455edd89e5832e81e1223440d8efd5527d0fefc6bbdbf76e973f3a764b57efee76a9d81fc7fafe1e3960ce2c1d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61f6cf015a773aa93fbfe4d549b5c6f6e8fcb567ab885e0c94eb6f2b3b0938f47574f94e5be8474e484b5fc6cdeccf8911682b4f62068c0216454375af0d314e617f65064f83087cfa06338381075cbc8cc0ae7ed28bf366362bf13329227e89f57134419793ed1ee9b82102ddd1e90c290456fa9ab6c87c37067259e749ab87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e859beab42179148cf54cbd643c0b88fcd8cf0df5429073d7ddeaaf5556cbf714bff00e0762a31fa3186f7be25a30a56835dcfa85e750965d16937523bb1f3e453094e7589edfdf05d8d308c4220978056fe3f4f956bd295b87936859d2add27aceceff7cdf884da1d7ca0a190f7fc43ad2e013db77f8a36bd840ba31cac8ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa6dbc188d1f6159cd5446118730e18e451051c8e41c04ce983a52369c334045369d171d93d5b41364ebc3b0c929682bdfa45c6dda51ebfbad58e1c0adc8e1bead0e64cf85ec7b219b84ae25d55f4c1b389c88ffb466748d01cea167d1bb977b00421a6f466fd9eee9f709b9e553644d24a32732acd7a24bac5339aedaa309bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9101365ef17b930640029c1a3c46335b6b6b3854cc3f736079f63f60f6abf4ffa8ba5c3092beac93dc1faa849b86852dbfac1d8da52bba050af2533641b9a943b1f52924e56536b0652516a963300482961d8c45e2d9bb41fb0a39dc290351e125045a9da739b3c32de8712ee67d4dbaa377bffa8cf82d7ec9710eee89515d84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a52076fe62057ada2eb05ba204658e97277133a63de804efac95c64e3284dced984d46d25ed46fc6441e51bd575616ae495229b0682b0fd9096450e74e94a37a8ef9e39ec481c7539d9a6368dd91043eb4fbde89bf7377eed65d2116eec5e6ce00b12b466e1cf0ab884aae58b678976f05671fd04ee6a00c751a8961f819ac7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed517022ec0c897239f0e4e507203c112e6e206955eb1bba1a868c6d89d3603f37be0b8ca4bd6993feca8a95fdf5659793e754f60571f7a55e6c7b771c827754d6a770ca1281b3f7f16f05910486a5e91af93685fda3226eeca4fe4afd1320fab8bf6de1722d0b434f873129abf4e81508627be567054430fc3e02c3c2c6dcef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15fd26507152f3b959ea9766f412daa0081769ce70df54d3d8942b563655ca578ca3caa9525e16e7ff5c032e5f4dc7cbd47b57a8716475687a9a9bc0719fbb8beafa97974f4ad43b195b0257fa2e98cb390aa4d1dcda3b10fb169c8111d523a3ed468cbb5213e90d24af3ffca545dd6e7f43acd6275e72c8331b8a03e6f1b0b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6f63b7ef22178b58c9c93c673933f13deee520a2d70b734d278f733ba5ba0a92647ba186e3a6f444969e0da545d06508acd7b5e00f19b848e49f36f6ca1c371d81a22cce6d6f6ef494ba2f4ef91b0b04274bd3bf7a4863e7bd8ce6a3839e2b3c3ee5f8948b1c17476e8f98d56e47d68003ecec3f294d4a506fd69a0b12f82c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91e9791cb2500153b16eea359b59fd102c5690115a622fb492582ecee15f21a2b9086652eb9f4eae1eaa89540f666da8ba875f82e149e84dae2d10634a77e6bfd1c8d8bf571addddd83ba04f757c48e770bf37e1f6f6656f91fb915ad3b24492306fdb6423e3a69ae067eb63bbd047cd3b067b67409aee950a8a604c2dce0b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d4033bf0fa4abac3257ff071d41d9b2a1a6be80320a09bdba1aa8b447c87abc571b115c8db74b83e862637004b75fac5a7b416e8c3003db0d1df77eb4c7b14c20509f33a6444e7f3a11575e57f26cf6f5060c1d29ba8a111c56f15f7bc19068a20768e8d24845ac1cb46203cf8100ab6f2262f0c4c7b9d6793b423fc9c24879;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb0dc7b7ea0e9b42e513a67fdfc9581ce93f7373c414124fba2b32fb236ae8b81553dda466899b0031c286d3b7e61b83ab436d49e50430460a29c898a87939641756dcfbeb85396503d914bd7047f407ee00393a4df70304305776f985ca04edce2c4b6e1a9477d5d71538bd6f65ae396f94caf61268e2373cfeef3d2923632a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h167824e6ff14b6f12c59a8660db68e007ff5161ebe482ae53a75fb13304ede40353a3d12946e065b9aa05219bace09a7473630d4df7ff82696905718ff1eea062ebf11294b40523c6cf2824eef344fa4bdc00b2af56d20acc7146b06bd3095badee7304c41e5c66f29b4a975d4dcb34d94df6ca3d1ba73e15448744418e5ecaa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf543fc0cf35ab3320fb70920470a3dd1a6f62337962f55ccef12a90941594bbb6e94cf623db0799ba0982e1563ae24ef5009fa77f889dc69b655eac794db2f558a2511e4f7b9846717a9dca634e9e98e73d9c19f96307335fe1f7aaa9e79bbca119a10cc709cbd0cab844f02e4568317006afe1c1ff6338ff433766c4e60754f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4646177ec2550a56a8c0e3dc32fb59ec1a928088f04f33558b5e6c4ff9244846f7fd89c8052db6233987330ccb201a4f09e3cd4225d8198ff3a75838160c2c154f2dde19e7bd658035d3d7e98abcb0583e16a1aa920b8a77dd86583b117a4a15ba1c76ffd26460396d9ff1e378e69e10de1642ffd97436cecd60f3d0c7630433;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h569a345c648eb7c34c6e4f2ef6aef35c7f54eef31d864f421ff7023826988e36f425c0ca3d86204704a9df576185a7da3042b3d5bb3c189327be8c5f6ed4e1724c56df15345c0840587d568e76d690fb93d7ec9b624945f407cceee7e63ff1a84208a98b2aa4bad61ffef7da4ffa25c0bec3147f2e22381db72019bd090ba907;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc174b5e84f1023e89102df42c301e2748f1cb454e2c98facea9ca2fe3182fe8bf546fe6806510583f7101ed8433a381986a78fd34bc97e26a20c36824d53d4819677d7e6963866e59701a94611284acad4d438139ae522da8170991f8f5b178c1cf46997a118249cf554af9fe1c73459811fda4a480a2b45335e519c13384d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40190c128f36671ecd6bd68d27cbb9826110419fe15f42027c2a390d06c402fb3eaea935e5316e88054712b9e3a5f774e15d819617ae9b245247a5c63d3c86ab4396d31bd0949a05d0f0adbb049faf8da71b183412a20cf764dff8c916d5761608ac3e270d2da68f4ee27391709f6d4bf909e31c3716ba5af2ebd6b5f4f8dad6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6b022c2a54697f8b97527c615bb616ad2c39b44c19eab21292eda61e765b2b785b2292174070c8792fb871bef0cf965d967d536f256296570692dcd20df3dece87334fd2f3bf9a8b2f86df24fa76e90b264abf5665cfb5c1e51fa0316e040ea85b03d43fa324479e9cf65481596903e8f15f7f29f8395618a3c7aab89dea751;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9438a4a86a5d8a88a32454609792de970f1437c7dab1ba514b8cc7e448624f884479ae7f955c0ad4ffdc6bd4b2a38e1d8ca20c0d70a7cd17675cf6420a943cbf4fcb108900e495c954c2724e77fe4aeced0eda8a2a8608272fdf97be8d92b8438c50db38ec6986ab46fcacf2d5eaafbdc3aa54c025f293f936a6282f610bcabd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68aef84d23392811dff6437a2dc4fab478bfd2f096d41bf62b2b8f3ab36d64159499def7ff7b2bb3acd813913ee06b24da0341619d5caf6bc2c9698c035ef703a6baea9ef75d4ada713534afb8ffe545b256634219249420e2e93ed6a66d54a4f1467b4dd9abd5c8ce5db4aa03c800722e582f3278071b3f3ce44650bc9d61b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he72b9920c50e1d2fb050701f21b3b28cb59453e7ac85009377727cac6f3e8b34f4acf6b4b3987005ceb23cf2b34859f0315c084f3f00c9b052c7283c0930023b803b63cbbccd35ad424ca0ead930608f3bfcc7f14d0d01daae6676bb978cfe7f274336cb15c787cf14c8396c028f2afc2fbfb59ff886fa7fa534a04ffa7e6100;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2e2ff6110e9a7f17a27e779d5e09188002577da3301761ec7600a610fbc5b0596131578a81c169885c11a687cfdbe5a0059868578df27983da9b6f8c993b3eefe38b97589fc554006de79335222f155fdc7338191fcd2792a846016268a1e28281ea91e334b9ecf5d496fdca7a986c2f75d4255428aa15ab213c17beaa11854;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h443532466202ef51157adeec61dff500d07463efb25853c4e44e4ca6cb782370487c20d076b090f2e6f9205c04b5c36528f114644f4a4aa643c5c5d558718da3a47a309dd7802f8212ca641df5c2f2d44e9ecc542da825204b72fd65582a62be0cfef5d3ab03b7c0164940466c75b9a0aeb8a20baaa7e9ff5657a7a5fc23044f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69f903ef74819c4f2b8921628f302e7dc2efe00cb73f2c999ef5e073d55b4fde30b805da2c6a66d8898a6ae8af5f3d66c8df1270ccb446a9bdb5365e3fc2ab492f5770a43be1bd86012ac43449b6e064c17dc8451b8b1929adf4441f678db8db79314c0a1e3fb4eaf82ef5bc2f0f35f6d17b6f83fe3a00c3ae88951c718932af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1af70c18156959957357dc8be0e28c1a9b007e515663b5cb99a2383d7fcd8e0f9100ec005700a806576412f067d20d937002b84382214f170baa7a8c27f68e052070dfd03107e0d2c5845ba8b10d7a33925f6bfdf7cf709983b43de953f754aafa9774c87bd228061295142cc24a394c8a3f07f02ce59a92ee008fa2dba2f786;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef40489f36bd151b4cd9c94448cea0e5a1b18a593923ae8d6eae0014f5936311221d20c640eba60222211da883a1ad71063e062681d59121f9926a5dc8e56deb62ab8e85d9d519f9670bd484d465b5c29be9a04912ecfe6a9a38e2ce659f143f571a05ca76418736bd057bf3c391e7300e7dd2a4ab3a42bdbdf77cbdb0dd65ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haee19af2ee163c2eaea33943cb46f1a02923efc313da6856c9b6fab0f71f310f8e2de9bdbcff201eb0cd35f73a53eb9d5f216c8588a618eaf52c77106e8bd109251d57d2c212e01f76043638c959582b77669bd5d08fb1a530017308918d99231562dde621aee22add3e730040bf9544f3221b98810d01bed4fc04274c397198;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16704e7e80b0a0587dfa9cc2853bc79de7ed67cb04feab8674daa741f378231b9f2a67a5226d1d59bd445f65603e4cf4835b3644f7df7b52ec74ef37669025f011388c9ce2e3bc6e22f4f1952990a94cdccdce1543488151cff72151644e23514fc564f50417aafff02155774deeb59e1e6b6541dc67829e8fb5ec0cef697864;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4c6a6dc22fcf9b7bb7b64a2d3e7d0a321360b455bea9d739b447374138893bb12e53c38018ed96b2b0f2e465763ac508a970dcabb28dad23a0e0d2a6987bfd7218a85f4b05eeb2a6152c9d897924a41c8dc6e8a40e28db0d5b997a102034db746a4e738f9941ac4063c8ec85db4379583f60b41ceb8bad3ced96c5d1f3f2ef2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb4258d6c4a62a5e5b1053965bbaacf9ae0983b73689a3dd8d8d850e7f94f658463aeecd32569657ea611b5d15ed06910ac34a5a6f8c35b168e8eb5b6f95e0622ec3ca3891fc77210c5107ee031c9c9f4018ef1ca9584a24da7d450e9a344f16266d4d2c0aa371194657233884ed0a5f5fffe83662096746aa596f0fb8fd2978;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21ddca6f1b93114c917224f259ec8de0f7986872c3b3ba305441526a2d78bc75b791deeee6b29ca8087e271c7ea9cee512370ab5258ded37ac08062b95bb5581bfb54bd94c9a989585efd6b5b872399bfcbfbb00f56ad4e005e370c2add6d959410bc927b076a53894896e58f0c26d1d7420e2658cb4a44ff0bfd6f9f42b1ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ac1d1568d63538db72538034ec33df05b16093a743353a3b6b2473601e963f85317ea8c662f76eb5e02784f447333bbfdc0a6989955d03e72a553f8385b846d48f18afbead8e9e81697f6f6d2e0aef24ebb84de5c94f7d8b8350fec5200cc1d2c21a880d2df570a8cff1b3ba435f1d1e46c53fc028103f89d5620162ef98f60;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95dd62951e07eb0aae3ba2dfda1d70dd9c4bf5f05323a4875fdaf0bdc61c631a86d7632390e68dc21b7f68d68fb35f7d9af704bf487d2febd7370899f20d1415d23444a0d3e20e3e44ff61cf1e4711fb5a4cc67e17c05e9d3b35df1ec9a1010a6034c01a8ad901b5e110fea87b35b4706a0d2188c8cd179028de57544c16d0dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80a8c7a0ecbed21062b3e76c1005bcb11f75c5364227a09c8ed2cb233e4d80b98459ad36eafbd22ae1e450e5428f9ef7c9f9c2b95c55fb509cdc74894cab0fb842c33dc78dfcbf30f80a0d6a1cb95436c546c6d4c0168845f08c13ec4333d424b9932c10a1a8d98c25d4f34792f8bea8ae17e315050f1189219879d8a47d9022;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e198d8818977198102f4c88263af226494f2677a09e4da4b406a25117cdb76c00ef19522d8bf9bbcd22ffd1cccc045ab7dad9ec1273a70079b67569f95d3153abeff1779163f5647ba27391fc32e7cd51bccadcd46b24c02749024d236eafb8a3694eca2836b66a676de6f9c90babee1898b6bb880d8bf83c77602dde19962a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c792b68059b60facb94261ae9d3763b516d62ffac10cb6888bca91d3cf42c52f1575843d18dd56bb0f8043e6c93e9013800a762c63c2a16b19e6d0f8da373860fa0405e60b2b41fd048ad83295608dd0f38fc04ba59cb278c66761b59d9db44f0ed9d0adfbdccb2c55c97732fc5321b4b420634d77a736208c40e2d5fa652d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cbeea1c46eae74f666f7536ffa1441d5eb9ab55eaa7a6d7080b4cb044e4f67bca8307da32d22d43829d33544b698d714cd39ad599d6a510e68cb9f7c90bd74cd3d32756ec01babdbeea910c9ce9cc5732336e485b7f4412fe05322b97ff0dd9210f004d8f7ebba1cc46cda32bc830c7e25042232483466786451416648f34ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a8675844329b9fd0608ac792580d13b386570cb30fc4b4e548b177e7a79b4acd735c12891c08b18560cb59ac5fdd6bec991c5597f7c45ebf76571e5d37c838a1a37e7b27d4837d74d55ce8245d1d6b9cd90df5ea4db52475895b7c7e3a0fcc8ae54037cac5f4db25eca003c18159a5648ebd263e11a85851f2d1296e3cb9e49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98af7028e5226d4e5534865cbe2bf553a3c2f8f89a32efdc69d4e0db815d0e055e4d8ec4bb1abcb744287f3f49344708958c50f2681e34eb07df92f7e7b61e90695434785b5bccba89f939d15778007843d521f3036bafc8648e5a22c862b73dbe34543eb11655866f5e039711c75fc8dffbe95faf90acd74489c3b18eb74eaf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc56ea15e6161805d3e1957f4a6f68c90ad52a45c1cdb4184f7901a45e2743a85c783c7481f1659dcdeffdac3686c59a41033e1a9623274b3ce14762c8f67e415907958f53eb49a23c1975b07cba265f7f751060a3f0936d402a0e878393ff8b2f49fd8d5ccb1372144181bd13f7b7dbcacf612cb95012e8b14855d2c2a381676;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99505cddba035584f6dd9f8758a9a723866c766a5f468da1c305c07c77aad5a6b9545bf5efe95bfdf60a04098fa27bd2c7bfb4866269138ec7046e5a33705238d1422e3d14dbd8a6501136948adc47a10ef5fb7a6be1c51a388a6a9d22df7bad24edf496681ff0509edcec8f17a869d28d2f3a538bd484828a08ebc34d7a73c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf15968bd63ef584a0c15111dd4976f92e9f18e76433994ece04527b34dc06665d23db9361c9b8827aa748416f6c16520fc3d770cdd1bf174fb7091ef25ceaf9a5ca72b5e8d8e36b0a44a9a413968c826cc58ae68293f7d30a5649ceccd955cd10907c98f3445d77a0359306a5a4825d52380f0a8fc0adac08915fb6af668f587;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4efaf85940d24857408ccb6f4221e7a2122c98a08c3fa31599500d501f0a016b4e7211c7b498b6ef94358eaf79b6192c7483122d8bc9a225ae0889edbe4a54b3c11fdc96b074dbf7e2e8740168b3c2eb344207318f6d3de7c2d6572839184be1d3c9fe2dd63f043ada75492f682d26c8a72513ae097b445a2edd55d67399efc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61906bbfbd73957c9353b3a2a8790a18d24262c54d648428d852e6e312ad8d1a97d21c105167c3fdea672ac33c6c55731931397c8c30357405081916363e5dba7a525180faa2d3bc00bdeb26e3297301d544d05bb69e72b48a07615d04e5909a9adb3280b764474238539989bf9ef7420bc8ce4b86496e1fb66ea59e5db12307;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha376ebcc90c1360b60bb2ce1157b4f726de428ca529817c129a88776aa4a1cbb6a97ca221933e7e292b2c5dc093e1b42077dbb1b96f37f42036f8a3e1de512992bda6e22aaabe24bc058bc650b34709d7a71d952b45519e3d0294eba7dc627c2850c4e3cc5be83b317b0a9e3f157f308f17aa57e4552d2d4842077328cb5967b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7aea57e6eeefe6e2458922e6dfd2e930d88400bd205c88e81a5ce06d3fb719d8b51eacce6ea5bc385e7a4faff219bc8f8ec53a4a9cd7935adbf1e76534346abb80295f408ee83627208e8bd1cd638318f3a375c36308af168ec4af2fa15b9701b0a4148de7d83d05dc55f55fbda83df5d41aeeaadad118ed0e833f1af22e9b56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb812bc11525e18420d31b556a035ec90c82f19b21735176e6207ca8a0c783126ee385a7064ab789876c446c1e80b3a4dd8927af18d126ea4491889a8bf88b7d66709e5d990c240b394ff1c6447b070c9226d6bc1ca737e123ac35059623804d089ad97642d1e9ed9fe4031cb52c846e12385e88d26c252d3b51dd37f93e75fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13f2d0b52a9bdb95f730b959045e7bc98cb899cf05398b6fae4aa3c2e4e66c0d3fcf8628068b2a64cce6dbc838b3092f5027b4a0965078ca9125d9c9368199b561a9fc7f5fb11354d4f9622062469d69623c71f8da27b9afd07c374a42b58d5e81236a5c1f988fc9132d1fcacbc11b8bdafafd85c9d55df6c9ab9dd5723b6a39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8db5be2600d57988b4188e63e4d73f697c8f5f404831ceca5c1e619643c96f6d6e81ee9f39fad88de7c82742b966553f3e3d978d9c4f9a44cfacfde2265c04c53f01a49f710f274241a3e342f4ca0657fc3e1e7b8a90dee251c9d39feef8b6aa7766d2ca92f31836e5fa44f80e214073eb8eba83df07b897da18d78156d6c868;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9b40a266023b7c0c6b78fe4b5666816eae5cbbb162fbbaed9004881ecf4e3ba85d69c6673ee776f96b1a18e6701c02ad2361fbcbfb9856944aa66cbb35bc6ccdaa425f474d9638f454813bdfd8c64f1ee9c4d491da01729c71a15eaecf8da67453baf38aa4c1ffdc41498325585e058e7093aeae8b0308e50f0068966a6dee1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2ce9544225124ce648b822cdef6915ec154c82f7daf0fe090d2494e5836dfc6c6d4ed81c7ca7f5e5fe1cb2a7acb40920322bcfe9e5ac4bdf8a66b89d76794738af564d2616e45e73dcf4f4dfcb12ba0ff2fecbfb7cb2a3fb3fb517de75394c65510842a0c9e0e1f353daddd3e40f970f498879d8d227efdfeee22aa912a56d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb297f6dd23c14624ca5d1b9cc3d6e8f65db11fa2b42df85c502007662392f1310eed55de7630205a164b1cc0c82d6c2bc60195365b1f74f7753d98b7b182568c6a941712918dc67b7f0aa585e9b37e63c5d391c413499f3121fcfacb7849833efe743545b18aa4988569a8f31ddf83686c0be534e6e51ea2ec813bc3460c4919;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed7132b2ac65f9cb468899658f6375ffca85c33eaf371bab8dc56fe35e541ca14199004ab502c0dd6931ec58ca5302ee7cd124b1e0a5638aa8eb056af0eb3f0899d8ff00c7c9c67e40bb80971d2269c2760defa3ffb0f9ef9864a1cc1b903bad944012ff7485083bbe13b3e857cccfb78a316edeebf3414abd7694884b6da76b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3f21bfc4d77803bba1de56a89fb798092684e08cc950c9961e944a1ac6c3cf88c901012bf19f33575f39d5b6b5ddcd418f4de2316d0aa9c0b597cbfdaf8a32aba83b6d0ef5e7ec81db60e8cd15b4f45dd1ecceadabdd94dfefc29a640d6b3a95202b5c74f1abd0179d9f04f3b3be3ab23a7b4d8ba1a2f84d798d764154523c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6c362e2bd1035102a8617f61684979f1c4521b9294aa7a022acd050d1c0ab5e9024595a0046315351286db4339c9d2a97fc4c1caae168a31417b605494c177131e431e9940ae2dda1220cef5b3c7822cf3bf890d70bc6fed932368163d5063aadfa0add3135ea838751b41703d11e7afb10d8fdce5be6c9b3257b1baf7a9213;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5e339920fb5015e3a129635e5a4e1be8820942d2bcd6300467f8f3f20cc7bbd3378f8878fae23815d8d264e4f8b7abbe1560e69348f90bbe874af9421ff734150d52409ed787d435982f2a821db95cb1a1960658acd463e23ea229f70e813bd0a3dd1aa527e10e668e6a51597f193b8dffd30f50e1a5acf1f47d575cbcc760d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0b67ad0004eba7870ba78d5bf024b8351ab610e9641e7e65380980762a49ef139a1f4838f33f1202b62062b871d84f7feb99cb54fa72b798316c8daed4bcb59ee6f3b91f1a7e86eedc9dbdbbb12815328e5904a6b2524c3ee0009270cec46d49a4f94452fdabf4e2fd76906e555ddb9ff93ebe000adc33bd05d37ee5412c555;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f1c6204a32b94b29273c944d49092e5691c0569e3e55727a0d37de78cfbd1ce7679da8e7a9a51d5dcb76d25fa0d73843fb90897e9d36b1a3ab10a7b9adf27af61f227b3e0617665efa77236d9a61d9a1f6cbb37408ff80cbcfdf367023fa48abbd2fabfadda5bae3e52a4900b5a4427eaf12cc31900d11115acf71739333fa1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h183164a013cef1a935d569415580905bd51e64814720290e98831b95ed2ec1f0327719447c7e55ec3b3fe8151df26048d8f4afcc42ea1949e74b3a813dea0d5a4e50365d696a3b9f6472669aa8206256615c82aa8e28611a0f649ba62ce4daa1eac71478e5f600980e07cf27c4abe6cc59aeb58af48c164ed68a76d1ea759d01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23e162f9d1a888c347c4e3927872c82ba582fbb57dc7652fb1c3962a53653014d00800babb02bf9913f2ccd7728387831d2f5a333f4d034c0c4648fd3f6b91eed9a65c0a3e511712cfea85a64cf2965f75b5eac8e59886b22a1150fd17fe204697e588c3552f68cc3a534a5f0961d2d82fd2924c1a25ede9f9e6a6a646ecafed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3f4589e4fc646fe41c14c27d75141df03ad7c0be15b69355ba9fd41a3d2c886a11638c12821bed45e2c22ac1319841d7f42fb8489ae3d2ca2451c93e9915fe22c9177a32e949a47bd24de0c700bda554754ef1ece62371d71fff18ef8b5228faeccd2af80f5d10a738103a5201a3a9449bfaededdc511a947cbd82cd717d5a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70ae15b7d3b937b99c156f6164106fc597324e05c7db95e80ff59264079ccaee359eaa339481e666387ec81748d04f7f8be2dce4b93059914b409f4ce1d5e74731f13c4c27fb12f80c66d0eface631e439442d89a76f2ef568a046f5bb82cff3d2d879912e3645638e0b5eae6d782594c73035ea60cebfe136ead9e76a9f498f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0f82e72e22f76e4c8ba1d4b3a6891d554f646b12c521d8a6bb729740576060eccf7ed3018bcfe109feed80a649a9df87caea46a9677e2c4b412fb0ae9a336d58d6a132378b9bb0b35fbd151c9921270e1892d9425534ddda9d5b68c57537fdf8aab3fdc6ca2ed1b5799db6c572a09e705f5903df1a3d4bb05d25b27db0b982e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h263128653658bf30248e176d917c50eafd7d3ee2431621f5f3dc5bc57c6065cd57346003da57a4f2aef1a3ffbf6253528a985872f015b5e96dbaf7da65c842bd49968c4a1294a2f624eb9d1b46437fbbd1561e6109e81cb21c34267cb89828db78c94226c058e98d50e8b77848e171825b4dee72a2846b5af38b6ebf2a2fc560;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5e90581edfae57c292cc64e89b856d159e48ff0001654275fe22c009092f304c28b29daa3b23213c41e0cc68d8986139588af7f54b57058146e661af9b8d20aba4b6285e5ffbee08c1ff430ad5a34cffb8df94e3bd6680856ac2f2f7a9f77f83bed606a16a3836174e066d9c5b9b46034baa415fa04543e4297b856ffb0aa9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5763828a07b720babb09b7a58c4eea7ed3f8d39829a0c93d72e3fb2bd3c04fc98ad7a1a1949eb31a4107731e265548c728e12fa294f608c111b72934ef51eb6859aca908630a9be69ffce6835fe3dc518d07b698d65f7b5d3778d3d1f5706fb067296105a50638c7818eea11d0aa2179154024ec404a60e04b4f51b13052ff4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41b15b6c4d8e95a2e7f40d02e951df3fbd97a60528ddd2021c2bb9708125df845c56888ee78b591c62dba4d68c38743ae4c9f4a0dc587c9aba92c996257b9dc22187faec771ac75f4dbd1f13e24d53f34ab12f9faeb3b4870ace17ded02136b8a99414b2b2305db36f83a98f0d84101f8ee422842275165513250948a90e370f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h409bd56c1a71b9b362841d02108ce4ba18e9f38a3d8db75871aa21b147687c591cd9b4d1a632be6881616ce5e7894127824c4a0231589ea3f4d0ae8dfa8cde69be34972ff5c8a663770e253b5b62b617c38431679f6bbc2a5726e09cb5a2d714623f46414fcc3231d874741f7ba1eb111c64a024c8e942782fc3c3830f61872;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49f360bd3f7a2dbfbf8c2cb240faad45c76180e1c142e5e75a530625e8f339feea22b558147f5ff86390196ad2ef91a01172e4df0cac7c35aac9401800856a8a90c22ba43006017384386772ecbdb61c120ff7856282341c69a7cc2a7c5ba53c381182d10589613ae8ed065e470d5f35fac53b921c53cebc73ec8862916f253c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1456fa8fad899d49a7413a1d29d2cb75d9dea1468132c26ba21e04a5206de4c7ea26b9055aac119e0e1f4cb0131be0d2f48fa071615c8c106511a86a910ac55e6be36803751045692829e526825db70cbbec3aba5a2e57bb947cb4b3949598bbf35082baffbb8e3a6380dad014174b7b1200e62604705fb670cc733b12cd369;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h351737dcafc3359625a4158408f6e1720a637ae5eb6b7bd6b6846bafd946b1aa43237d11fd8e432feff930205cd8347c05e806e941fc560d26f17be1182fc32f09556bfa9a9685c3c9e16c3f208a72aa5233ea941a6697b397de494f4f12882214b7aae3637ac610605de40f5b0be79e05f92e57347dce47960804f2ef5c40a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2792fcb9f4a98af53b171e7f33deab38266cf5c689ee8ad4d4aa3881dbd4b627fbdaf5879ce47c150f1549b5437ac4699a627ab3d4c9f1e93d92a23342cb366fb5b2d030bdd42dd5b85aa29291b21c7a21fa6a051998cb5dbdbf5b87a93716302bfbe4747825915c6e7ccdb6d496a15734b772dc2807e65727c92e3ea10ac35d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8f4b1e052b8de5a515dc17cff090c937e8c9a517be76071c37545130ce4f184313a4fd89eaa2a037da61a0cb8f9ebf523567238cad224c03bf7206571f7b15e64683ca9995f1ff1e3c5aac46ff142a1753c5ccc95985b0c2f9f7a40a1f02b8d5897d5d3ab8398d6312bc257c1da25046adbe87fe38ee7dbb8bc532876d7e921;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe9f181bda463a73ed70852b27a398b642eefa4446158e7b050c8adc65132bdf0e5c3be1c879b60c620dab71e413cd511209ba78d464dd79feee46009094de3daf2c0e473b427e14d94294dfa3f6018d69647b05a1ce2db3eecf5ed32fc69d5f6a10a5bf8922adb181a1860ed34c55133cf91982ef781b1b3abc16ef2245d557;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71fc26fc33d48d6bf6fb2308c07eed1030728de9e0cc5e6fd5592f2edf4c0a55cb7cc9e4afdbde8036017df32dbbb0ca398a55abfce1a7f54cb7a98a34cdd0669c5265e856a4e0ae0dd7cbd453e95562a6e283eb753cc7b927683bcc06eddff3146b37f58183f598e4eaf6b143a2097103996264b36e71ded296488739114cfc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65670a31c9aa7fb1da6d79a26646f8e680fdddc9c71fb156a4625b07172e0daa52b9241578bf71ecbffbb47ca029d898186c70cd68b737be54903d4209d783999b050cb2a063f986eb01221a46ce8ac09e746a4e3464c0e4eb6876030ece6c31a41df52de7e8df9d483aac8ad2e6efd382b28910f158600849d329a97205ca8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70b642f1c8ce066df0afd1c6520973a39ab0e0dd9aff984fd94a71a4fb2adb3ab253575a6f10899700964b96ffb3773387c46762e63b55dc01875156d4eb9ca9bc7d0a8d8503d49fa5446cf6a0a4f20a3c547cc8ac3c34a0a83f89edeab0f21454dba91166c47b65d082e95ff14a9d140f12488ee4816a7b771823054874d0fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h686be4df0b9a9be2b8ec9e675340cdb9b7d89bdc38827ea51c7942cb30d0251439480557126f2310179acc030aebe5291c71f272f70152d07c358a46344792b29fcfcc98f892f262db7e14e1a391ab895eb325eea86c1031270a2a12ae3b2d003b57eebf5c9b953b805685bc0c43c8785f82668ea0a15d97abca227c21733d00;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae8b7e759d665d18eeefbc7c90ee22e7c5153c0be53845efb33473e7e2e932b7d94be63d4e6392695ea983421cc57517c4ad44f3f6fadb2c3f1472459ec8e187946a25d277b424883d76afcee8972b9743c5d963a43c55f6bb110bbeaea9fc01552bf32f08151fba40df3f9e2d6885ff50b308bf246f10f2f5545b1a0b9ff917;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9044cee9562c0fb2a3dad955ea6a0495913f9d03b2835f8c582005b206a39dda488d4929e3f6001a411f310c2faea7228dce766d188766ffb228cd69b0c9f8fc1bf71e42d71a471f28abcc05644f68bc298eb9fb265843c8b2cca07610ec6fee9cc37cfae0308af45ad1b14fb93ee9c0777e24baeb446ec7a952d431d45380f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heffb0eb58e8dcc28b31991a97729dd042d6450bc7f5c789f881887fdec37e4d5f30b036cbd09a0e7af5ca8782a1617fc7456a5e678fdaae07dac894ee5793d57dde193256e78928bf5a4a33669a0b36cbfdf67ba54438f0fe10ee3c0e97b93c47a9d54819348008275ec5784f0a02d4ce3d03d602b0af4c9b5ad1c5627f96ce6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f46b98ceee330929f87db76d5dce39b441866f2176fcd094780e83cca9f069f1491c257f24b1faf78f164576cda8067f4d2d059787fb66fd043f3a7350db825b38c897b7c450fc79ca4854e3e7931ad2796e8ec6d91d799a44b6c3d3c377425e770ae89dd478b5f366430b2be77367351966e150a8f8d740011240d4016534d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98a2b0656db777507726f67f8ff6d28fb25a2510245c39db6fedb1e303ed3ddb4c3b932c31aa3be6995946c77facdf6e2529511839adeb7a6990b9951875f058a11cdf8768b09e22abb1d170dff8b6a3d001c2c98608dd679f002c5ded8930ee2e5b4e0a8162773d6e9f35df82757e4b081c6e978f9cf2971a445b589643d2a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d2943eb99ffa099da23877adaa0ba35c314801e65f2756fef2f5ce6d86c3d9ce1192fb8bd3f91371f25d939c9b4df72cde2ba44a5b4852056a161355782d55e63ea75858f8e208abf69e9cc84ca500c9d9d1e1141df1f5c31dd27cf5e4695464cbc255b1f982e9f8dd3ac208e4fadb0cf22ccc8ac8f97fceb0029a12cdb6d12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdccd994dc3efd8598d516a85318f29bc738ad22606f3aaaa44e1f6c68045a4a30a29a12255651efa1f36e69c9428f94cfcb59ddd229eb0b6d52101c5fc7ae8fd80982938e56d8664bf98269e20f46307e8781841ee8380c3da88998f85f9c9e2d5e340a92173b4ef9edcfd41c386eaea4b5f55042804367ec5d6cce56a9e4ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dd50d4621ec6ce951bdd19bc6386f37581d45817f76c9b48acc0c853077bf000e4ce2bec6b073039ca6bb4c7b96a04e792dc5b9bb593c000615780cf0c9fac11d3c841b52f333faba3ad4d5f8a7e6de8f7332afb9aa9313767eb7bb709debb0d4a445204d6de40e294c3b52c0b4e6f99c500e8b808217fe43f60c5fa032305;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd66ce565e4eafef90cbd3852b01dea51dd196c86cb628e4f883c55c51222649209a0dcc4cc5ce5e8f0996ba4bc28f4058c55f9f0b38630dd0075bd3ad098e532fddd90be1a99dede7577ee5a5538b578aea118b69ce69dbb7118186177859a3ec6ec3b9d4557be17f3b8cebd52e6b5fff815739e50afe590b84d9f12d4be676d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h377543efb3a44eb2f8bbcf6cba2ede11afa2293bf19241e72e7a75360575d4762b35bfae109005bcafe8882efbf64725d29364c9fdda15a0c31dd6bc518077295b849e9c07da23ffde24a4af6690b37c73956e3d28eaf1ea72c38bfa5b78578ab06c813fab5fd82febd8dda7374a4df91338f49301783cfcfb0b6bfb5e1a2daa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8c8ff511d8688bc3e3dfd317289b3183f210289038eabf51baa003858165cec8e8f06a55a7b1e052b0564882f50ad3ceadbd5384c3b982d42d7ef0f744a18539bfb20f5e4819adae5108659f9c3060deb1a018470b467f16efaaf6de877798448b1dca6e1c78a6978c6e3e261e9fabb244b6f1d537fc27693cb9309ce9b4d23;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ca02b638405896924693122a2678e7fc1de34eed00c82015a7686189be4b0938b206f21c42a532f06f229ec0345bea31237dba63c3108e9151d9f19dfe8502a362d3c78d243d2baeb32354e90ad810be6282a89e74bef43785d77a4906930b709038dde315531e02abbf009455f1a6bb4abf2021e20628ec65a72d5ca91908d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56f6cc8f832dabeada97764c2d55b3804c3537c7c846fc995c21e1f6dcdc739cbca5336b4f513e4a8c59bdea26f818c908bcf6ae6bd29ba1790f04a8c9e280c65596a053233efe2c4e8f4fe14089ff28fdf4b697cc5e3278d22931d88c68766c6838a4eb99827b9b0185a72b0c01d1c2d36b461b97594c262cb2bf75c259b223;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dec45fe92ce0ad16541b08fe57a5a214f56f75167a50ab52898dcbb888cd9bec93f68c4be1943400f6bd8d7beccd69e4c5797372edbcb42bf6f1aa1f0fd8b7481cf1f73352c705e6202344ab6eb02e6ce9e1c170670a203d8170c1ae37f37c0790bd2d87bdaa756848b0cd7ae17f821c2cf4959f5963d973a6b5696645c7c44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e284496eb5a1b4819ec723adda750ac4f42c646fed45bedcb566974eb0bee9c2e3e8ac79b8a3f4fcd7b63d4e25af05ee6c3ed019574c6e7410e27aaaaf1904704cd6424bcec299be2ef7fa1ed063d1f7b79b966ae40de8ced409b47e8c89dd634c3ed3e9023d4a3bcd430728cbe0ce3005956e32e002144240f47a6b0ed510;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef6d75a6bd4bc72b271395f7a6e1d736b9b3dc635296d09187c23ce1b65d99eba2bd03d1467d89a64dbae38f67a119889c1f075795e1f8349b47b86e6e7af9a0c131390192102fdd3b96e58e332719f4967cb45b9aca0e60fdbddd18728f9de0cc40a0f740352f5065cb6545095dc233e32646c21aa14324d845a84848c04121;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43723369d3bc988f18b3dcec0ebfd359a4f9eda531c2409d04783f1cc81eeb08baeb66b47a83e67fdc5e92caf18b69cbcedae31c74b7199e39914aff008c5873bf6a63ba9203ee6c0d28bf317ee0544a05436de1745114386c3ff0cce20cf506e567540b7554b2f5d80f5a4c3f01d5a8ddee19514e7722c38826c1a760007d9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42ce887a001589469f472a02d2212e987c4906fe0443b5d64419ebcc4f0834146cc86e3e86298de664455f7b995e04680b41e273f8fcb2caff8c2479aad82ae43d02c50c23bf351a8aa718f4543574f52ebf693a9c061400c3829b86112157d6c5d93ca1f270b3fe903d4ff38adbffcb0fad7185eff3c7df72cd1b58a51e4bcf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h816df04cd038bdf6f1fc5e734ce85f4e44ee713e5e5c30ea2d2dd3bd2bd2d31d7c300636f3d660276b93d6fe3ecc94d524ddf3e1aa437d74230659555e4771433dc3ab79b719f01b0f295966cb9b7433ef8e678526a3e0339b3dcc0f7837b7feef1a0536cd247426a6d0a4d7a73a20105fad782a0642c25bd5fa70340bbef960;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf21a1d189f7dab46d97bf67fdd5125410017fe301b5f9cebfe911b312b86bf4d625663a8862e2fe9f037e4ec72aac813a79d98113f95b96566834cf51de2290f2bc6e81159dd5118aa39248d802e50ec17156b0be10a2c6b3a150ffdfc16273d7a85f571513f2a70cf31ae978988f5e4518ce2759a18f0aec7fba0e96732722;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc705f2da98877cb06122c94a873435a51a578a37dec545cbe035327419b6351c07bca21203094eac41a80991d3e55ecc9e7b0f873431f0f9f4fd6a55473879b92649aef87f4d97f0e58955579c94d4223bfa758b9fe954d02a2ef7ada83cdfc1ee0b70efc6e3a2a47d708431ad175ccd9a6938800dfcdc6204d9ad39d27a49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fa65c5a09f10b5e748333856b8340ea88e8d2347194384dd207eeb9da4db3cd0c1b14afd56a802afae7f5f96b533ce112bf567dc49e4bf39b37cde015edeb66ed93bbb221176a4b7afc0fd7356b1f57f8e58d2b2556b7390e2b32ceef321f5544b9a47438559ef9da6d0a72acc120b17692b02f5184f47a42721eda51e5110f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc1f886bec550c5652a2e63456274c0c336d1b0dcfd310d761d5a227f6d0780117d74c76b0653626af9462da890257eb25435799af78b7adaf9185491e6d1e2886bdb750e5d5288bd4108723c9d1dfcf1eb17bb2e57247944adcd284195475d8b048993dfad4945e5818bf892ba5cb60670f366fbd281211bb0f78e6587c26aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9f3c066e4f3ed30e2f0fc47ae0cf5b4797a088424fe20176fa8f075af25bff79b4cd91ff655da1245fd79e08ffe5679cbb6844651bb5cf8ad52c907ccb89c9a3f98f90a4981513748d4eed8d56783d074ac3e9b0274db3877565b120d2b43b7c81c79cca3d09343a921970cfde7096ce816ccccf05ae515fc1e4d567808f81b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4601b491546fd78137610fde2aaddf90ce31c7d78ec109c682d530f0618b4a698aca38eab72561f06d351e9ec34c6711db596223bcf200160fd12afb30dae1adeec8e153cfbb103ba1fd444d5c32a7694e36709402c360a2fa3981dc4840cd3c3c9e4adb53769fb559f0cffdf17c2afa84be517abfd96ff31dade87618a5ebdb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff8f3b6d20bf86880371f2ff5f6fad5add2dc2bb755f40d0c61c7a49d35ca332a392bcf2bc6721bbdc8ee877517b895645bf352bb9a67532a4eaef1bc6319d0c573a4689a23dfec52384c95e71245cb2fc78cd70f1a31f84f51ca0145b3b5a22af36f06a1d4e374629154ff099fdce688aed6fdfab3200234bc6fdd72f9ebb86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h591a6f304a197bc250871bacf6f9dc3e91f6855405653cb8094497851de562c91ec5e577c7f61ac6aae4093eceb1f35772ddac7d6f22fc7539ca70310a47574aeeab691b239ec0c2523ec8d9f160dded4c64e3adb522c2dd00934df5d06a4b6f54c4df36d9759669c179581b6b4b373fa8bbe9246e8330c269b0c2e072134646;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf290615028585d9a632dffe3712dd7aa9f5214e003401fcdc2d4a2ecc2775bd2b43e0ab29efd39a0cffebfaac5c3bd378bb985f6efb2cf54259b757695eebdc1df53ea5570cd4bc42498b9263087ce5e5d2aa85afaf7c271333d66a61ea3f91523ac0be65d0310f9d226d4fee4e375e2640e9f125d224ebb2e88079eb1802d17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69c4114c5f07eec5961a91afc44f942a66f2739090461c3ef0452addf91d098efb9c075ecc6043793f4d81ec44f8e549d86cebe4c0eb4bd50f70037c92c6c4cc7b9cca1229158c20e20762cf582b07a45cda4d7450bd141003f934dcd1d7f2beca4e1b7af7b668d38dc21d1ed42a18d2a45c7452e8a29ff9700263ed5d9fce8d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1c83149e61d745806d332887dec2f3caa473dcd391e3402c182010c405476301d268a56bd2705904661020a3ad26aade5ef22dfda6e08eae83c94afbbc9324085214765fc079132ae326cf40ebee729f0e214a5abc6b3e3aabad765b6e0299e19bef839b20f44bd5299b14e0bd2d15e883c0b9c208491989388ac0ec29cb124;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ef413b40cf5c58dfcfa9801bef2bca6f3fa703136f43366927682a2166965af32c895a864fc4548364b32f1d7d54aacbe382ea82c164523bc8a5366e90831b847f43b9c554e2317a6d43ac73879191f102bac5a17f447655eb959c787bc1b50eb5286f92136f64999d83df92bdf0d4194d096ed83f32a700ba84c5d23f54cee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce441241fd38dd711697dd6e146e72f74fb4f4220038778dd46f54109b0eff414b03e956c2e9f0adce940b0ec2261e35efccefbd8d95daa0bd9255fc40f5f0694cfdce2646b6bae17f7dddb5d31846d2e858036222a20726d148a3124309a929e8b92dfd682545b53f3957ea79ca14048c84508ad8d48b80485dbfaf21740011;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha50c8cded6640e3d488c6b1bb7d679ee77eb7bde2cbd3e3a8d67dc2b5dcbca875160d2ba228c2a98346f2f8292c9511dca31c8a128e6a9a92e84303e6dcc515e60488d4de00b4b87fd40a3266b80fd9aa917de12654f2fb1dbe6e94a530fad2be35b2ad493b562e4a465d4993de2dfbf0f76a419278dadaba3d690afe368d082;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dadceda7efae9dc70eadc33a61878741bc7f647ad4a58c29468bdd2be8d5d3fdd0e1ff2d6eb536b2496dd0f91a385d25f1c4177c5cb7ce1b9e88c6704c43e6b5cfc5f0eb354936f3871e555e28a1ecae77bc8cc981d8916df43179ed012decf0f1783c99eef9a3b767707bcffc086e8e855642f8ca85b0fdbb5c9eea8b447cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5f8943c8785f3c51aed8b37a3c4d8b6102f7db667f17d49791a3023fac50ae31c24b68e8ea8e37edbeb5a0f765b2334bde04d848c07e61b20bc1d57a022a87f58b20738b5bc385ec422b1a85d60afc8a7c1109afc7e486a3febc21e6aad8548de0f021cbb2ae74aedbbd05167a3854468e1de440f30c1f56337817e7d28fd2a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3aef390986fcdf5741567cd6cc33a5a3e389b7b4e8727a7994c995dffb8f80be7a592fb2034354a43a1e38d56282814a2d649ebab6408dc38fab43a685969145d5e4107f0b0358b8f90e3ddcf6ecdfaeef2f233ee2a77f24d833505eb01904cc3d09697fb6c0b7be1d658a3605e50ae52731dad2df5507a761b4167bdab9ef6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3531694003f339d7c16b67596ddd42eda681b8c54cfabe1ccc5f4bc2276e390c63bb7ca214557f3f556ecba27b4214e70020adae1ba481e89f89783127ba89d00da310d03f273db02a0f6594542fe226cc8f9449597f3ce4600d9761a94b2a6a813bc2d6958f8823da5032a82d791018e6c5b6fb73f5728ca1fb431a04cf5911;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5459c8ad0adf53b025cd84e0487e93ff47f1e2f7e678a99284d5c5ff776e9552eefab5cc35789c68c044733ec1662ab474a967148996d5661744a474df59456b6c78e3005b24d9437aedee99fd9e0ada6a1c465871dc03b6342e88ab6a8b0ec8011dbd22df4bd7c38d77220d5302051fc79576c2af6057cd4ecd16fb7d84ef4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2009e12f00ee81e05f8e6647bf8681d1563518bd2f05e90e3d9a912526b86929a26469f08169825f54ad04a44d13f9ce460760e52a1266441d6feee4d85ff40840de9a2ed203cf04c70cfe13a36283cb6f5bafda34d855554d553d17675a49955efe7b8fb7efbd4daa83c0a519800e308a9986b3b42aecd9f09b873236ad5eb1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb90f8e8329f2da87ad3d57183cfdc48da8c450ddb3c0afd54a3fcf5a705883a0c3da9815a1e0fce0eb5f3fbf331e0086ddda19b106043cb631efc08874316769f7bf6f8ebdeae948f972ac08e19f061bed851a0b119422f9dbd79f226e15d1ba494de67dfeb60b43a8a84b9761a59409c35dda00b26a7e2577f47b9c7af534e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51236a86acd030b2a16ecd9047e47b9b75c58d08381ba72f80cb78981e1c29501bfe1d2654bbeba117c37e80168bbd6d8ac5b4526339e231ef49526dd2db1a3af64c0765cf713afe0a22d7022f503e7510fcd3162a66000f2291d119cba3645a31ca31684fc21407325e1da0e916ff8b9bd149cefd2a9a99cea736bc9a95d284;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8db8b03e326f96b50877aaa14d58c21fca2fb11403d30ebcc7d4d773d085047b93793049607b86b33d8b27f1b24f6541c1e5989343f96f5f9a64709358655112381fc0b776d6991f503dbc7e430fee95fdb064d4400b839165174a3773f53066918ddccf1ec3e300101c6b29568e4d3357944c2c59430b1ad0500406a322d38e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd22da2d666b0345f4871fe4dd058cda62532b7e5ce826ec3f1cd6a1e196ce8b7cd878e79e89dac9e39cdcfeee868baa9a68c12ef020f59dbd8b23b5fbe11a0bd892aeb9e6afb7e1c9c9e05a2946c3a46c585bb7618b1c33da264ed284d57e645b014a8a49f9005bc23f50042fb3d75662a9991633ad75ec5fdab5516d6065887;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6475a99cdd1fad1368e5a0e8506fbd671f95e0d23fcf5fd099ed75b2330f5bbee155a9661c7fe68d832a07c3df3737bb8599a2bf314c29996194996db849576cbe844ce4904d01721d6f08cda5f7bf00731df2baae92137d65ebe38f9132e03e67fbecd97f1e7f8808a85b7035c78212992c87c267167728632570ce4699c3f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f555db10a16cf95e9d14d6cca6aec311e82f1f19aaaf4cf4922d82f48519ef2a4f2251472b82e296401349de01ad772c552bae25e42deb3e989a3325a43559b7749be80e86c07fde649f086fb6e2d2860c3dad8ca257637d015f8bf878f8d1aa68bb88f5a50bbc56ca902c6ce36d71cedd706c69580861e7e5303e802be16e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha94782192546e6446715965794178d6cb781e976eabdcba16427e6717724599dce8ee61e608e01083104946c69ce355f27798df088e78471b11ff0bcb1a0bcff459e99e00c5a0d204501c2bbbda56314666a188b8fd00d78524019f5b3bf9e085c69f8af60c22e4bf5edd31bcaa690eb10c81a3edd30e0310df1c7b43f5d42be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33b5125e54e889f7946fd3399382e453a40d0a9eb04d23c3cb0ab3fa4bdf3664e2817397e986ae49ab76fe9b28a3a693e24632f920c76eb2556d8f83ef2a5e016136f4dbf80a904cfb7407548049269a56b0fdd05d32b9bc6dd368257677d97144bd507203b42a148e05b0b4bb8305b7300d953dbc4347ab0c412242deed87c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb02b25b27438baabf7e1d99cbb21bc6c604d064847d1fc3b6d5ef48f34cb16924b1e6ca49c31d9a7b4d2275da342bb4c974bf94ffb5b37f58740f8d8cdf6616f86363991e891499ebe543356ccbc91932f82b32da3a099333402a47877720cd7ac9822035866d0fab2169d9dd92397c86bc5ce3b6d436ba62db0fefc4d504d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3509add459002b6fe88fee11b9a419a5af90a065dcb1d2f22476e9cb2cb6eb4d57a595497347864a0bb2a73e46f6b894ee22c434c80ca65aa4f528ceac7f9560b4b0c10a451e09a932a1361ed4c5dab4057611ccb18c690d6dbe08316ac61108a450a461983ad08daccbb9fba55362e2fff39a69459b21d4751cd0cc7f27b44b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf670d72750bd2faeeaf03e1838ffa9c6629e5b02565230f812a1de63eb47cada5fe6a5f9e519e843031d8971f78831b182f2c8ba8c2bc192ef53a660805f8b31b31b11b9129ecb024de337b4e49ffbdd7e92470f3db41647dcd80a9c5cc54c998a118bcd6791c0557b61b689c07d1074cd23b4a9fca937d12920fe6c2a223d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf36580e4039bde4b242b45bdebb6d8592ee5619f3453b1835e0d63fc768c9ed7a0b6f798dc57f41fef4e61c9df0b4aae3b839dae3c7b1a05cf873fc143b0b90cf0937b4f250e22c96dee2c5d1be1e948ab02e9235b78754fcd3f9d0edf92e6b234c5b4c68c1f0b6efe8268d57d8ac359fb9ea02edefc024465f75e73f30cc8ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h915e4055b7ebb1b46b246e441c63a17bb53df3c9d59340572ae28df8ef6f5d6a1f2444db6a14535b8543d83e3b27ac9d773e85eb6d33ccbfb4d2595822162d5ecdbe043f1759f8fcd5fdd8f1d17b215acc264b1dbfc559e0e6f74befad31ab365bae0a2b9f214d7e255be24f41f9cac043ee313a3d9acea20c3ae006617f8438;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdae042c87cf1b0d7651e0eeae1dab79a372da99ae319734d502ad7572e1ffba655ac2b39c7f4f4ec3d6228054de163fadfdf1d38a6a3f829239a2a236e69688a248dde21f8987c41da0c60300ca3580d6cc5e9a8c317d6a609c32977d1a53fc05b8510b04205047c0edb5edf65f524a7986c1cba54b812e6a666ed2f9159855;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf238082daa0916e6b02128c9fffb683fc787e2bbd31c0ba4e55a5cf3d7dc8f79085fb0dcfc5d9cad7665c211359a0d34fa7658d3f581d71c140f190e313e54057555cbbbc2dc578c1c8e22984034187833d91a801d737988b7f032320aa36a19f7f0f371ebbc6115075442d58f654732e91b87d9e098cd8f2946855b442aad26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce45d69f4d9d8f2efc1fba6277b6b48f024eea7e25e488f2db7b5cb1e2abb68780c69e997ad484831c2c7fe86010d8b0a0b93fc0e83cbb110f93f7142d0b79fa55229b32cb77410e10b0242997ddee324ecf07136577a139bf76447f98f56ac92af27528647711f45f52747dbe2025a81009bd52e67ccd8360223eee83941cb5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab34520786c33d542224771c03cfb1a779559ff7509e031587b01a026896746ef9a6616f14e47078e4ff5cf1607c0e413d2dda8814f5eb0ec5c2aef18e90a913961ad3e91fb876948d355e467009f43df09d3399cec943d59c728c33593dc8e6888ac4a28f618415bd4b2f1d7a81680257a05ffe4f9ba852ddfc0eb5d65430be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf966baa118f3d3feb1adb29bb9754ee5e686c267433184765bc5bf96edef1444b126db7d6a051095930a8af54b008b656e3fd6ee9a984544c809a9f63523cdc0be8ea12304b734170241c97d01f9ef758635f85d03decdc929bbff4f24f6ddec7e63154afc4f33cc8fa592796791885f9b0b0582973366cd3c58f48e93212833;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha03ebc364a056ec7476b18b7b923564dc61f3de5ce2f2de538591f8017a7cb368362460bc8e08158401e9600f8f8c28357de06b2eb38bb2a9f8b6e4bc4c82766e6e7d4ec2c119e852bcf9d331c38ec4a679aa8558c3acfa4848c6f610cef4dc6d7a122153371257e62fbdbc5940e226ff6c47a2c7d256997bddda8830570701e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf46538fec6f327e49077dc4cfd042f1cca7e26beeeda7085d59ad73e6b8ff28ddfda346564967460a0a408675237c6330a0a8d5084384b397bff3257d3c4dd3ea7e05d68a12c6912d18e211e08616de4cae94e8ebfa07d245ea982ca124dba640a59cda13dec0a98abea691b1a6627b4627038a2eb711aa7262646e452b46d54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9e9bfe09659cea0690354dabd5a8321c997e0bacc5691b40c733b4e7c8f5da307c8e64c36ee27f7af62d9463255016a2b6895ab2d098997710f553e4e6eaaa088f8a5e71b3a19b1435b517bf44363e194dc9db0e1eebb8ffea0310af6a89ce437efbfa74b034da0cd0441c1944d9b3c1987090e3dc5d99c2438ed7d198f92f3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h531374fc116e2e70d55eaaa1b6e26453abce671b4bc1d5d3c00ac3de27a892a756abc947ec49a3b9cdd537dee71ddfd602777964a9268b90426c50c1afa3f26f150b44e3ff7ee9e33ca7a3e406517966a21cc78d93f0bb2e8fae4492949adadce39e0c6ad0fcb0ec95d1ff3ed83948858157f5457a19490c4c50ee29ea0f1c45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39cf11a097cbcb64ee297812d2d282a5981edf486922602d02cb32c975c29fc6e4812acaa818483ec31799342a218ab5ed9b65cb967f703c787cfb46be0c6db53391d420de9557f789e4089cf4fdff961a4832aa50da9d5a2557dce71ad3e95321975143176a3f719988082fcb904ad79f771e8bae7751425da8d51c4ff9ec16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb21a0fab1056841d8d58a5d747542858da0fe6989efa1902d46aacbf546b027ce446a381008010ab74631f6f4c29ec0a5f3e20fcd35a09ca9cdb7b8b79faa5f895c68f8a17837c1b2dfbd108bae37e9011559086f986beedc8117fab59e29905d203d409a59b18e6aa0dec5baf276d429b83fdd0a1cdbb3f469d92884b479ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7985e3ac1027068e5154edf20fac32485f6eec15080dda2f7d682a37edffcd2dc6d8df432362bd81a2a1f11d34782330119ceccec6bac7dec8b6f64f370036bbd5ce40af42c22fd6dc21f06dde7d3aa3224b68e64f0f4b826da95938ac63f19b03e259c4093f429bc95d10f476e8e279308a273b4f6f51508d2e3aff1096d64b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81b90e4ddc2f100e9686fc72b9c9fb5f66d71fc3fe92ebebf877cf50114c94c07f723e0283ec329493e38e9a124e7188a1cd5683c744e9e17f26ea9aa98f546193cd7a347955ba8379b64d06ce15aa178debec2f15aeeb370271485a73a4d0b942cb5de8f5e067981460ea797a50af5d35d7b67b696d02bc7f5f6940fab4987f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88a5aac1f5dc466644a2f0c180134b9a0de062d7e1724cab6ee1ab58964c0fde0996f749a57160ada3cd62b20675ac3d03af259b618a2f19c165e373c43561eb2626c9d4c1ccf9e8e5676cfadb8a61d9ba4c9117b2029acfb2dfbbe4e4f4b998b55c818736c2afc3f1b5ae46afab6f6cafcf1675a4a2802c9dd960ba4b14eeeb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bd2dff5f013b9c270669f70d4ed22e144ed8573f167323caed78afc387db9a07b07e19063db070d9637e13bebed8f733fdac61f92c86658275d1457e58b8b045d28ef5010668f13e71fcf11ab2e885482807447777d83e58c12101445261bfced76d10ac1f68d5addf5851738f7c87101fc7565d3502cb4bd7247c84d5032ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76a939cf2e86ea90681ae6a2788bc99313a5244942f6c090eeba4ecab88f3e6de048edf9824f8c487a451c5020b2a1c0237c089ac4cbc57266298a5f85fa126b67b493db8f44e8946ba125766a08d28bf7eebaf4c6cdf699fe95ca10e187452c248730cfc224d4e42b90603435c7b2e6130307815d913d86a7ba9936d9cd6f05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5830b2c4986313f75f0bf9474dda8dc4715e423e16e7f260b8e9ba8e7e106015fbd88c1b2c9c72ac0f16575b3e7f3d6d47824ac39cfa0dc03c16a22e0b9d57c627858271b4a5e66fba6e7a8151dbd62e8c981f6f7402b6718c1e8d4e977378288aa1d551d71b1e1d5643c5a271ba3f5edc53aa17f6a6ebbe21787b81dfcd78a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2750bbb6077b281f649eb897418b430ddd192e63d2afb018d11e35816444a3b374f1d4f4a79c46a73dafa100dbe526a5088457fc3e6fd36be7e58a77cc56b07a7ec387666529028460ae66eb9167b2c99caa516364f6fb8d59373baca9a1e347c9afe188a506dfaca5e0483677fe4341ced3958403468ed758612d1591d375c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbddfe5ae6e7e2d1243ef4e94833abfacdb9ef5a3e9a12c75be5e4a2dd23d170c25c1848150f915537cc9aeef001efbd5774167de359ffc50f1a6333696d95bb2b71e255ecac92a2256251910357dface1e0e1d04722b2d402e8af30dcf4ea47110b3fcc013c2105b3972f6ceea9126fb87da2c2512b7d02902538a04a55e376;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42e2b8003ea41bbc8a1d90131efbac1000a8ff66c633d73f00bdec0e895e8aae2a49275527e4dda6be0bff1bc2b34c3955e7e4ae895fb390d1d76b458e00b27b699d697dc29bf3bebe33bab5cda92ce431775b0973527338ad7018f0fef9cbea1951420e960bff1e9ff254109b35f5b3fa003734c373c124254f45e5cb499d9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d002d846faf43e4d3bd67dedbfebdda8235b5c3bb648bd7d1eae9f25085ab796d59ee15ec2c37eaf286f0e382f78ac5266327bb23df3fb0f397117eedea84e6cace0d11989e9f29a90e824c0eb7d46d08db0ad81d2a35b64b3d94d8d8776d5e94f974ea0332797218994bcfcc390d21a3a164d0a98be032e93fe37994e8d85e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he75e43d00400efde0c0173c5ce11a3bb1059b40e55f98291a64b012378519e2380a47080044fbab60496a1dcbc5c4bbd6dc0cd0987981ae9baf988bae082272a42020793876c968d81b213621c5928a2b6588a91867ea0d6fe5f3fd7b5cca52a3711ec6bdedea4c20fb5dc00125946d916a4321d178474ff06ad5fa624591e12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h461e20b4548a8b72c9273fd95b1a481e2ff62b1bd464b78aafcd7d36c7b0d6eaa9823a763d4655f0f931b9514f1b4935401a3578ead3889c1a7f059968cdba45d7faf04c49dd24c9664f9887bf150a84f1628eae83dd1397b8d7d94eff63d61f4a4bdd68df38d36b4664e6b215300570f7a4737a81cb6d9fbe0dbc571d0e8a73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he947510aa55024e129ef66cd533d7d8c5daa43a690d3bca04fd489d5701567e447b642ffdae822fbb3d520a42ff4522bd23b2adf4c623fffdf70a76c1104134df3bc038066d93a452f8a208e9be4f3b81ebcf492d32bd7df07e7a398ef37b6577ed5a36a973df58d4feb9f3fb515454a7d76ec269996910059c75101709699d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha32e4de5fd2ca545af8c41b8b47a34bfe3dba5df7c5b7e32fba6234bff9dd4cbc0bec22ffa78fa2990b2edea2620fc8e38cd409d51867ef6152265b5ed17fc2786595b9231bdf82a43c76aabe8be5ad832d11f61acaeae4ed8c958a86d5e51ff6d6cee9329c30da064fd03ad970f10e01b464b5d66b7dd0634ff1ee344fe9692;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1cb64f01ecc67a64eaf16b87403d26aec1d096e21414185f5867c91afafb0037ca1130e160ef68afff248677b95eba09492b7bed1f10eebe5dab50b23e1b74f2d0761504bc5aafd6161141460bed7ea60bac8f583976482e5c6dfb1ec13c34ff720b995e060bf349f794f6d60918c5146678f67c5444a1fb3aaa0f021f0bb4a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6635430b5d985ba2ec02c833914297b33552e94109656bfa82630396fbfc4b7f6a2e04ee3824b3bcfcf04c082378ab59286b7aa0244c58714bea2d2e4e9441ab14b779ff92eabf3220c6ce372f82fadaa009e04197db4356f6557c0f78c9bf5ef3e248952ada3a88cfb158835743ad0693955f996b71909832c2e2f8f3abdcfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17244d260a766e01694867e3dcd7ebb2f54dcac03940b8974c86c9118c73f9e1fbaa2110a2a8be901e17fadb7cd522899c61fe5ee7bbdbb4a469b622b509e086c9da3aaef7b520e54597cd29b6d06b875e2d9654861b1f8266fcac2c39251134abb8c94e664ee48c09dc333b7f1784ca8e813429a358d0a635e126e120a404c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4156a97c0af431eebffe05a362b531d37d99c6aae68d4a72afa4b82d97289236d61d07dbf3ef4e208924f2dce3c23e7af67652d713f02e6244affce7a5deba283278e3e360b5da3e0dead325ae3276604ce999636cf978406087307a96bfae387c0eb787b62e7f4a4a07e88ba975c83fe4261858cca8ee157cd7c94a21f5253d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h687da5d8e3775c8d60894d3820d2af0d9f93c588291c4d94255c114c78b38aa8ed4f743e49ef68accba6b048b22585b0ec54d654bc545d5ffdbff40d3442c98744d74fbf571502db6bc3eea0f8169da7661eaa3cb1e16685193ff74f76f947ed585f8a13365c965e9689ef1f78225aecc3fcbd04c9104bfbe3ce2657a7e87a96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0b533e68a0123e81fe5e1a3c70d0a73c9089dea93691a613241886f3dd404a6005a95013b4a20f60048ea060b5b084f7268dc25574504538d75fd6d4b18cd4038c02dfe8d8d9642c815984034b7208e0c7e9d846d6d9a2bf4d74579f1d06527eb3ff98c15bb3d5d94c626b2aff7339776f63962326de7ba9e333cceb3eb4ee3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h392339e248153894199cf4f866d65fb57ede437c39f1297a5dc72452430b0824a8a613958e29a94eff4ea0f36adcf0b3a9a5589ad7cc99a9a774b3a2addf9ae97eea7d944661fc7149cde9139b82a1a2575f7b78dc223270084e47a0900278d393c964baa9b455ea32b7504efd68826a11952c6ab0a8299465aaff04f8de30ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h232b37aaa0f28f0ea4cd486d6c3351846c18d9380f9ea97a3d7e24eedf2a5a240059aa470aae5da16685ec346b4ac4f16bf251a0e219f08fe8beffd90aab3f2345ec25af8b53ed880b83c212e8ad12453c475c6ed3dde8cf29df7385dd9047338333a376698897a72a1a64598b257143feb89dcec87b9737c498b7acf7b5f897;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35a971cf131d37e8732eac8e896be108c89beae57e0cd52bc5c36da80c71e181d5a7d12bbb85903867deb735087a249e6830edc5238eca75621ebe08182d78ba8f9408e03414bee3d67c34654c437f1b2053a86a51f92d800e9cddbd6c798ba8fd8e16c8d68e0730d30aaa3fb09ad27d4e90581aa2819bfe7e9201c8fd915029;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha58b84ff7a156705c68196c4d02664326d0a48be7acc2ec1dd2d4af671240ff0b278e18e34716f62d0bc7ece0d122c0fe79b239c6c80a6ac9deb47db394de61e419b75323243e449e567c76d0554d96c4e76843d16be8a0bc7a4d57af136964ca381fbabf5ae319c39489308793b413b2ed8c8620c1024b18b06b981f81f43c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7260ead04cd5c979e86a32b763977839a1e73b66fa53543812072f8ea284a80bcd27da87fb5fe5cf2a9f9d9898bbc46f570675710a95674620089cf8c18bc6e6963c1556c1957f516b9d4d3df8f09902f34592aa9c286c95bdca23549a4459c79856c67ce6fcbd994f70cfcf13c55f09cde16e9dcfe513c091f1f85647adc36;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b1c6247a5cb69abc8ad691bc29d10da2366dd624246f342cf877fab3260926ae4c11640c3871f8b19c34fedf78a4b6458a278ac88cfb0c61955ae01d7bafd7a2666211c7c41d9c52937ee996aaf7ce2d77fef3816f274bd5715f5de8a9af5a79d240f750f3676f079b11b8b08a26d694b899d0fde7ee167773742ec4e0d8367;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h238c4e5e22fb99a2c64b6dee675e940fb25c8cb3a4f3af4a992ff356b90a928634b855a6b7c4a3771169dd721cb2792b8a39000bf6535ce107be54f2d2f2ec5251be1332e8d9913e2b9a31f3e662c515e05ec36147ddc00e74e1685403d91fa356e7db0f958ccaeb4f3e644c246061e540c54b0c71478fc8903acff6cb2094ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4f90e19b7c4fab71d2cb47024094494848072a8f4d87d12d9fa8fc1c72b3127d8a6d7eefb06e8c110c793ba4938ec730375e657f7af615c2c58daec14872a5103b2e5e72e5fe6ec3e39842195dff69b82ecbd0e04ce6eb4a9edc1c876479b1c0d4f2b2fa03e540719dd1d1b44ca15d756253e3ec92e5a655a30ff545158c829;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he93488e01cbf09daabcaf3a492f39c1214853d53428428a2c73283755cdf509c884f29a4295aa39322a3976c86a4e413f800a71258f0a6cdaca13a8d4e87c87557fad32e47ea18ab23ca41aaedd5ec8f93f82662d0a219bb7a4e2664b29e77bbd09fa478a56b64331954fdd4f2121554ef96478e022667c7a6bf9fcd8ea59f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39e2f3140b9c0b963fdf2e10cb7ce1112dad40e846fc3e7a652890e69489482951d1a212d4348087a0e7f50593cd1dffa354d423f1c5453fcd2333d9e2ee299e0eb7adb10d0f5e52122366c37efaa9920e5a11d286af24dd144e1a0aab88d11b1c09d7c799609837053f98ede02f892c653b179837245aed0324e30051c60aca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda07366fabdd0578fac96b962109ad24a66bf099866e25c819d1947fdb34ca0cc6573bfd3e26e75d66f2651c1c62e9ba3f5b61f7fc0626f40be2b8bd670cd1c65bac1071de35b7d4be1d5822ca742fa440a6e8709f22901039be5bd26e64a9587fe03c294e32ee6d218461a745dab7ed127a5db3ce0d0784d04da9ab8bdca5d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h485968b8efe68641967fc4470125486c5a4e1b7ed2e318976fd514d2096ff845c4ffeb0f629586d5914d21af1f73a23ab08ece10676fdab1acd9f6b3ae3930b0fe1c7ee22ddc37beb21864c5f1fa65ec852f7e8cafc153490a38780151cef4193f9c901e16ce01b89f2a9eccfb08be33a93eb36694f97f1ad7576c408a33c2eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f95910024c2c61e2bc6b4d8587591320c23c76b7fffc71711de30d958ed1a9ed4a91883164bc7e121e554917fd813417da65e463c477d04aafead28a5e6008ec132d0468296eb7793215e35a8aab6e3f0e08103c98d420643a6b5b3f598d1ca0489dcd6551c9aab6be28830016ae0b2486679a9406efd67acc9c86f4009afb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf92aa3de4e086baa55ea0404ac8987267e0b21d977e6e99135899a2139027b63336b1e8ed5d323171193b643979a72ace2efaab6f25dcf75994ebdd4476a78e6f4e1be6716d7c30661f1c24c5f491c61cefea6ab04c5820414eecc212a8741a90063859cbd508391fb3b0278cea4ce4e7a410922edb2ebd868d1e6a498d6ef41;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5322a63258414f69506f72ca26e25876e4ad2f87c34e16e95f7441641850c322370b5f0f3c6647669adce45e4b28263ee7f714f65a8cc52ca2f7e345512a82ea8b441e000063060bf2f64ada8a6915206807d6b5bedd085065c17733af4c963eca0ce584afb717fa8de1f41f8af4ef1105b2c5b8dcb823800ba668ce051c23b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c8d348c6d02adfab2755005702b60ce3b66e32efc53c68fcc87e8217ec1aa73d4c68930be0fd9b974db9c003acf31068bc7677637d7ddd132c8f1fe46a9cbc81c6423856ecbbaccc26e4b7b3179d0fd7ad1db5492b39aa65b88fbd6e2a977d817be98749ef1dabb4f6eb85910da977c50ac303e8f32cdda9c68cecc94194900;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfccde786ce63e9d2edf3b63c466ef8e0f0a641b32f39c5ffc12c4fcc24713489ea17aab630b481ccfef3aba4308caa5d747d466eb7e0e997fc4d80d9b663a5cd70ef6ab919efd0b076828da53b829f86ed0f2f1d377603c5b463f0ea9ee17f7e6f89b2ecbb02e73f5cb087b01fe3a5f9c5d40f4b76b1033cd3c3920b70a23ebd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52186d7b0e2048547643103379ea801bf6815f4d3d7997a7f7abdbebb2ccac8876fb74ca406d8cb9de57a9a1240bb270707ce3914e2136e3c3e4a031c00e36a3f38f347bb06b9152b85af873cccc056c55f35fd2534944b9ce09c3fc7ac50d582dce01581b1f1383a3d54c5e67c19a793fec04bd780d69b2d0bc4364b68bdb9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha51bb37536aeda4f322761cf753d643c78c7b8d45d4417a455b3483e04f5ab7c0c1a6fc2f7c11f691ee253beae4f1819bea643b6a7401e337798fcf95272064227e0c9d8287474527238ec45bc967695f20618bbb31bf13cbb90294f71dd133dde72e0e223da81acde35c0e8fcea2a3ea1b2dbe18de7f91937776bf409f10073;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbc8153b8cedc14e19546d786882896f1d34a6637f5d7e61b5b6e5d3de56879cd41d434316abf3436e13b9a84bb0d3072ca153d3176342c07ae89e34529b597af2098267fb78f61c4d9b3bd167b395af84e45486ec2a713db2485c7ee13e5cd98c3cbf22aa9b7d12f5c3a17be471cc16d61222c2ae56ec9dbb8e93091c3ed6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c7e4b0990b070eb643f1aa548433a774829396c4bcd73f31b6919fa903c52119f03c558b9edd29923519c3753668559e4ba5e296914efad0dc4e1e4dbbe596c115e6c4b9ed367044c18ae7f3a5b2af662b1463d3c3b5d4d94a7cd20081f7b91ae42364fa5cf377f1270a66e2df0d60b31e8b73ba2ea7df24da376f49de39ccb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc3a4b0c36418acf5baf37e3bd2e29682cd72988de0b9ab8be60fa3d1d36a62ceb6f268cf6fe0bd310c80171c5378f54cc408deb71aef4ec25981a18b58214edb277d9d75246b121ea6ac4738ee77f256892a2802ab41d63487e0bfd5c09d12616fa2c2fcd21938c92809ebbd4cc7750f9793b52ca36366bdbcb120fc34e0dcd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35ffb96f18c369d8b9e231bea04757870487fe2261b3badee962ab621f99f6fa7e9d5275ae6ca30847ab43bbd47fdecf2c098ccb5a697477093735cb04697ae20907cf826c59325e4c7028de348de4a4868450642dee177890cce09aa5c13f49883cfb3a5be4c7da374d6ea4d5a4995aa99c7a4b19567c14acf51ff0fa92f8bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf94cdc7eca13b1bd595c9443d6c663f16436b695b90f1ed0360cb656c4c68d7da004cd89cc80297fc3fdbba95e6cc2aca8caea7977526dd30ee8478abd0f1a073dc64675096f1e7cc6458967701dbe2209cb4aec003a00921f5c7782aa758346adff9f469191def977a82c3c2596ff944a4b00c015818f6a194b3c96202678dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4807f52e863b5bb609e06920379644b5f609c5edb5fb3752567adb1ecdc9319f942da0ab4aaa834e5307f6133571eba3287b0ceefd6e13ce1065ca4e0958084be3f71b73343bce6b3cf0b7ab28ee289e23bd4ec3f2a3992ea48f209db77558ff0a9ceec84416f6c19fca0010404138eccd1948275d6340557bae22419a30072;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fe9d2a6a33273d817e0121b26842704e1cbe3df105434640994ebcfa7a4ddc87843e743d4795f752e956ded4fb54123ead3b768763a39667871b5e48327b830c392d46b42984b3914ef4ba6dfbe30679f706b47ffb04f87b076c837cd12f7f4a2fd27ef7ecd72554860fc7d2355ba6346250002be65840686dc1e981b624fe4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c86f1410fb681c11968bba3d639e5cbafdb1651b42886510459ba143bf6d32fd546bbb64670cd6e149c740854f5757033a047f98551d77f904498a226a986f8dcf4cfcd40fd69f655322d18d4b21348c0a5aae0c7110847bbec435bc4f0f8d2cc9a0349ab996777b4dfa777f873915289c70d0044797105327c465a83a7447;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2644692a3f14fc55787b54addf77980446863b1cb432865eac2cd0805788c33041cb0dafccb3f4a8a9bce3cbb4f7bc71520686395a73c4b864d50a090a72da483901a2673a9297404726c339d836c09edd7caadc4ecd22e7cd156460f2b81d5a97d5c0c4340dae08890dd7500b712c9d93e28f43ec9795b981e9b1e11e0e8551;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2c82c093a849c7bb577fa37d20514172505d1d7f693eada39ccd069a539a850becb6d572dcd6b5cf2ec10635dd69168f87efa03fc341cb37848601b7e87b8ac3b485c5fe8b7eceb59cb7493965697da7c8b022422db592b7e52817641d39f02d9954ad62fc7ff5363957bf28909616e67ea500c22524feb4f729af18fa25adb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc41cacaf31bfb4b30538ed71fbaff14877f2cdc6ea30e37588379d4204f1b1bf1b094678b2b0f36b390fbe070ffc6b210000e5ca1e8c177d1c71d6f01fafc4b3537e6777465ff49e0557114fbdc2f77803bb5992934ce4f8eb6d6953d16b98d61b61dfe8f303343d5a6201fb064cdffe874a31f64cceceee754828e2f9433a02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h134426ccb1a044922cd50c64e7b065bc2517377246e33d1a2599c5a616d8937e43562e9ff1a4cde628816b71385dd3b5e280d4b052a3a2925948f1249df37acae5273a8677ddea0f772f42069ec2211c4a10d18bdb5f9dd7945e7185735e2d95294923c099fa8b15aee93ce4cafadbad856887ee9dd6a1d20ba65a9baf322812;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8efc9f201711382442b6a1d0c984a01b13e991dcd6303c234ccaf3b737ffe6d297ce04c56e4aae5d0e4298003f05ca4259bdea4daf58a1f2409ecae2e3b9b7b24e6beee313b3a74781f95327bdf1b546b21a20b30433d60fea68d4dee42d8555b2f9877d7735aa1ee53073aec38fe066e74e2e8594221001f2add55f04b0ea5b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68ea5a1c113ecfa3406ec9c6b0c1dc94e9c6aa1b19578138056d84af2010825444113dba8cd81023520e441841be3d0da115e67ea86214388cc469cc6b47da0766b4f744ab556239cd8c7774fea5e3f219a4f6bb5c1c990f57468844fcf1ef60f8a0c19d64a638c208cc0016391dd6ea4fccaa7aeea0a97b5febf3e74c7cf966;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hada33dc00904f92d46147bc530f7086dab9d41bf26443e5c1f473cbd9cb98ace838e01d366476a39d814633eebfcd7eb9ac3d5ee0d08db8aa60946d98a86fa8858b0141132f56147ab4bd00c8d78e15f67601c253b8ceb38488f04f48fe0412c59cb74f64f55dcd20e1f3082659385881debc3e0f93c8c8cba6ea20e962ff361;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab8c6d721d47e3d3cda47d0f2ab6401d0c879092eb31eff5f5d2bc5d944eb218636182791ddd0fad0a11d211e6b5287c24066a6b654db0606fd3d981ab71bad007e18b4f069948a1fff9a43d3d71579fcd3743058a716822acefd6f8fd3a8f6f57def4758f585d6a3802f54eefc491a24439eb34ac609c49736590bcd00529c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdf841dde3102422181a9a2a52d497a8157fbc5cb705b00bc9a3ad9bd839e4ac68dcf8abec244d229e92e6d7f96cbb64b0cc5d9dfda6d43a89f0c5db568811cf09408a04adbc3a5498d157dacc89bac2465128cba008f7b88de003a668f79af5c6ed0767097385356d79ddb328c79a3756a94c9fd8668348f0c98ad9ca6ee8c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6c6220248f3a94f27322f5d2c64450337c7a647ed0780e54c21cf2f3c44cd0b11369ccff2db25adc996a796e9d2c45a3d09cdf0764ad630b4acefc75cc620b8d1ab481f814bfb114d9d5374b56d339fc379f4910c5f191fe1655e6bc662d4b2f0038675c2a234fa3ffae4d659cf40e0c16bea859dd2662d007f2dbe48f2abe0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h490ec6a9d8509a5d382b88bda21a5e566d7a466c0f4ea4cd0e9263d0267c061cc1bb55b0f6feffc2ac4121c17ca10e5b3b6f5afb8244d111dfd483b2a4617ac37ad2802086d5c422efd8342a1ad7547ae8669ba6c6b32eea20bf85ae52f9eafcc5285579cf95cc4b9407a6258a0e4549b5f7cdda04396737b814d4e814c65628;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb15cfcc61bc5312253e8a218a8dbd3c39e4171cbd93dcc1fc864335a1f7197bc9bc45bede228775244c2ff0cf5bfdf0b904eb50a3e49bec69f0cff071ded5d63cedae17d1c485012641e1a405c6a87b0a83940d875558cd8e38415884ccd3db396a3303e2568075c560b5447bc45a413b76abeac4ccab51938aa43ae9c974f94;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75b25a7369e6f5d66622637223c84e658506b729cbb86cc28634cb1f0e4888d7d55e4d0636c7b3af9a6159bd490e80b7e3ce9d8405542e0a6e4f0cc45c787744503c4e1d24444e83610728d710300fc93f3945de61e6111f9ae64fc791b40735b80ae3b0d8daefa046caea48dbb57fbf99894a7ab19949f0edd27dc805b35893;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ac7e7632a1d84e893e0bb1de016b4f7a6ebcd65077b3ef0be966eaf388a18b6461df507cb21a30055a2c24b5d0dfc4769a568d030a37af79c19d89ba144992d04a7377198f440f42b4229661e6c4b91c0a032c413aad416cca51b8154baafd206cfbe6b26580d9bfa4f1d33ba3d9d6751e624efe7f0ccc644ad5b884e415d92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8d3f9ccf82a2129a34e347f18f324de9d2839372eac515dcb95363d0a697f86451a771b3c5af55b19283b71ff826aac2515034d3b99dc6b305e846687e22ce9ff48a50aad93a7ef14e33542b06940cb9efb9ae99407e1005a342f7878e083068408406dabacdbb94f8b9ea032f7770301f22d3fb600215da1426d72a9d3543;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h606665679e690e68f1bff415e2d17ad65728c5b1e26aa914b61e65914d557eb133c1a2fea743d7c1ae387ee046a51cb17283a18140a8ff4aa3a4d8b7426e25ec805e88132ef9ebeacc13264e4156ec850cd5cb4cd2acea54f9ea8b4b52b1c5660af9ec5cdc5d8d40b297a3d1e1f4ea17c8fbb0013b2e1a2fd2feddb45104b049;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd24a82ead0145ef5a567551fc1e5239fc36e1dade3fdc10b9378165ea579e7929c6d03c3d947016a63666a8e587717504b9245ade803c00996049c62941819390f7fe695819b2f747193b289f1a87f2133081b68545f75d76e26ffb16ec1a991818c21f2edcab19134a05bae2dc3ec7c223bbddc86a66230dcee85bf6db83ff9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdfad5061c5eb448c3dcd2bed1933f2e4cb62801ec7d72ada741f84fc2991add0ec970e342ca4782315bc7effee7eb9e3fab99f34a38672e13a73bb665fbb577f461071ceeac724e7cbdbf40172b0c895ffe647f019497e63162921567832338b2f702892eda4d38ac945defdae75a30abc5b03418b610af77617096eb69b6a6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2e73a9c9baf2045445c575e551ac34f4e359dd7797e42f155f66162b5e3a8d2176c641dfb50526f73cf752d425d2d46b6a70c39722ee8e710bf3e0697731270cd7e28d3c6e42a76635d3b30194aab614210ee47e8fb99b4fdfc81e85ba6e64234a3a7e0f86ab370ea08bc0b1e00186516e8aa230744c2cb6a22c046e53e3e07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69868817523cee8212a481ddae0bffbe0cdf400e8a4f8bacec70baa4f46997ea0edaa77728427fc3be2b8e74ab9e05e5ae3c23501ff003209b8d97449181187585389b9b9dae0a2854227735681b1f03744b8bfafe0fc8afdbf433b8bac64727ce85c0ca23a0c3a427baf9577548458373cc08c56f2d5bc62d208c20f4a7d4a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd7af246cd66e7c977873edfc03572e60e2ae5259357fb6b66cddfa8ecd25a7f425c53ed8674896b80ba2d55117bfaf42afa51d51d2362ea5fbe46fbab86f1f12e6094d5f602611b3c089833a9d13fa0d5915d31e969dac3c6651fb7692e2b24a3318c38cf3c02130c332ea9a96e99cb85433914811d84828b97a447c8fdda6d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8844bf4b96545cc130a63f8f6113df5ed56cb47810873c9835ab4ade2e142e4e4016cd6b3426a2f8dca212fe336b68db45d2ad93b9dc98436d63711d85d8bd94f4b533c6b9446d1b5c4dd351028cc6eb49a1f52463aa446cf4b4764812ee2863320d8601a6cbd70b1550d2fc7578a8594b68b24b1d5f563f473c4372771b2743;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59d07077cf8611144ee3c94cb269192bd1c7626435bbf20086a7118113a5c13c69f176e07003bcbbe75f6c91bb1b5d77be9fd062e3f94628feefbed0adb765ec6f2874b1058dbc8bfb11b6378dadbd88d47bfdbda479bb123a8f42463814d80545d317f0fa44482086a597bf425b71df161c605b62585467e14d34c115b77c27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4af55c2442bcfc4f3ab44fb6453da3992fe96ea7b369c8b1ff3175e794f1daadc1f7c962b011af542389e6628fcd70a04bb11d0c9c4a77dde0eedaa0092036ca3362007834ada593e35dff6de994c2af11c1fa542fa1d83782e1b75643d03e3609c063bdf91fe95d8c66db458908ba405abebe2cda9ab4a8a03db747fd758fa8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39591f4e1e5494eb0fe81de03499b3d0fab6dc2a6e157324fb6d43bc8ee21b8adf5adff798a202b231f4ec676a98ac995f2b5f95854ab0f015db4ca1de41d9fc920f7738e29d7382bd7e193861dd79eb7ae384bfef6ff0c6af5ca2d1ae55a5eb93017802a6800ce71e3a11ff53ee1fef3596f987cc0603a4d4d6ff096a3378a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d3e8016b593d2d4d6dd7bbee554dd74183aabe1ffb78912a06ae83c372692eb376a4881d3cf7334b7e5a9907c21f08bce2de65e93247287ad6ca261079c39cf6862224330e8c37d439c9be85722821f9c5f0781d796923f2d5ad287e234b76413c2e91964523b2d045327527216e8cc0f144e9d480b43e80062f1c2515fc3f8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e86b4426fd981fd2f8005401ce38f03bcb4e87b8e492768b657be5382d68e70f4e84ce5f33143e487e3c045c40e60f0d84b95da48550a6b5a856147c5bc7fa6d0da89f5c65c9be44501cf208999ce84c3ef0502ff7be4f0ed7e253920772b9d75bd66b880c0572be69480b4c40438e990eba9f4a795c1ef332d05a220d9245a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadb42f5d5471133cd5c7d2326f3e4e5dcb6b421d6ae42f19a842ce02c3a629dc1f08e45e58f9ec97a50fb977370d69209bd856b7fc8f3f07552ace51d01d5a4e91f2e747224a24edc365824e5d17c47d8a99a27d6e56ff6a4ce33703594688eadc7414abaad3f60de741f3f1a0988c298676cfe259ce3f65f3cfbf754405558c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ae18c725947dbcfb115070b962c6ef4b2641cf902e3466d3ce23eecce9331f74138c8869556100055f3266287c59e9803f56410f5ac013e71f1cb1eb19486f6e99cd38ee9950d726a91e47cab25d3ed0d42126e347736f9425ebb21860bf15281390ef5ab2838dabe0c90ecbdd8233aec866132d208ba272d14d097d4073d10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6932d4610b352fd681a09972c91634d60ce3dfd42a90ef3caadcc40f8cb66188389120424c07a3d93eb57cc626d1f50a4bf54d8ee6664d94d7ffd7949b67846c2f678a9436e98031a5391aad4b7b158368b261e0eb318434b388f027109f78c1c1a27850922e77342d46e2a3a888f5b038222b4d42389a252ec82c648ccfdcfe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3afa1cdc07577c76a9a17d3d1aeb842be6c242a8c60c68dc7ae2c2fdd5121626a57db279b82f08410698813fff73b6dcc3703b1d2e7710cf574c8c6c70eaa98423b92c723f373b49948e4e0e7b485f269411e1cca45c4c5ef51f8ce005d03e51b2289d920de625cd9cf729e45744248bb7eb06c8017492bc090ca31ccb8b93d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9baad34f4d228bdd44bb7d0797f235b72ecbd4355309d318d1d8baaff6c2ef0bb1a188ea9f78862aace05891fc619dd8014cba7ab9d1fe996eb512bdd85ede94d8b6e4770717c6caa1f2071e8550d18e7fbd434085821336045c2b10b635a5e5356fedeb22915899f2dd4f18705a6539ce133adaf5b52fb8b582002492423839;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf97b7f336ddfbe79b498acd6994108e3df94b4b88ca4cbd26bfbabb647facec703f1bd0422c1dbb7bf025c6289b8a0c5308bf8130e98cd77355870412c6a189dcadcd3986709b8e7ad40f3c551d5dad356d1fa8d58ec6661b4dc47982492f2ce46812d6d06d150fc292d7370588107df050196bb8f99021589807455acb83414;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f115596b6214a21d16a388011a2f90ed7a13ca72aaa824d55016b5367aaa58f386c75123257e13e6a7d41c4f489ff15505dcc80a4a93357989802d4da5e22034592f8a4709f2f008b9e63b10df9be3024f96fd70dc3cb3cd15bc90cfa5df5e3c7488e0ab430785c3fabc2e13ea9302cf72be0d0c3a413a9c8413398bed64db4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfb62fd27d04b580e8dfaa3b0d035ef425b08a46f8787eafa2055358b398eb240b21d5f03bdf51152740408f162baad497fd13d51dd5a960284cd2f18eddb679e3d3774f11aabfcc8e493bb97904634d4199944e8fa7502ccb17f896875cb03775a83de4df6da9502ef9e9f5c4cd427e4ac05aac4814a640285a551ced4993c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9bd28431ca35978ef24f3d79b353d6b4d615193e19cb8359b0266f90824d6258a91b7c5e78a50f44f8213f7d9a55d5affcfab1a1eec1b0c3c14a22825e7fb722d5cd85aa9e910692d0b8c6287f9784e98b2ccf2b704c6cc645f5510cca81d81448d3e4ba9f61d5e2178026bc20dfc7cfd0bc4f7bd12652350046906436d4075;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h632b7f2602487c7878df50767f4a2c911debc669a6af284e9276f33152120cab56ba537fabac7cae8904329bcb5c071ff0ac64b242503e6b6ec91a1cac388a47400d6410903ec5afe116e6866434f7ea883c5f4ce971b7e59ba6f594acb2ab565f3d505a192848039056c5a47ab9f0f24f427e0a0fbbb0c377d815eaa4d4476c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15588409d47966329db8eb936e5950de4a8f8d20159287f339218fb00a5b4aebcd8b67f4a8a53f49e1c54b49994c27a839ae4df803d534ff698f0d53321c6322b309c276d4ee1a2199394b526a626c62b0acd8146daca16d58757ef8a001d9e5eed05e1161d9c459c85838423c7434d174be4ac756e5ffdfb4876861df324645;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h271fcd65d7b717e52e923291584a9272320b15271f57e7a5f2a3e414d36e9447f492e94b1b4c64f808efa19d27511a8c972f67e96279bd6802dc9f4e7a7038988ba09fd3a5baa5e247fbb140d9f8b329632080969125e70b1a34183252ad48da9803f7746e367940c8f026b01e6c88d1dc8bbc4fc5ac42719552e67edb86a3f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a144a3096a80edebb67cb3cfd4786b2e24a9679e457e5226b8ea76d97308cb0cb9faf045d60cd2090327052a32156237c856108783c2c6989135656b83c21f3e8d74f093985709d477228a0c78345a8c47211dbbe448edeb9d12cc804c6880e84fac74d831aca04408886d4cc1f43262eaecf6fa9d34cd63a3adeb36026c98d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9e978f400263577174eed1451f6066c4b63434355bcad16af282d4ced07ca8497c0151065259ff20f5f7deda6504aec7259656c27b269051ab467f53ff1a5186c37c494654af20747290b1ac489630d94c3052efebc4b5e7f7e08bdc33d6e32826cdcb7c8b7d3626b75948b4dbe422a135c806cd5538bdc4a6e3f8da3a56eed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3004b32279000e79970b26870cd9b278e1a7c131f6d92a271de37f26de8a56a3557cddffdc5ad92695311f36cdea8404f69bbd9ad7e3ccae306c9ea1ba1ee076a2663742f0d1a8fe5e0a8529799e4ee37a41f8ab4130fee1dec8fded24b3bdbad528fa9728a90fbb004e1d47ab293ebe27322274f03f40ecb2709ab892f01ca7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h682b045b0c96a58a0be69f50bd20b40c722b01dea12e4c0df055ec91998439988d6bdb58a2cc753708618749aeaa5da329eba9a06c45f179811907f832c5567c69595b6596bc263889a03393b63b96c0c6af95c74490f133c444f8a559c688bcdaf1e07705903bc299290462e42e600fd3f7bfe67cd15014a128ec9b89417825;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d012c423b223e3136c5cd75469caa813c0a8130cc8f95e47bbadebf4c484e4d0c4aeebb8d66b58ea07f4427a2f80476ed8f5757ace2e150d1f353d52861116db76ea15b3bfcfe88c4f4e98786a4619287064b463906caf277f413945e5089935d46dafadc71760d0d34829421a85c5b05d216a996a8ba57a9b0973084d133b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee98b6b677e8bdec02edaf0c7b4713421dc8d26ea280f84025b30b2dbaf26525a1c973fed65e615ad8401057e35ef6d9043c1461bb914a89b0dd744db1974b1c86fcb61de277ba85adb4a4cf92ae041d6b946b3990847fc7bf60638fb51cd628fda161d2f016686cf382947113d735703bd7162361168c2fedbf2bdc2e3885ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d93c9acc287e98053dd09ed6136c517234278616bf535827684574eeec1e628ad804467f14ea8cb9c36f8831d1bd9b8e95ec3c596f6e4b4ef983c9ee8e5ae1a1ac060ad2b2b9904f1865810a94dfe99b857b2f203728a4b963be13cb9dda0ec9d59c48bb44dcb13bede2984ff984a66bb4cafd53acf68097a142fb9fcc75fd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73eded0ec654202841cb4835bff0af371905654efb7490b94e77fef936224f772877d39e2c741f1c1cb0c13f67f8447704bfdf3f3da55bf72fc011038fa41eaa8732133a6c192b322a87db89bd220eea332ee252ddaade6b1c03921a625f00ed5364d0ee3ddc44369698e9212155e3072e8b72b8187560ca2b499f2ff8a1d8dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd68a4e5a80995db82e17c46414e0bee60bb1cc63764d65e7fd6405882f69aafe3b66a3a0bda62b33bc2f68582ee700694a00acab2bb0f0f00fc7c6186e952557ffaae8ac00b6efd117d58f268aaa79221225de7a61c9280184f0a251fe912ea8ec94b4adb2ca26dc38c89b6e293c484483721da2e1e0b79ac2e28525ae2859d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f0a819d722e9244642ccf2a7c30ef8c9070552e24825fa298b71bc9469fbc24f3d766bed09cfa3f710d06ad6730f291e3a7c11aceaae836d6c1403e6b53ffa83362c7fc29c476db90865a7e6dd81f0e2a2046bbc58cd4f4d62d5dcbb6b05990d81d9858a7c8e6cb22eb1bd874696217dd69847b97f93a913d4d117f809c47de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfbc1c583f3d274a929288e43967324c232ae43187acbec849bafc6d446409b38d1607326b54cb8f82d05abd97be644a1c55487ce9f63deff8b8d3f95b3061c9b3be3026a00138d6c4b7cbd2ddc5cc848ea928b17cc07e27cc4de41f456d6a66e8cc9393a0b1384ca057f90a2d9ffb9ff4e736b0771215dd371787899f98d52d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde9d1e1101175b18fefc1829939b833ed235186bacd91743d1a48aa6eeb4f5eeb92c7b1d1f8f415d9713cc852563e63a9f9f1b9254fe133fcbbfec375bfdc15575e02d2231dd68eee1196c1e3d3e407256b52f1d7d0216cc7f55a764749f51d63e0426be5c2f55d7e2a7b0a4fde04f7789e0ee3cc68bab74cad37f16aeda791d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha74a6b43250f627b2a881e91654697e57ef10f4871ad42eaba8af8c297322d91900f8691e3cb63f1b9c744de720b68fa5435e9fa8de06a7492350bb61fff76f177cfe301ab6131fd6f820776b87209523d16d7827b731199b036aa0e1abb5cae161eafeef1deebc1f99fe97de7092cb9bce8bfc9de9df9c68e7a79da5c7e5bc5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfa1d9e38dd60d3a93eeda28ffe3ed4247604a5424a48532f51f3168be9fed11ed1245c7b63a5593085c09a18b52bdf1ccece2fe3efd3004f3578f544458db555e42245b5e606f4bbac042d1f1e15b5b49837e4e622ce02480001d4a513badbebfce2d61e554340d806d493a1ab1d7540d37827406218c4ce2784f652cc25a01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6a3dac97a48d722fd56b5ede9497256e2c8090ebbf7cdbd75beb3ac1e9ab54a3f78b52585e2a8e644be9b446632acc881541a3afdc60d41aad9dcb229a3283ff160adde133959a11c9eb1b29f49089d661cfb9334870ca57e1af61ac312c17be44293dd09a9a43787aefabf975c23237824c13b61d5f2f93aa4f445cf57961;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf499aae22018d7d408d58c85617f6f141a365b3cd4e6326f6d863e4c5e405977cc03a1e93f50815fed4a66733ec61e87574638b06c09cf52d70073862c18584788b37c957b31c70b4d8401f8f3b47908cd2e977a98d2265931096be25e42b419e82c9aab40e97a678dfe5a221dd9699b1c4d63fa9695dbb4093833d69e599c6e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h180106282f4d8b1d431540015d574079629487c633fee93243b1fd620588c3c79fcee58f35fae523e1c7c9bb83e672f01d194e3f04b9d5b917541740dd04b6be26604f73b82c5e0f36b81958e90a19e4ad22952b562aab79469a8cffe1547d6ab14cdd00acfe23f62d452fbb66bd18bbb881b8c8bd574f4e44067957f487969d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea2e0c34bfb2bc1b56feaaecb5c30506b0b41c92702cd3772daff1d02a0248175df84cf2d35476fdddd77ad62787497fb4125341c0ab5c9afc224a25613bd0f402267c7d83005f90d270c58430aa5cfaed8a07e682215bfe3f90d15b976c160c3c10c6fd5b498d4aae030675182a1db75b8342d2697b80063e2c40ce62ee96f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35ad0498e0bc2d1322a49a830dd4be4e87d0762b7d4bfe307df2d0372cc2c96435b74845381acfe637e6646a67bd2ff465f08023eefc4fb8e41228336a463cc9b862f9923eb984ee1f834d6d913156ab3e25f1f7b11b213cc9ecc039a6d718ad9c46c0d1eb825bc500ed7cc7280c058c98b0db9d5b47c72358d03124487b0f32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5d2d53b7b9321ee69169cbbfeb4448bb800ac80c80f50c5533163da30fcfad7aa78f32c0292cfcec01497fd23db4986aa8682faf2df3360b361df916fe2bfde2681f5f44d54688ea018ec9d0b3e114dc3392ce365885eeab58bd11febdecb3c2e1b45f40edf502c41fbf87db3aaecec8668385af1356162dc05b3a8950e8dec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h201fa6c8fb48632f8e173ce84109fcd80464b89bedc005ce4ed4464c663b5b496f711ba4402f690a1f33650b3e426f7cd6bdcfc19278d5d6f8d786360e66ad36395ed179ed1115d9da460a293790fde221233f5c2b381a125711e5fb0e08f2735d0db8530661134bbf6fab5b3979f5024bf918ccb803c83689bb67c23d5e7b95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3b296c76c8502da103bd2e247b86c7b86600e12163cc92bb637c0dad6818b5b530c0fcc1d230743ec6de3da12e9ebc02d94381f8708f7e6d8d22cdee95e88bccb76766dc4c7edfb5fd5a875bc330b82d4df550fb7127eb640ed0f99dd86ffb283bc561ce552de02a9564d4432d55d86300867b9877320eb9758c44cef61ba6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b6af368bff03146c0d76642494eeef2514a5d0f9543fd69fd1a4df749cc5be0940cb5cc8f8ab3468165769fb4a4ebf92adc479127ae6ae677d7aee1ecfc93798741d6a4db4b5f82a13cd0b5d0b0aed1ee59ba346e579663881f440213ea51cf79ae2966788234f0f4ef140845d3d281c016b543ab97564441587405be3fc66d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd50ad8f7606b230a2c15973c2244f34fecaeee94edd16e379291fd5fa1393201ab16c995e40d228181eb18187fc50fb24eaffd37c39a17731707c7d3a2e7acf5e22c951c64ea937ea0bb0de7fd5f4d195a11c7231a96345c8c186c7bb0f4dcd94f247bceba3ab159b8668857ca99993ce27e5d26b116a3a0434731ea75854e72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h701cc73560587ec4ee4b66769ae5951a6e873c80fe8ede1b7aa5f3de539fc07d79a4d9b04c41282d7d346c6b8dc784fd07745086246a0a6c7ad7c27544818dd122feea408fa65614f9dd0a478439a51bdc77e3c4ac9bb06a73f53414831b28d17a2a771540b06ed939e8c03728ce7d55b4836e6f26fc7527e892b28b7ee2845b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b3da9b228ceadc5275c4b229ab0c6d90ae40459f416cde01e32526524fb78453c0610e5ce1c1f3463f99af6f55c743311ef6da7266cbd1a4432b2ce77b6811e6159c278826268e1b32dc428baec581502d9a3a3c28dfc0fb3af77620e0072d5597d9abb1e8c23bb0f48d0919fa51a3f8a4ca4bdeb14a4eff9365b990d87cbd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0f57afb317c58f070f4e4efb376a7f6b5b5313356e7adab66564aa7ada12a5b292bd43e5e30fa2fdb7258c468c7bf63465c84c03c8a34f9746653dc5f010ab670a76eb80068bc9cc4bfc11abd11111868ddee931f14e30ebbf842ad43438ea86f2713b653daf23c7dee3e99f808516f383be23e60ef10b48fc77422c22b638c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h458cb4eea0451aa02a2c40c7e904d3d2de360ff5b2fdf943eb5680025038e4278703287f1c1a65a7e4ac330088a537b0f5f029b256020996eeaf77e4b4e5c84e3ca1f593191619467b4e8522a208aaf9b3b47e9f65a01a7c0986b5b48c20885e69b872631130f19abe701e4dfdef3e752d50a0522683f448addde405e638d812;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb4c494a9b9e0ce3572e2b3e4866e7c04f2df30e30387080f927e3e5614f0499ecac45f2891b0a7d3a1d1550037abbf2875d2813ae1ffdbce4ee7150fcd845f13ab70c1739a5323ff9444c51bfd779dcc9d594a72a0bc02fd15e60d171bece9268e3fc69d642081d1701f6556584e040748776c6cfe520b513a8f49357632d0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb58e930d4a744c74019c95487161ce9880942c7250ef79222d2997dd8db060ebcbf3e4c05ddeaa0ff638f2966e4c0102dd1b79ff4cd85d0ea333dfc6115e8c6eb42334f456c476b2b3b96158af62ff4b662fdb1f58d95f092fb91497f1582c517e3370f960451090dc1a717819c74e7e1932be21951b9bdf3d237984b7fd3fb9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc1d9486ede0f065e0a09e071dff01fb919dd9e0e149703f49d9534fe9c026bfe41c2b7f4d75b2d1c24cdc7ae34de382e62647e2a6adaa4b7a03fcae9c9ce87810f412646b65f0b0c649fba1f658be5209cd57b15381226a4db995e7c37ff7c62b857c98e556b41854eb634483b049d17f566ec1e19c4519ce373992597ed5ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65c9dfd3a0ff90741be882f49fecfd502138c50db57fbab42547b20a15c12502adfc4ea7f3ae520c6e43d90566010705d2586a103c6b4d808bcdcf7fb89147dbcea2d2e49bbcf5269cfd3064e44d47c164f02fd4cd024fb16e186d22bc124aebe73e01aa3ecd4515e5cf9fe561b47acc8e1c2bc5c3f5942ee0f61b4cc9d65c20;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9166b80810467c9adbf74848a5db0388337843fefb947592cbcca3c290f8c9dbc4c0afe386e8745aeee1bcecda70f4b7b9cd10566c5b861b462a1362c48b4df82f0baf4a735ab6e11fcb9a2a952e14ba163e586fe39ec92ca0721803639eae646c858a79f9dc5ba3041a3d1d8c31812ff498d4bc60948c4930996766da460366;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf90388c5d348c290e867e18c6f13723cc00bf04e6b5a956f87df7771cffcd7f55313cd4bc27f029be85d012b4b242b26f10d90b2bb24c556de445db57f842c508835da1fd16480b528c38d480052e9939fe4f0a366223f167db838de1f31c15a1887faf6733b893df9a46e42d1d03471fe10ba2540d53db14fbc523a44b8c21d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ce99b74a863cbecf24d060c76b92b83839875b4665b0b0335944916870dfa61431fca5f39e99c761458215b3507ad69862316580b094e0f15736d0407ff624fccf69f18bbc5fb9b22740f3a2bd9c3c62332d8d702b3bee7a1b420fa76b9e3844094e4f40c6e30ad71bac0194e0c95e8145c66ad3d1b4d6962aef93b5aaaceda;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h713a779838e3b597db654dbd33f5d94495c83851c649031aa945ae23c2e098bb508b120982b9515ed90b45e4b58eca59268871c4ebf943aeac3ad4479dbd2b248f6f7d738477e612a3b2fc56dceac564041003801c62d36de3735c18feb1818102ebade9789e24a777dc908fa467615a2ebebd20b170283ebee537f5524d5842;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74f6328abe725b9aab00a22783ec45d4a86a98b718703644af41b375056ad3ab3558aba2baf6829325bde7e60e1a2f42505d757f397255b5a9b40c042e52501ea485621f739639148850d9904f89803d34d147a5d0707ce6fc0dc2f414b623d8838285106428ab9ab164fa9e49820f431f4aaec3a2f542a8beb0e38143ff9d62;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47187761786b342f5a0c3368349294965930c8b9e4b8bc3489c488acf8e8a516eea7b45482e4fb7f01031633db09ad17418491e808fad9c62f654c2410c99d65c13fd50688e82c3bcd47f374fe9029edbcf4842030d4c7a9025d892e5cad4bf675cb2fa22007218db48b632786ae806eed0aa31c66a997e51f6d224c9c3f5c07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fe41ddedd4a7031ea6d3ba07326bb6825e41ff2d5b815d177eaf016dc81fae8a7179db5362c00d9ac84e88404c7b13f08e026c5b7b2073d89ae0b448a11963a11291331367553c41059a5f2e8e875293bceda4259cf9dfbab59c138f4ba774ac48406d32db28c7818fa056a06fb8baa76492e2b09ec6e4b562f757644ec8380;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4462ad1a6d4e8c515a29d231cc1b8f75281ec8804e38da347459cab554d198a9fd5093d3d2f3a4616099f326449d112cc50066899f8553268be9f4c408efe11f0243a3a0b8350ac425354d8fc338e52afc184a6025596db190119a1a11061da081511826cd6d356d8b9a1165244837f0c7564b40c96bda5c604824653d80c3b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ceddb2e9b4c5ca400ef574a88ba203adb83188e5623ea3adbb2bc99fdd40485c7328573e688f4878e244588c263b41394a5bfe80c4769113137740aba16f9f1a75dafab1c23b04989959d0f67e092c01151de71c4e727059792f951eba51c42057a7022fcfb9a2eb781675dddb6ec7ccc9a53c35588de41e1bc059cfb79c6c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5cd4aa393c829f75c1f529f3a1c4617d592bf4bc639b5707f60c33a16faaab2f1008c0e06f5f9fd8992ce2079b493599954d3266bf36d079bda629a9dfd8581439be436e7d7f0da452d4d84c9562658955ff7a0f50aa7ea3d1c9fec5536adbf9a861a6968d675e329663636da21834ee4851a5964bb2d050b5b155dee2a9ae2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34f5e08b17cd86dde781b35f47a9398b0787359fe650475bce67a46cab82e8d4ce1a336c5b5870156a208b407cba8b1645cde3eff19fcacff3afce0d5a73fdd90e38fcf97c6bb006cddc58d7ccb1bbe4c7c1072dd3bb5313a4737795b6373c3ecc8ec4e6826f5c62a8e306cd4942330335881fe29c28f984e3c0cd6f7d11ac40;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82db0e710045feb0a834a52e60d076635ad4ae543105f1b466e633e8b644efe06e2f8c33056ed5bbd7979c47682a396170fb695f047366e125cbd0218a19a353303a5a69a5f920bdec84527f60257cd6c6a61097174efa0d19b72d840308f5244a7ceb395342aabb50e536174917005a16738ab7211587cc906a89efa4b3925a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heed971534d201537d72898cfa6e651f01adda24b4db30d70ccbf82cf19277f71edc249fea56391816637b3f0db24fec1341d51a643a7634d192778693796af72ec1eab5b719a918eae5d07791a24dba62437f6ff40be9a09912ec2e155f5e9caaaabe9af6496b9bdae2c186adbe75b875e9713516171b0b4f275bd1f2c04316e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dc4881c9a62779e8a01d79ae963f218b7860218ff773d8dfcb49d81c34c7b0cc9f986ee5f8bb1953ca50d065e8b88c4fa06dc2862b7683d4375be6e0157d1aba7840f1b22487911b8d26ee8ba7b3fd874216fbe3495229c2d32104245a4d98ef51451a25cda69a42e7148583b5767380c72d7a07ed8ae68c9510b781777d942;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h806537358dde15f6fcf425a60d5d8bd8a1386aa0e2944af3e6f85ed3032ffc6e7fb02eaad8d1ffaa44059da7446400947fe81a7dd60934b7580e42926270b996e4c1ff96b91d741ee5ad66079327fc248803c4c2a2639a70ae10ba3697ed6ebddfe081f8fc233f0e94e75135e1f89be5fac986f1a18c5edc2112a8b0cdc4ac79;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc5300fe9ab6d4b965634072458b85395121d987ca1583ef9a67786fcae2573e9760a1d3144bb2047a1847fc3cbd19139bf39c643740c2af471f94af1bc70f0f8ab0572377bee17c784352e7838554cd770257b1a3f92ad95145100d93be2a7644fd8899370e89e3c3c0c9c330f022e456c8165b0403b48bfbc8f780645c5e58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ac49cb499987490c6c4547af7fff8ab60beef4ac3e59d3b87f155427d7bf5a63f6c45698353a3242d4cc02086dae49def2246d31cce92cbfdf6d85dff2645c17ddf8848e0a84df636f14e99af2f8da760036eec72e5b981d981f76309395e9937847a1a087c7c7a633b799a6d2d4c58cb6a0d404319e4303507ee23fcbf8406;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9678fcd53f5772f32675066c449b6b23f8efa11bf79292d24c6ffcdfff04a25e763c11b27e4bb669616c8f70f79845f2632f25880cd6d18780ad6ea1c00fd8ced8a7fe93aeedf9f46134dfac280251604fe03f32ae659c4d586c665852e0f2dbed585c860855d63e96791f3e6c02ed04e9128140dd0095fcd721ab0bd500ee0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68970c827ace815cac0f02a2c89d95e0485071d0bcf55c934698e538d68fd5909ae4a34fec1cc47cae719772f755a04df89d0ae5cf022f3af7d0c5187fd3aa0788df68061823218457796933cc08d0c6ec8a9edde5b0afe95a4ea63a4cc0995dda9aef959fac8f1f15aedbf6811f78f21438b09a32450e1d8bffd0cbda1e9835;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdc7bdef75ba963c8ca9f14b6365544e3eabf047587079c71c91fa2b98a2dc467bd9a14b3b68badbbe52aa79212223bdfa4652e2fafa37511a6b81dc27bf1cba3c0986e829a722abd5bf4e0558706932b1f3b7e377fe9dc0add39974efce80a5af9389e2a5bed13c6aac2fb11edf48b92c74efe1231dfefd2e368bf1326f99b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h934ed0001473e3b36222911f617c577703ff95adb9161e0a998b60d516d97e35ff12c035e2b531fe416590ce2139a03a18ea27d71f710fa7ea269f9e69574ee4444f9d17d14e254f855e4d230cd05a8b95eeca77bbbc3fcb602ddffbfd419ef6ece469cca72cc3e0e36880fdaee76b6390b8b05f28055912de5403f81ff42fbc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6af62eae317c46580fdea2c1be80a3fdefd8265d01f296ef4674a3b626815bd7dea0c40e9b2a2830c4f9dfd762c654c367e91062ea807a62627a5ae5396efad19cf18f019145948b86c9487566e4c72824dbda70ed105109b11860b51be4bd820573c1b68fed587bfcbf5f46ac408b43e3187c451680528bfb4dccdd99566a2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfb76b241b5c79d9df10353b3de03e1403cbe91040bac916f891e8f5ed806a9c8b0ce6d722715a4daca0eefc20c8c6a65a0601bc4a14528278460a2cf2c472e664c74d8aa6c1789e359e5455704866f9f088d7f46ce4e32dae8760e91c4b1419d0f277f08d263c6bd04b9a8dc5995df82dbb2750b3499dca56681175bed4ab01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5014799beccab656f6ac8e30646b75cdc0a6d5a2ee166bf17b70f87bfe8e67456861c38b379333f07efffcb43dfc982de817bb1b1901d0ce94a533a1df70cd7ddd03165c0058e1a37ec1bd654ecaf8fd1a5b5c31dd786ea1d91159a42fe167b6bdc8952f934a70dd84736419e6db1689579ed1552f362d0e20b9be097f50f6a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h144f3175fcfa2becb585eb5bfbfd6b491f200bb53f121966e948b28220bae395700c68670083cb4a295e24d3d3265cb84e690386dfb3d119e2047b6a8f191609f3c95467835cd186aaa7e3776a46ef10cf2e9ca4edbb7172cb3b14f36c8982c6cff77b776ca59f9ee3563b15849ace8e68d624658becdab82a3064b45698eaa7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca8019bdc4fa0de8a6bbff7dc7263803ce273e1238a62c66a9a6a2f960e65f20ff0b9063f3b94cc9c82ee08f18f2dc83405429946909cb056e72fc3fbe61e36864fe04bf7b869e3cd8f39fd4f6c6e927f0117842da422e492c85d93984033ba29c1f9e295fa8450ce25e51ba55001cbba063547f0e2df9375978d9fe07dab71e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd7cc261d0f8db926908131938b5ae77f4669aa5cbb231e84973f4b6ea462059b997a5e9c5d0687915d29417f4103fbb91cc82a22c2e1298976545793a93462ea1f6134543449fe0b361a251ec475970cae61d05ad5fd5b9d040d699e99bf39b968fd70d69494a9526bf00807aa5dbe7ea480944130151f2e45a5299e148a2e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h810e885850ec170bbf3fa8012fa330ad595f2e1f1a62b8f164eee8de8fa76859a020a88be90a44f076701d63b69dc7da9fd6008f0d342a2aee4f68264444b68134613140182fe786b18d4af0c5e209688173cf93f460256ada5ac5a769131e73c6b760dc95ca9b7415e6f34d22e5a2cc7858e0d522444cdff968b857aeac9bc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fc54ecb605a74ee95da523936834746bcb6ffb9cfb219a76099993d1943eb632650839bce0bff8473d96cefdb6cf8eb9cb03b063712fe76e8fefda5bfbe4cc5951bcd3a43e7c7d2bc4ecaf7d3b95ba1abee39858c94350152ee2e6ed1bc83bdfbb98519cd1e5764fbe5d4363b6226de52d82289490c9ff31497b355c027958c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2163f5bb18e1f6546d8b9ef89a95ee7f5b6d260be6eb4c8e69e83e5336ce22f54a7b040480d92206de6775870ba4d58c846d4f9f0fb0157130bd5779ddfcfa0bfbed159e076dc6e05d187c3fcca96e3e17d45524f6fd5e1c3463532745023f09fdb726eb9a93d970021eab56925df38e16b825e8e8b1ed7b7acd7a91c745c71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ca27b4ad7149ee25dde60b23d34555cdb0e68ac646b47f7ccb5839e9d5c4db28b5af84e6fd81b72dcf334dcf5e679a8c7799a9970ae46a761189bbf9b10032e1e466101ded950ec4057128b3a25b04e3f33dbbc0f2dbbf263749bc5af2e0019898232b6608f4b790e7a10ec4f79950acea80eb40c640594c3c3d8e5c4914f92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb995722b0653a4ef8fdb62b311cfc8e6a0543ccc95364f47d2411779d7f2b11141cb64a46401a8ab0682a8501bd1c588c6358a554f7907df961f15500ca5c302da4e9da33558aede56818b3be6880a0b02cf3b4d32bddd217fae225a950a5c6ad558b1b75b82c16a32a2d3e4c13bd410851d8ed8ebba50d0b282facf409a6bd0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb483a8bba086bb1272597a635551ad01c5c79aef03d9b0bb541e86f3e4a14b4bad2318f9a69f26ee049222708f5739481d4f3cce7f60047096b68eb8dd001f0275e708bb33921973d38574c3276e14673272d627c2b32be2f16d689e763d81c15ad21348972404835c122ca729cf998a85cc5880651ded0246d7179458c47de7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6729e1cbbfec5ad4ff6d133587b8ecd61de1a7d63640cd9ad2403518c3c0dfc18a254e337c03a3a01270e2f61c7886dfff5460380c9dcc2c4363c8f3478dd2905dfc7f3b00e04d4c905e734bbe8f572734477e00af971895dcb725cb751164c332b2ca7b9cf8312edf2efd0422bbc4f77e39eb6e704979b234acb303d1a27e8a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he809e7fba0bba0a07302abd109d8be98672f23563f205db0335ef8224a811d783090ecb0baf24ae3b44daaf9ad1534db3e53557753c60dc94733422daed98f4f7dce82c1cb79660b8be5e2186217d89aff4d2b0a7779c5b1990f513bc196b30661b1d47b27b51fd20af6ebd41813c02fa082ffc17b19a60f67fe48647d7ade2f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8525763bd4d2de5c6f49524d4f43eda7671fa02dd344ba9aa9b33e157b7598cdd63bcd773f5fc6f1a23f6ec14dafa19d262f1ea1f6eae9138183ac0469f0ebbb71255e5d363ed076b0c327c6b88296d836ba5ffb9dff7fa7b0d50fa1da73a490c26f7512664107609bc32e00da78b40d984ab48710d6fd72dc7200b4882985;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35def0e2a55964ccd78cf3c65974d1b5e1aea4120fbebb1fba593ebdcdb8f356562742c36fb512bc676376d1ef6e3a6aecfcf418affc0e161437b66d8ad08801f378817f16f867ad2a4b30886737b7c0695e20dacb31095d876066444071132787b9a6308dd344bb0da4f8c2a6f16433b44d2210e3b11abd6593422ce89daec9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3c43f89ecff5b7d4d607c267ceeb80e19cb5df049254ca73216ac2974cab9e34bd50697bbb9c9c384bc4816bd5b9253daa7c0a7924e804b909e4b7e2ddc411b62a334aeb795807568f3c85f5fa7ed59221a03e4882464d7f6361f80a1fab4206b90d2591ce9e538e31f3ce9a7b3296b47195f7c7be24c1ca35a4972acbe84d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf55c5bdb9b50744ce971af5c6031a890780af9553664a69eb1774ed71a83f19d5e56fc07a5959ea2b863c972dff17d0c9299d425e8692411ded6e19d6f4684eb9e513a0c6e94bc492becf29806802641dfb04296d42c5481759b623c1a935a2f10875d7eaaf94ce29c66e7c990d8dd9bc069651ade043b2b8e26a9a2f24b9b29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hada30ff71d96bc81e954e851baaba3f475dc5b809665116b51ec71bc3218967800832160c354a7e740a09b152e75a870be514dfcaea0f90973571ac101906f8b6e886b9509af3e7d841f620118bc308570e0abc68c4f2ca6059bb71a6d9b9588e6594eabfb2d8ec0c9e66bc5eda11f2918c68cb2ff5cd74fa7d192727cdaabd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79f5fdbf5cc79c2056d61ace5e61c27d19677fea20ff81db4181a18fc88c0f071d345766f66483d711819ca159121795f0ca58f501ac8c5a75977e528d5369d1bfb3d479ba9c833dd67da6ea3d67c8da23816cc5ab155c70fef32188e79bbded693ed7ce59f38440734a9a5ab9e508ab9913520abe30275bc812f723b249b5af;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8be460e50b712f9d555dd43e1fd6f9dc841f8517b6c0de2f69c3235cd46e1d58314149ef4395dff792f4e33d066290a9baca03cf08346a5ac983d95a9422fcc88c0b61c17fc1744c92fcc2a326c62037af3a1a93c300478e68582c86ea6486a90df3444dd9d033cece82e0c0d7397aedd821147ee7be84f991d7a6f243c77596;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25680029edcd118680ba86c52cace91ff497f744a6824feb72d3ab2606ad08c9a3fa2d60fd3d01d1f318e411eb664a6bf5606ace63ab1c8fe4a43bf8cd376aac110645d89f4741a64facf8aaa63e1e6863dd6153760dbfb545dd09992f14d1b4e5967ad9f763dcedd4c885a22ce66a31857db64693d529c5315c60d7d2862dd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d924149776c51e8100d900dbc81d10a881896be34ee9421df9ac041548068f0974aa78f4ddf8447c779bcfe5e5835048d79f73acec5de95148b773be550306c525f44dd37022cdcaf932a947500eae5b64e55d964391986048e68de39a65cc2d7851c273782f6c438b9100269ed48748103d20314fbf3a4576823a832405f0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e668389f5b3a5aca2c859ec6ea7af62811c0f6b8d989c5aebf7ec81f1a2d2943e72ccca27c8e8e08d254dc2785f2390265d6e5aa225defde8e1accb6bc460d51f45dc14fb41f32860c633b6a20bf4fa56195dd9df520eba5ee2ab0ee2b087e9d7dc75602ed7253cd9b57f13d3922aef6916dc3e62ce4f5212f4197bace5f0be;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc420d8b1001c8b3a00a8dd6c3b0d6d9bd73c20228b7bdda9aec50ec6f098cb01eedfad969105b1fcc5746e2989830600e6fa501ccaff5cb60527c4b91ddc7169222015cb6e80b6e9f2d9c478ef5a11890a1c6fce2729ca2477041b82a90980473809cec15addc4489a86119697a1c0754bbfe6d5a77d02f42284caaa440ea3f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb717dc4fdbea7f5bb47c3707cd5be5bc46b4d22952163c6f3c1875109cb5fd2a81393b37429f9d0bd1974f127ed3ff7b08e32eb050b129a764149c407f7d4a0cef35aaabc1f691f7d31180dc3cd9e48258b88fd7c7cc786171e9081dccd9cb975b77483033905acd8d267f87403c6c649dea43c4647cdde43f6053bd4d552243;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71066a672368f866dc524c9e7c539261a528b93ac4a5229bcabd859f65688fecb0c704592d508f87e0a6fa5c2570604e7bb7c4e8d00341942a972915ba079bc9db56dde9d6c5cfc9a6eadfb2b2a3e67ea04c678de9cb78ba1de80f7bc3fdb4de957ebda418d38689d9eccb1fe9a74109502a74efa14fdd288c7b578339d68535;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bb09f679dc850aacc1b2df66375426fb10eb9529191cb9bbf7ae03624409ef6f7b7f9d3855aa6de116b3350056b3b35a83706f1feb8002d7367ea0ba6fcf86600d999fc9272716e849b7c02723562a6654e3fb0d13463c894625ea3b59a21478d1b010adcf91d2af1e149e592a2c0ebdabd261909b2eebcdb2af6603ebf8f1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc39e7774fbf87aeacd24c332a3aa7d2b1eac6e64e58456b2e998f70e7eddcf6c6619efcd49001ceef70878ed93a92fadde0bf85339bf425fd68834b37d764844d9643d6b21992e3a0844a0157280af24e4a7fecfdcf9ee5a3555065f5d8cb0d566110907ddabfc52029df865717a2606e882764669da5b1313f71d2971349379;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2207e0e646c12045c836bb769ba678e53d1725a0be83c288e0272368eb65b0c8828c1787e46910d1d6fa4fdd31d471e8fc47bbbf79aab0e7f0750a4a21de5f7b55ff88356f968bfd9120f157b0396a1cd948af5dda9549959c57dd63c3563df5d049f4352bbaf02613f75d4468aafec01894fae5d0443e50ecfbf9d750aa8ba2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78435feebd4c1a3c4f6eb43711292c9ea8cd06eecc8df2dc9c0ddd1e902aea38cb040cbdb1617aa55eb7f03fe372ec39b19715070c9bc85e490919c994d17f438b737cc7965e99fb751ecf451590e51803ab1abb8d24fa22b22606bdbf95e6f0cc2db7e218932716f1f4527d5fb4fe81060c58e03f5ba59e1c1f101cdf0d040c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7abad1c84b82e0c45ed7c74c55d7f587e23798de1ba553dfd70980f0276901199b00e1a1e588985d900fa3c99ee8c8325f8d2a7aece744f11f857d7b177916d2a4c5a6687f97d65b0adfa2de759d77b3ea35e5cb571c214e2cf6ca854601830039dbf61674c9adbf689effb22cf0ee5c15eb8643ce1749d24edc1624c6b1858;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee1519176c97ce453c9d44e62b54009b7cb4e86a05228575b478f8a015edeef5176565b006de7abe1b3c30c8d5ba2103148af8d68101ea344df3d860f755006f6fbc370016e31a74970e0f61ed1d2a0d978fa31cf6ddf582f0e17eca675fa549d11235c1737ce80d711e965ccd5780f839ec6549dd18a6ac67d187d47221c001;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54369ef06becc026886628dc34575258c2c0507c17fd418ece9db5a35fa3cf47baad6db2493314f5f71027ba26326fc224f5f7552c79fad66d192f8c70ee028c3d5a9d1d28ed345351c78ef7076fcce2cc2c1b606b2242adff47c1b2373ad3ef2fd995b207e53c5b6a725e6f9a8e789aef66d64d116d4012ee187fabcc7c180d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2525ebf9b78ec3e46c559c04fa10ff3edc720decc7084d09642d4733a01f7b578371b84045fac2e15e8ecc60438d3c00d0b0733f8ee66795ce08b4029a56b0d53256443cbc6bf1feb3b51b2b8b725a6048c58be58d14d39f5b9074c5ed7caba490b9f09a2284ff28df59fe6b1c6e640ebbc5bd9dcf125cd374f35eaabe8e04d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb640b4abee7c4c4c8447b6d39d821af2b63e27338aa7041444c8a391d1cca19b11d2ef67c389b3440f4ca6a0a3fdba2eb1f68e060834e5f48267582bb2f695f03f7dc658ae5e3c6529ba3c544d1f39e20ce32dd1d7dc442a094fccd63043e65cbf67965df0402142657641ace559c995abd54473dd2c9ded456879df759d6c9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdaab2beae68952dacf4b160695b68bebb2dfbb1f26633e2a25008f8c404b979a8a563a5ecaf713e1282b1853121b2aa9741375e2cc933691364448a2f5bc8d6d9fa50b7f9a18430c8a0dc0a9430b36251e5274061251c288d7b8ba1f724567203917e79bdbc0d1e088e41bc69b95fc0691c9c3c552795e1a650ca10fd01fee2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe2e7563156e714323197bd9749c769f7facd34975d857b3fb2e8ee6d024882020af0f932d940790277d57b34d176304f8590a22fcbf24f8c0bfee6e1fff2bb9d2a2e734183fff9db35820ec23b9c6b917143603d3448744ac2804cf6c6c99189e2be732673fcd1e0db97a5135096e7ba13eae007630e67d2e7e94031efdc21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h138b4e6d501250fc2952546cf510c07ee116bdfcf0f8207ae6342f280375bbc74ec8992cad2be1e1564ca056bfba555a5b8a90d23709f08a6edc5e6a2502d1c0acbc0add7a3825f3fbcf08f2c469e8962eaa0a1aedaa63a0d029868732b4999a2bc0dc1e0c5b467e7078bb3a42706b7531d1504144709a405e5d12cbf65d57ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cb042462648552ada5b3776c937b29debb798d93bfa16b9b3fb085b079d67c9120642388890ef51e54d5c289d7c686a6b01f4d338c8f2e10127c9fdeeecc44e84a5d9ab6a7884f5ef19a95f1b7485e2785404884fde9dfe73bc0adb0e4493bd863484de03afd5acac2b3cfec311c7b383a7bbe2dd009c08cb6f2e675edad6b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h125cc9732b77ed44e4c28cca111fb1cd7a7de58d05c916691034e488d8b91afe677019005d621a3679eceb666ca4ea5a16bdee268e347f913f1439b277e041d839fb145d0c7308ba6eb6538c625bd425f31c2931ce92937e6792c024f2c3a350fa7b81f14c2836ddd47a37997813f76ac48212dc07f292a9dc587c930cbb9d64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a16520ff06567576b8b1632ad96b8e90f05b63b36ee6d46410aca7709f0f8250bc693dc0dd5dfeb743d9fa7cc137783cde053493d58250c9ac48c239c58c958845c30414f44b1e350d610be1109d86fea05011beb424d0c41f5e632ff912f0dafd44ba4dca88da0c8a0d98a8e50252e280630f375e2611416f45f3f299b660f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc36b17904c42a96513edbda4ac2d188745952995d1a26991c9393cd52228c749b2ddfffb1c378e08c68755fc1a4718b57ae0da64b6605dec4d3ec82b48c9eb20deb2b1d86e32682cde5e447063b7bc621416ba25f6a8417537a75255a6e8ac52f3c7a63369d60248b5ae12a9ee514052b1c4fb95c9464daf3c7f3da0a470fd9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h459d88252a40729d8f724c739b56d9e454e138bde7de190e23ad7335ffabff758147a658b65b57cf0989adcb3dcc0649e1c8859c9b548005e35c648e39b192aa6fed3b745fb4819d4d3bf67b3549273eb77dd4005320179527d8c35525ec3c4a74e1ed5bfc435a9154deccd55ede611fe21b5967b1cf511b70c9350bd3e35f83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h195abfb3a239c02322492e90452807117c984a102e2393d7aaca096d61cb9942ee8b6ca43bfac175870eacc8395e0174928060d723437dd09a4211ab53835ba96450f94abf63d5d2d8b45deb2cadb3ff79ee86248614ee64ea6a947aff7087f3e0e2421e744c357fb3bf462f55fc5644a8d5decb194d62b37bb2799fe5a11bb5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef580dbd0eef80dacaad21b5791e3c277c814c8833eb081135ef90abfed8e45346a553c5cdfbb08f4f7db16a22cac00cacc6fbda434ccd2a449f1d6a260c88f1ff59d9ce2a551a31c423c42a11fb9ae638638314656da40006dd018456251f2d7f578eba7a626bbdc906a37ea6dc791a4d7c15937223aea76e6b251734a9ef8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c23069bf05d2305a24f0fb931615299e6899066688f64277fde9615b91aa11d212c035b4e13ad9de113c646b19be5b8a1f7451702d36786dd4b6c6aa24812fc58c2ad2a4f5fac7fb12fb789e5cf78f028f7d6c95010d4eaba6f93281be8c34f20e7dc80ca5e43b4496c86a08030bc95778c9ce87ebb226c9cc7a5056e0b711b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5b14ed5f7e593cc104e009c80f1bb111c2fb694533aa9bd32bae9b106d2a4a52d4c30ec4c44b8f39e45684088c2e563536a19cca165ad220e0854b5109e69be4beb6ab744c797829e89d2efa1edeff481c27fc1b4b035d2113407a6d369cfd211b3e525bcd3db55db353e89c2908014ea7024490a4b542506c94f17aced1c82;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h776398669dbef822fa77cf08cf5451ebf7612b631fbaafadcc46b39ed1a0bcc8540101ee790e66d026d0632ff68a7b5e0a8f008ab81512c98900ca803f5e74d7e4eb1cb9077bb28c67b730d5e399b4ed26875927221062abd84aedf98373842fa06c6c7843f66022fbd5c43d608ed088913d7ec1ba2ebb536762d91c5d64dc64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f2601dc6320943db813915efaefd76ea0ead4ea1f5fe6739b1813a5f3d67199efc9d153825bcb30b0e4c0eb03ba79633a20798a5981caa659a6ab12dd632ed6b2159ca36fde384962dfe7481ce6a05bcae1a438f10015fee1f2c10eb30858c346073ebfaf6f27241e961b763849660f8a06c0d06813280a5b45522416b12d7f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59b5be10fc9cf0585de8178244a74b91ba6b0ea5dcd3414c2631e0494a1b767f5fc11ca2394bbddfff198b056b92ca590cc1355bbb753568afd61861f43f517139d8c234d3e08d091ed53a52c43afec67515091bea962dd0b745e1c81cddc42abc3b8bcdbfec25602a8871d6802fcaa499b582acd40802b42780b92a63e56077;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96444d2d86b72e3d70951930070d123bf1cf73b12bc35b0caee5180178c4979ad04b199369c819e47deced0760ad596b5f535853b5d43c6ccc8905fd73a370cb3c454720a889954156114b76776c5ec4691f6227563620a6a8b02e2b7156a258fdd2635da01d04a3ea8b95051809c775cde0f8fac60c3870e3789af103ea8ec4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4214c8921469e7ce8a283e5dfa0d38d6bced119086484f0194c41ba46a4629a44a73a958a1707e6fcbcbc01ad21501f9a10c2fc75ff1ebcf56f817ddd3c22fd6c337c9489f88586e4fac455f9a0053997ffb32d0a1ea0bdd3e0781397c1751051b069699ca5f7b2ccaef90ea74486d5cd911ce4d0c7f3114f186180e0889370;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2271d7abe116a8bc5a452ab7d7815a411b25d5de89952b393bf06dc1e4132ada059e76603c564962e7f7b16bcd0c963e2a930475fe764172b85bc086258583885b290bc304e973d9782212fee4f2ceb37ca37eedcae2f63517722c66535a53fbc9a2ee9b70be69db0a79a1e18e02940e2e4b5b04d5dbcd04c26ca48c0360816f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfa4ea05bdf2256d552c6dec0eef5eb6e02ccb4d458e449989122c7d9154ff707c737e47a83a4fd92e6a974bda31d2461c8defddec133f425650ab2205024f74bbda2bc276030e4a84f2fa4d86d6aac91eba98f1ed22049c8e71e4de48591b99fcb7fa927eb26302b8028d5f9ff66737ba779987daeb76f43fcd6eed2232faf5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2920eb9a544e3d547aedd81e4a3c910a4285ec639fd90eff595ee67e6a8e7c32fadaf93ce3177e65f50631dda46c0e7738ddc1060eb00d2a71d39db1b43914e51abfad82a2c664e2558f4c9599e7b0a9d32e0b8710fad78f22c3b6571406cc8b9439c34db1b597c48348a5b12a73e1e30af86f3a61063e67f6986ecf31c24fa1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h385baf5c9a5b78a5c349e8584f162a4fd7b1373d064ea7a7f89da6e687d403dabfe94c196dffaba48c1d64167cf6061a542c2f91a16627e3c1adab57b39da3445f95a3d56d3bca2b3ef6ac0546ec105e4ad4680b3bd43ef9113fff861ae34e10f44ee91fd4059fefb1ccb2adeb1d3c44606af10fa9e50a6fee7a711d44c7be49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha92fb211504b1ecd3203f260af7e04f225d70651500654d6550cba7e4e0e7ffda7026d69d838429065fee3bd01f637f6b2b596bf8081fefeb5c7611d32767236603759417e319e65de9deb09b61b4301730e7fa247c95b346b9a763988446c6df3bbce3176956d5bf035f14aa1806396dc5e87473a3fdc077e60476f718ae876;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39135ed83be48fcd9efdb64ffb635c5f282e2e24f42dbabf4e6b29451b348ab68912f93642d2fa58387b351fa184f23dc54eb8c41afe64670f3b30081a1bbc340d9b135dc1506b86f81603ff7871495495825601b49b2826d6adfcfb9bc071ef0e5aa4626cfddd8afcbba89c51f104e76515412ac23a5cbb9e06fb731a831ece;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51a1700aa65c630486538efeb2f1f4c11d9d72131fd781f76a88ac5213f8695a5cfab133fd21bf91efab23d295d21d334f7137f060046cbb3a02a2c9a496d4dca214b6d4ee938b6b824cb2b3cdf79c9e4d0281d0437665be49c21466763aa96b2e1dbb08608d63d85f06d1dd4d1ccc01e945e758f9b9fe2a48c6f80b009f4017;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e3ba5046ff4fa651f5a6ca3d410e898140ad900b00d1c1635074b16647601ef3e43293d81216b1f58aa32558294216ef6485825393ffcb5e54d5318b14d76bf6d49b3ef5c80a6a8b0e3a0772adc6a527d2df7049516ba73015e2daf9b0a636d4a1f9a37c2d13aebeb5c3055cbb78c3e35a147089163b11aa6bcc3a79794195c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e012f5b1322f87ce2a1b0f3754c1c4c49a0355d194de4657c8c628012af491a5174f9352eef58ea71a6fe2a567870e5f2d4c6749141e8cabe8894857362b3f676710caaedf270cca8231fbd5c91e16c673c336a575ad37a3e13ca0830358ee6bfc348207a6b64e015b85554230738e38272021733ab2edf008e30af28c7d92b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbe76b911a2e0df7060e5df850337cfffeba4a328ce9d402e9078c253486ef94ff76b74e8a66426bd94897d4fccbfe0574c4ed3de039127b904b15aec78e7a421802f17c8b34c066606003badff0bea67ca52fd1909e57f6675129ac0235164d0376c854c6e41890ec0f2740d00863c62b8bd46aaea7a951475c401c78a42d5a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f87c8c3e3f67a4235bc5f3aa2f18371ed85fe1dd389b52dbb17883a4c3ee2d64e831bb8b0ad6e4e01b926b3efc93c4c5c01b5f158a87f9055555685a975058946d7f56bac44d96f2b79d734e52b2768d7898ad3817195cb6ece847b7a2f4ef81624cd8c3b807f27f0358acb114fe16d2ac097b8babe7c434a9d7339ee39a54a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd42b9426ceb01656208da99633c3967dff9382d06fc54689af4bbdee3e8868a19f6f97f8680cc4ca78bf8f35e71a2682b383eaaccb1f5383a89b0905a7670935b03d1104164a838fd0489032d383c09dc0ec9cffe2835197b66a48507d1c8c8a077bd48eaba36e9463f25980191a9f7e950274b7d32577ed6d22ae98f6eca9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d5a53d97fe11f035fd5e8cbbf08cf4e787c01feebadb1954052a563a7a19c8da43d9a7ab4c884154e721d67045e28085f790cedfce6fbd2e33ceb4cfcefad588684b714d6be55fbda8b5cac9935c1e9fc5ca68f167dcee41ad0b051c1fa5087eca3067e575f4fd8de7e9bb90eb1c8dad92dcdf32a95e6ba1f91deca23887a1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea05bcaf7b1d11bdeae225f3f3d13a2afccc581232b7d5a3e1ab698747c4afd4b1497a8fdbab9a35136a20dd4af695d651dae15cc7a3dc438fe26c46b0dceb2d9dabee0c8ef9a73cadeb1525a433383a3f4cf4849bc64f18bc5bbb3a82df89f7b5133c960b9fba662813f03d8f5627751209b22f313383b52bf7f2b174146cbb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bb76046274abceabd7643b52775ce099ca4bcdf482198f8fe833acbf78fb7d43f99cea76102783c9b45816c69af5aed89cff7651b6e21b1bb296773caf5090500933880c0be2cd4ebf13bf89abf773453892294c17c108a550964d7c359645b2a9e68d23c304435f0c3708a0aecf1b95a776f672d0257b1024ea3e7bc36dee5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcab4cc43699d9e5f25411d5d7d807e235e8524aa30f2958b1ffc3a7fb5c24bd7e2ae8a3050b44f8782cef2a8e954ba66abc261c4479a3d2aa70e1ac635d59dd74945ad75cef67351301481cefba6fe4062e4f908b2d32bfc3c91420a4dc5d06894317258c78c29665b366245cc6ab63c900816f6609c346c2ddcdd71da48a492;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d49862bb9c71432394c08acf2c75cffcba31df42411130386478ca95844fff4fd5a83905d6349a72a61afc0a10f382a15987bd9523894862cb5d099417af42d5ab2bd3e60650231faee44035ee3d69bd073f9e842c58e7d538738bea55d717d519d1c56b6c6b99ce09aa49034c6e65cbae2fdda84af02a7988a67fa8fb7b03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91c4200f0895794f7fd13dc4501e0aa818b47e0b4bea33c9c631fdbb04f36809411460100ac95788b6177623990bac1b9a3a2837abc0ff643ab44aa74817802df196b1ce4e93e42e733a4894232c6d76659e803be41800f5c8ce4ac43572412f1d9617aaee41a00468c09f3e60b1fd8c0b42dd70f9b35a700ab7e8fcc2191a85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd92188cd0e9238089fe57e2ea6867625ed5ed5b6c43f16e63d9c2c5f0a53f066ff8cccbf24ef87797e4dcbc39a0bfee4cb13849216f7a13cb99278542c875c6c1bbbc1dc525e402dcee480c6ae571af7a06933d542e74127f7c0aef284d2c22183b3d1a77df479f9752bac76951fddcca61cd41d9829be7f1482bea09b17bc0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c7560ceabe9b7ef9c4c5c2a0eeb3ebcc217bda07cd0179b6bc1c4b55a870b93e299368f5a2fabb73641a026aac072b250886d4a57a2fba8def90eb933b8d6a17e261d1762817ab1019c17a1dac7d6224c11c1cc2ab6d549794a860196dc2b7cbf48d24aeea9745d579e4a9134922e36c2507a71bd06f1c581da870689994194;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5de77c94caee799f8fa8b7aa5d8ad108c2142ac21063227342feaafe2876601ae6e70080c7419a7d7e1628108677b8dfbaacc64d5f28bb86fbb2ed8fe78b9377e0da78dd20ee433d313facf6eb1d86228293be3a8483ed379b4976eb47c811472fc131da6642bed8bb713477f535714cebe5b46dffb2c3742d5b8b83c186528b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfa77c5f8a9be0b8049c4fa752d82a14189c7421ab6374c22d169a2e46f81f6ff562f72926f177ceaa54388013156d7d600b4a7d453b787c3f0f1e547acbc59597d58c8bd975baede2bcf3265ee60cb937c488767ee6180b942e7bce9b284df86e5529a40d18f07346087a09d9eba6d5c2668376fb92dce7bf5159042c4a3a47;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h741ff0fb7ed2f987199caada014894623122c15416e08d5c0b3090dfd646e8ba54702e08dd7387e1cd1a1924b79c388a2f752a6319161b4b3600c221f55d3f3cbe26446a14222e9fe892154d5293da02b6d29e0f50346604b0234e06060f94fd153f9e72bee51c891d76ac186baea52463c9ef12782e4d12b71ad7c66ad24f32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ef68db5b862e7dadf959e08606bb8002e72a35a00258fe41b16fbb7f3e1dc597876e9ea2a781bfb897304fa1fc5be1f456a30a263d0d861c7b05cf25d5faa20a9058d90464eb5d1831060c6e07d7943a64e005ce35f36c544656705cd9c8b45c843feee9af96973586b2091216443f2665bf4feeca2978e601579bcb8f2b6fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20faf550ebc75a48ebfd5d7073b06589ccf7480abb862f4071fbf1238c0d33a6207f152ad33e11ead4c8c7ac35272b3e5c9ee1748afaf32a1be32000801a7b027f437d8f5487b9e14120fbf7e977d9e56e27a556978316fb55ff94012e8c9ead9c44a46ac2f3f5f95f58a38449e0665cc8630d825af8d553fddb03701a376d59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36452248a2a9a0537b20439b7f8cf15ae9e1e3e7e6835a3c6fb196a0ae8a820fc63418fc2a0fc1c63ebaee3d9e87a68063fd1ad60ade0f0793616ba5449e12373c75888fbe761e4526cb6545f253ea425876d128a70b88a3dcba7eeae70dce8e1476508a2d987f38a80459d1381ecb2c866b67bba856c19fd274d6ace08d4623;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc58f49e5fb705128e0253650ffde2dd4d2bb21f9ac56d89835d4c938f2e60b8a169eac981f0cd55a91f4881eb5549fd991ef98d307467cc0cb272f0d501f7cc876e619707a2d206055629a58eebf714eef7a6288c6c57e81da22e7caff067fe91aa8b629a4a7c90da75ec9523fe9161a335e70f13849f9a33c39f34571c587e8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cf0aec55fbc66f08fcab6a8d7602e189a9d92ca15149f3a0098551c3e1c6f4c69238d8129c99da98af10d4adabc6517e1c3fcd67208741db7597f1d0259440d2548514f693d60b9201af745d96c8d1737b9542a44e032f6ada581f1f23b641e22c4d42ff48c616d41fa22a6d5aba60a90ec6fce21a98fdc1dba638860b08375;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he34a56df1862c8ed4a3585254b25405f0da40fcae686685a7207a8bc97bae81a524f9f88e357f8eeb6d8fa8dad9e61e50fd6294e47e4cf63e305311cbbae3115ad9a161a99bbc3be22609c0abec315acb72a1d8f7fe0117b3d04168ede76fb6c48f8f00ea4ff6a0249a2040b8b0c263a64cfabc4bd74f9c065a0b5b43eff761e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0140288275605057a483612d56b4fad63e402d6210679d70c31e267b5b5b058604a5655baf048fcdc83ac6096e0716223271c5d30fac6f49e6b76fb7a103c245b1fe37c55d8a7ea1845e73ce8a6e02100a1e69887e992cbe7dcb71842b77839c2924e7a67e3e4cf2e94f950dcb71db2f514fe612ba41c89dd0c7cdfb4465f7d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d24751df07d53a30b3804a33f0a343415801039c6c4bcc243c7de39b932e1ab75e75edbed28330b56370a1a9d383b6b8d67c1470b792e818a162b5cca771d97628a046974368bab37c97f1e9f1db3c9ced359a82cb85a9acb05e30aa69c2f21af2db7f3894da3d001bccdc6da1a74f9046fa6fe04de8ee764689d55b2d5a999;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55f4bf22d029f97c86c308b85cb535737dde64aa694f46eda667f07611210c3efe49a99c9f84eaa424eb060bb5849779dc911ffb9e804b1d72ab2ba25edda4ad0d60195e5b5d2c4e3bc3990fa1aae8f21bf6fe13c8ca63080a855c9b7fb69b22e95f6d87be6bc3ad644c8adcf6a984461e1a41b9cf565af857417a7f26fa29b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba3abcb7f5c0f5f3f96c621cdc67e781c0959bfb91c705ca11fb00e04d5238e892897cc997efdce6875398619dc4a14c615c35df047f8d7c8f6e56f8797616f05bf47c08f32d6a03f2544fe73e6b45dde3e0c4969df20c2c5cd3f4ae712938491c48c6fdcd563298a29925978dd6a7150532f885f00369438279a0c127233faf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f0b14f0253d32fd725fc3905eb57662fdd0279cd9dfbfe7a58524096d43fce6b9e99315b8a1d956fc3dd8a258e9695e55d98ccde30c9a9d8aa9a619e4e75cc3c4f6bc6ea5ef58b84dcdf89cffffc261fa99d00925c049f76532a835849ca301cc1288ab68b8b93a3f214ed8eaa2ba4523f0b29723799b3ce0d5e513d5abd926;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e20bbdea2076a61c59a7a873dfaf1a23f3281e7e76e162348c8353facb9e298040f04bd495567cfa43b0ddfc23d66f7a1802ded0dc64fc029a1c13c2af2cda47d8d19dd2ac59f12bf9755ae346be64dc831adcc29a7bece69d546d35d81cc6279083d0de16edd5fce06cd011dd8d614a70b15a7dbc1521f81746e2919b736fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9ba02e96d81e525324b592234489f21bb16ed33550019f62c69e1e05b93b1f842871e53ed3d197a48879d03174317866be5ea753f91d3e6c681f9c257b4711f4e3fd10dc16736bb72fe02cae696e6a9e5b473df21f61e1084ac4c2f89ec01610d0eb6c4d293c1509a10d81accae4fc3df0da459d480415791e6265c62b35667;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he28a6d148a65e1fe2baedc8390d4d57d7bf712d006feced1987ddec568d6cc8daa2dd5f5bc9b61d99b938c0118654226356296349a6588696697e22b307f362ae34cf4156adaaaff2fb6084b94c7bf5687a0b86bec65d3c5873b26f447ce0a4a032870244e521519979db5d22c1d695f75131bfb28bfde115cf164cc449b97dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c914c9e8cfe51871f24c952677b758ac9d74d1acc33fd393927f08a754b4e30be46511f68319bef3ad6efb81c4be5a54ff12c288ada7a4a63a78cc06258d63f4b5063dddb03d7b04593451ffe18b3abbdcc438318c04949168c29a2b6219ba0968ca5a6061201c01e7ede40e06c4a0d4c2c653ecabc698c41dbe689a12e154d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0dbe97097e6d68f1d7af95fdc3d6732eaf878ac2883bfc761f7b5c9ab7dcb8ac178a3cdb1a86e13c3a934d9c40bbfb6f33c292ce69bf983dd751ded392e97529fa0d7f1c33221e42183821258cf61503c009de95f66243a29f347b9ca643daefd77791fb7f389b228a103b0737f4fd57c2ec95d7476bc3d21506939b6ed5647;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6a0849ced42fdd00d1aeda5655a8bda392c9e8337f2365d05f525dbafc8137cc16653c18183dd1d78477785bf8c62059bd11e1c4124c39de42ea3eb2e221722c983da51ec58ea2ae1423b6889dd8d95afc64191573195f0d69be07194e018a00c587595d62de1a0df23ffe223bbc5ccdcc11a41c04f815e07575bd6518c72c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9ed5a3a4bc454ef5559e8d4fa894c21bfae7056ae9898316f9c99e990ce1f7c98a2698e4baef4dbcc1eaf7d5160f3e3ef312555fe8c0a5203abe98a9ba1fcfb1421551f63fe465a4d14c5fd8bc0de41070c2de160568ffecd02d9318b33e8a557fb5cef8b41fb6eb0409336b1cf1181bad5e1366f02974505c4b09af755aa88;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21ea24e0bd4c816b8a41726f02bbd691d700cf5d1bcf68025d6f92c98fcbfd82cace2bd009b86bd0ef3ecec4a0d816acfbf9f2d92f3554e46f358d3631b2f846915883004f218a42fc254b8185b408c3f4a2ea7486b9151b5e7e9808306cf03fff721f1ea4716586abbf65bc902b093a3dd65b71f454a1f77d74b8d142d023d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20f5ba7ecbf82d9bc266515fc643c2f5c66b44f958de59e9b39ab45b90a162d14e75e472bb5c06c22be45fff95f373e7d7c4bedf67d6672d154ecad354dba88ff0805bbde9f0ba86831a1e38f65e572b0e8587e3fc5531dea853e50768ecff3e06b8d9dab2bbbe32355c25ab983a24379bd8ed5847d1c31c8cd52f2828796d47;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fc1bda98346e7f629251d7fda94b4230b0ef09490f40da8216e55f0de13b9edea97962d486b8a1c7370c991c74afb6c4143793ee12bb72c53af2f38eb0603c628f081b273c45af2673495d4a8e7432c42153a265ed4a6633c566d5eac9e505fe84daa916890bd082fcf2b92962debc57051e1e84b74d7aa69a15c1d45b0bf85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72c652e12216875b05ec50f7021c007c8d0dd9e0ebf030db24b15c57cc64debd22cd38dbc4063c2334e9fdf221d5ba6196cf5003d3600ca5ceaf29f96c6a4b9dcad86fa9ecd924df12db8835d3fb1c28c60d1a02ad4b22af051d5a1a4a85bb32dc0ea4c1ed447f29131cbc2c6816a82432b9f091aad015c15dc9f7142fc4d37b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ef2e82c7761ed218432805f75a4f0625fc42dbd8a98ffe5df2c363a0126908423229d45c2e5ea4a7930f3ce188f763a830c50b26cc4b114d26760cd96ceafe62ff2c17660d74056fa885ec6f67ca74a12df0b4afa4957a67f648ca52623e8c83bf29b1cb71dba6de79109d100445020b6c90d843d24f285ba3e73a5fa50e5e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2bdf5211d20f732736debf0ee76f11260fe1474ad1d7413e2425c920a597dfddbf9beb6ba70393e8089602dfcfcf60ab061f7e6624eef6357a5d9df8f3d66ae2359750e5298a5f18b2f855f1539595a3d82064453193aa17d812e6304e849954818e1ed057ea4ae980f8b55aed71151542f5137b4875d429fa3379a94374e6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c61e300b2574bdb58c82c07b68e3f197ee090b5bccdb5b1f7bfdaa7703ebfdef6b2d4311c46c76c846f4e88e686f07d9c9adcc08a56b786812bc1448fbab828ea9770b6f43dc145855b0c1909543dc6407015c7f1ec8f2a9549ea6568c45db1f45ac9a6f7b2baa440497d0f18b57caa2aee2d7266cc4ce9e3fcb93b29e2519b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4228209f0d9f17bb2e96c56288172fbdfdc4e3c9a24a581ffcaf1746a8a9b27e35e354c87d8f15f1c2f52f8b532c1259bd59bbc02b6262a600a4508ef8ddc67e53a40647d608de706084cc064476cb19f5337c0de5a412e2fe442aa91a9e133db0f90b058e0b3554082b36a5dbb97c89c82da2645dfcb6484b4976bee2032c77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c2d32542f46e4331a6c35ddb0c7cf56bb64766a65f818f53db224367520a0545073de906e1845f6fddf501531bd19489f4d6a1e7ba20c2ea027be1be915a00685f2033c75bfab514e742bd829efa8e20391436b60c600c69d304bd8fdd366d051df4abe0a8dffefd626515709d15c26f20ecf8b439a91a285fff186e3b45490;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c2d80aba72c22208256e90b185e4a2c1be33692e7ef6d4b6dfdf0ecaee25c916bb9d6157b6c916e54e44170fca0aa641ea7fb46e5254f44b0b4e5dd6cb5f96fd78b4d100a2ab30f710bf69d71af8da8f6bbad46d58873e923b2cf11fc185bb90aee024e33218ddada35746d9803df40b175c561ccd8fac4d48f039f18866389;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f6175ec659eff139e5ed748f897dd94e6eee5bc6748ff9c8bc9ee67bc7e7304c88e0feea5cb583276220f6686a2bc4e11e95e27bf8ca5232d776e5eca45a64b5451f9e4bec88b9cb6d8339e8421c745ed7d5d06111bc0111c7b8853d438a9e54b9d0b10b4e578d6b79d6243da74fcd748cdaf25823db15f6b9b5c38938125a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80138127608ee6dceb1a8d8d48a56a93df50aa7493eeac77c9c50047e09e01491e9f0e7d02aa3b2b1c9fa810143ff9af8e01d1e111958fcbd0ca105d9822fc70fad30d2481790cb1d9e1641185fb590e1fbc0be178894ac43fa53e49cce35dce1a43a2712afd5c8774fbc3aab59a85f2cec5db9d36a37c98add34945d0027900;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3144886e4ab2b411733d6d73b4f681043291a2551690e44a74a1170c7c78e6fcd3e212dc8ba662e8c700a7683374723d0cc2cfa2fc645427559d8775cde8033f954788ce3c2f4b8fea0acb59c808cd574f05bf0128479ab8986e5718c9d009581daebceb90cb050f9a724e6e47046add09ab789158f71d7f2e446540c5370f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb45acee13bd9f25a9f1dc7cb1d3f71b012ad9be2defbc1cfe4cb0370f9f8ead783900c7cd5dc4fccb7a8ee42dcd2c1b581738cb82a1ce39cec992cef2be40f9e5d0a1f537b0bbb7c21eb2a9fa36545844d17514abacbde471feeaa75a690189fb11ad2416e4b99733144ffd45c1172810058749be5c00462f25c351aaaf98d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14b9f8524af10a067998200901a98320896425230d0ce6f22db3fe3176434b7dd399f5f7c7ad61ea1af74bf2d093764cfca203e01fc694022b4e7e577e409721d93796b758434fac05898b10764dfa93cf4ee09d0915b7ba7ad044bda9848c7b466e1acc6af92f2247db7c87a49dc47624a9bf2255e4f2a39051e8ba27237474;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8363d39f856144ed8e46dc6ed235f631e4d5308c74c43a1a012e39188590d9bcdefb9908c9092a92bda16372328ddc33c75bee075adc59b48ceb5a0f527b0719a467ca213ae2ccf28ac6688ff7428e379115dda4064c41673ef445fe9b4935a0b309af34892aa30afcd1a50f8bb988907bccd4f8d711c5bef4724c541a6871f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b9c10c9d44c911843d3a1901b8479304414e38568286dd600d0800186365c2f8ddde4d1cf70cf4a041a1b288d91a5f1e8f5aba89341d44d2a46b62d8e82f26f48a0aeffbf0c13f75151ac900683174ce81651fc51dd9d59a2a852d9b7d9b2e9ecec7d7300c1229a08825e6fe62a1654483d7b44d145859ac2c9342bfd12022b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58a4404d599e1b98fc6a36b8f329876ff6999fd970acd60db56f3ad1e75707dd11cfc800168258aacb2ac80e0575e059e178b531c704bf9ca52f2df451744ae277a4a9178996fe34fc0db2cb3a62526113c79118a058aacbc0a7a34cc819528fd1f2c63f8f77e9acf678d5e1b22d4552999904c6290f17c2246aa51a28f00041;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28167157a6bee01eda4574cd910709eb2a3ac304d90822341c81d7d7146c43579c5e88d62d6127794a584273e43aa01307810d64a5e678ed12267be45b07739eb86829b626ea8b02bc382808cf230e0c22d19c9d0bcd042c205f653fafcca0cef1f6c955996c5f40f357dd219faa986c81443ffb1deb17aa8535693eada825ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8e640c17a1ed81734d7c452b3f4bd6da4a45b12131d78c02a4ea7a9e349df1f1c5ee3c19b0aec906add0822afba6f3f204f1d26baed1deb336d151ab65db36ce44240eedf65a3d26a7c50c9fe41b898002abf55a9ed8be5c31cd9369151bd170c9348b1e5c2227c94d752347f83946d41323a2eb15dc23a11ac3f78c9daae1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h866110e49477c503d9aee31e1b1542ca92f90c2faa4c7ee3c1180ec58c2e5ee6c0c9020bffa2889d54cb8d89fc1cd363f00dc8dba530bbb7a8cda09c94d93985f03ccfa73d2c5f5ac83673997ff084b5633642b3089be5acea4526706eee2385175c10e16879f655d952a0fbc2c0b146c25dcf9e63c092e1611dd615b12b2448;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha521d0e51e115c6d438b6075ba999a9cf980ad31c05b93807b4aff64e4b2fe5a394150cfab0bd2fb234575507588574d8b9698b5c350bd3c9d65b5a7224f630e1f70e49374886509930d7a3d9cdc5b457f54ede7eea8b06b278c987feba36b2e5a578715bee2a92b97eedb06aee01b8156d61fc07a0b0c3b68ab6849af3508b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99ee54c086dac216e1986d4ea82308fc0a8384a084f2fef2639526fd55b7712c892d6559599ba0344bc1a4af14dfbb76fde528bffdc2dd7e69c5915a18c5d6935bbbf8ac2e2943994c5de3b5d593e66e923f391ecf3a02f924d65e5c577d27bd64492f409b70ba97d6429cf51864e55d276d2a8d4e5dede8e5e7ed38628a2019;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1c8bbbe971b5d73a81b67ce99f0554cecfc2e8dc127e022290e9b81d1815a7368b0f89bd3867cbc7620f8a6ccedccfa5fc157911e33e5f197b9dabdbadcd42f2485969ba71c4a390f8c717b3592006cfd063cfa8cfa19a9362f8af73dd55cb15025542d74c4034e6cb2561cbe4d2469d6388c40bbacc78dcf387d328e2516e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94e467efabb0b486707ced2001872a4875dc0edc9b648e7353ba656f262b258229a7e2d8595fddbefebd719f442f2942732d62f2d3e8c34172aaeb81953056ee58234e1a7f3959fe4816d9859f2347dee1fb5eb1a3ff322a6712548653ef84dcf6980595871282f88d0da91d9b983c59ebad750c3d5632276f32a21fdbcbc8da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h450b4053bc3f9d20ff8ed92f4a34f1619435d52e9c0575b146a6d0b28c4414aea05f14c86408ab1c114e097ab2ae089c6a1a5ac7e0cae09c4c7aeb05f72119561bd2326493190f2b6f6f98c6b8e00119d0f75f44ce80e5903eb14393aaa2958733702b8d14e249c9859bb908150b2aa22ef0c1a4716ad8a68254b52cc45561c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97bce19d1c96df9ba4481c77e6668d6b3ab92908e7d30eeb21bba9e80e2b4e68ad1bf4fe154b38fd2f0c7f18b21e014a31edca7e8f35511880d178d0135b6bcb9b185467fcf09cb6ee491e3593e92bab2be5bb15160b4d272080768ba3f297c91ddb5d7ae78b493a291abbb99a69b6c85238abfc23ae0bf00f2ef0331f16e401;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd187947c8ee6cc1657a0b18c371fe80ae2330eed4572d0802c7be0dfbcff2cf74a2cb47cc0035bf1b567a13ebd694894808e8b0ca723f7dd975d8b06048e379c33e057c2181ce522c7584532276a3b6042b782fb80acb726db99f52b0e66682daaa03b9eaf7033cd4a758885b2f05cbe9999ac7ffb6401de13dba9285fd0b96;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha62351328e3eec12c4030619295cee47086c6ff157610785342f358ccfb7a074940f15142ac7ff36f54ab516853da70125cff9529adc9fa82be08f8effa706ec1699c3bf9e5b668240e01214b42cd284d098b9b070abc349c61e864396aa8c67c721484ba2e65d02667557b3a7f756d7ba2f93377b64f028191c48950aaecfec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb857f39b13993a2d089fc09f5482675038170094fb4d9bd6a744171d2950e8d4f919bf320dc67573867f926550d9b103241d7ba7eb1cc840aa4a6352f2c0925c71815e167131da27f422849d9cc94a6f5e8e971dbe6ddfd99a48bf9242b44ea85248f954dc5fed810370b7de842b5d19c00a7efe2605a6430134cbde8456df5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0f84c45324b389970effb4b90599f9dd850e6609d25b3d08a2b06a4e7c74e7aa4bf75192d92b3aa28397d6a93ad1aa2386e9b86f1ddeb0b7d8ab3e15cce2fb6d9caec0081f53007e0a383dd53fe9dae0e4dc70a4f887a499f77528266140baee3a3228cfe648474e52747118d5ab9bd1315628b8f4422cf074903b727421a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he768519cdc666fa452c9fb8f76942a7f97a08145013bf80d4f709b32f24e5efc90daeb31ef23b89ca6db956b808753f8e1cc4d445c60faeb009c8a7c1891273eca1f68e33a1097ec443ebd14bfcbb061b1c15eb69cf690626aa8adf21dd12a9c65a4085564ca917ebbcca8df865d92881768f716c4a9d3327772ce1d5205b08f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1f28ccbbc08a6c65b59d5e28e481da7f1de762bf69b9668faacdf56b52f698a9f6e2c685585028067efcc543c390f5e2c0a478edc8bd3cb3123bf1b57593c38c42f595abeff8f9753521acb875094d4f38d59a7552fcd69339dc6ce70f0707e5affd6347d39d8a6b3ac059173616df73822de993d4c9d5edb2dc734ad387850;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28e01e372a992fb54ced4354b5e87da2ae3386e9fe1cb8cef4aae2c490ecbe3878ba3e7f2778376ca692171f01fd4aac941dbd9dfb383afe2112f171c306f56b798f52569bbbd8c8e88d8428abe93a10cb88fa76cbf478da0fb452f242a684932ccd6c9c1e060e96c6e18b1e87a15ba4993df24d8b7c378f311388115630c65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fc4249e2dc57482f7fd69abc5dadae76bef79e7ca34b1494b2c51e51a64478f9cef310628235a6b0c3757e8868a3faa6d61ee951e6212f0efc41f15e9847b1670ab97b79bfc41d6f3c949c452a091d9b2d83d418788876276ca1f2e985c62677bba63b9bb6e7b3ca2c3b97fbd226c98ddf87c20ef0d613421bbf800d8aaf25a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had0749eeebf714c4e50f5337e414b526c5e3e13788af5d706f30f8037196c5df1d68bd6346e7eef55b6e5193b17175b14d5395c6ca37bd222523448afae30becbc4c6cdd1ffd4937f88f33bff40982f193c77d0e2741d8656b49738d7916b6a9c47765bc977a7206a8412e3c590b4e2b7f8bb8ab5373b7375b2e96d616f76825;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc8702090a5a804f126fd087bc1cb149ccbe3e17e022b44e95ea5f21515c60f8fc7309c61e0e9b4c29577dda8d8f50f4f532490d6e5fcdb2f6fbaf1865e6956ab91168802983c7edc9e33d2c762ce00a2ce2cea2941f3d6dc94ec605d852a0f25ca49f7855cb51c25333970c0b6a34372a7f1b43dc7d1c5f2b3731c4fba27f48;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6099f2d5f83f1ed4cc3722d68734fcbf2cb8e787ed7a5d8a822044e71f2590f8577328d4f7928dfaba0bfe25803c4f05fc2d3eb9723ffeb2696b101d1f39662d076ce214faea8835ac2537cebfff8309011ea3f29eb65432aa5a8c05c23c73a728528fa12633b8de9642a532728a2a69dab04950db5f31e906f9877a189812c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7adfd664dfc6a405294370ab0b5b8f57f378a54d317828dbc3bef52503a0b92f65d48789387ef0c6a4bc43607ed19ead294fb1728d0624860655b879fce8912a54c91287e52334fb1e88ed7fa9feeb356eef69d27398a6968ac5bfda9fe84ae8d5576b68a59e4f278cf96f51014f5fc2ee9068588a5d3795ec9ec87417d4b300;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4964bcee88ab28698e66118e50957a28fc63c0dc60d53c1a6e49035bcf7c1c8b0846af1da35900f1276cf23f0b8b3610d8cce122ae72d8e39f81c6306b779aa30860d34ce03f4fbed7230569d0965588ec5b934810c3520ea571accd255065b6d37ebb80155f29bf7f82d97ea7e561ef4d29f975c83bc82a8939af7f12c125fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7b4edd264a0c07f6522ab3914724cfb4632dee6e85a95ec439811d358c800fad2a5cd39ab8e168394a36fb4253089fe432fa23f6015cb6888acc60b23c67f3edbe0fc9ef030c18131e6bd9959fd0c3b57af002fa39a252a6d1b1f6bafdc7e85386a90f463a04441270bc9289e9366f568303b908c8598c33f2fa255aeab32a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4af0eb727c3d6716318695d64c3c1741dc70ea65b48d0e585f5f56f79b3d9928e8212be2bd86c01840913deaa09005e0bf8caccaa652aa0572329b59b722463065ddc9600443a91f7d9f6644afd759d24ae3e26431b3a6e9eccd79ebe960a8edb54ccc82fa03eb9b8b2c58b2765eb2aeeabcd24900b8346a7d4d200aab24761c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2aa94b71023f956505d49572e73e0aa35b32ab16df489561dea87879b919b129fb7312df136ce8004bc9e3788d3a7ab254c965f5d34fe6c8e5dcf9d106c76d0f34ffe695703b88d10f50f9871b5448773bd4a1b13707c63e7f92fec8a12ef7d39963c0b325a7495c06b44da8e98bbcb17e4f066df6fbc26233777d235d612d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f59ef755e31afc06ebc2c99e68bae9968b33bdfda3fa83e5f718bfc1640663e22e367bfb21f1582d92170eeef4a00d9dc2cc3f75a3e6e884e22f4be66f10482321279351f667f8420c483bc8883611e2a8ab3763393de3b8aa4686e32e5d957d67cf140312d0409a2484a4a8191aca28670b1fd0b77d153adc593c96d2c5c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1815a16de9379e11046c63cb37466bb85aae719e3a5926a3b85451f4d8a1eb78588e33efe7642040f466e9ed23ea9cde7713bb66de80bff6ce2c66370d1dc2a3683d85dbd1754777c92756e48cea147268ddf09bbf9400af3c04cc6ecb43c72966497f04c205cdb3d8512f684f953220be44d814dfd1b06c7473a516aa6b3fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h207679b9e566b515d2437e83156059c7d2a7433786e845c745a076704c5d990f7cdcdb919f69966fba8412244554146b7db17bb616f36a2cf17d4a85ec98ac220ce4096b461df6243e26cd55627b3822095ddda53a8ec9d8d66149b95d96d32a60236807d4cceec4f06befe29560d5f2fe455c2fa2d01df87df2a504e8891025;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b81dd61748ad23a7f9c07ce2ca4315f814582364ca23669cc2a26ad4b0e3e70dbe745c3647ace8a5aaea52720362329ba7a24fbb83111d9e781740df6b76bfe58d0272bff5d204ebdc632119c7c99dc7f97c1ca11e5dec25ec9ef7e8ee55299b2c0405b1f8a351b24e6a350980f5bf91b00a66fd287e5fb8885c1d4a2a39022;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f3e1ea07ec87fa91adc0ed072287ce3ced82b3c02d993fd8eda0385da0bb36558abe8105e654edf0f23a312049cbc8c73aaae3ff5f66116790427b46c586b3f0539798bb17b9e21f1260622e70f51eb1708971ff940d130990dce2800680e80c5a996a1c8523a780c850115e10298cfb4826817c64b167d3ddd25e87897123c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba3903bdd4dccc45e196d02e8d80ad8004ab4f36d1be1c52205f58fdec29a9a94f0b3514ee5e66768406222baed58febc11fc597cc56c6d8357a6078a6730c40d4a30cbcf18e0c6c1a226571945b085625baa0adf0c4aea43f643e13b9369e415d49bebf95aae77b034aee4c17fad0d32c0c14509be6d44a4fb43a5e8d5a063e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18c7ca0346f2be09fa51567c80e123d5c066d2f9d4f8fdba02b5bbb2e86104b6ecc3db0e1fed69029b32874a3829803580acbf30b5a5b603e3ef7152ce76134621a97d6713f08725be7d2da10e2d3e797593ff2300e7f620c5007a7f41daa3629e510f91d179a4d47c630d1f31d22ac3f5f0872b17dad6f2fab4c7cff45309f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd58d84511a0afe0389ef31e45a56f095bef7cc6fb42b7ae1089b6f5e467035160c4bab689df57000cfe0aff3405a8f89e2f99ffd0b56820003a2c1b96936d534c4e86672d0e1b41901ebfd7325eab93f7ac4a8dc5f1b5c2d62b158563119a5a5f0a156d0ce7c16730372c55f71af60a6427b72466584036fa3305c826870f31b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf158dc8675b9ce88000b4487d4379b6eee277d065e211a4f5e70be78330110b5adc53d142ea3c46add8e415182567392275296d05e84cf131d01a8314ffc8f3d96d24396bbc9ee92347511e39963daae1b8833c7024067d0e1f67a71a3efc1c097e5e299811aa380bd45effdbf9b4aaeeb831afc4bec9c3c89aead5af78ea6ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedf66cbf6df4818100523c30b0e5624e860587aefb9e07889ce8bb61dd0cab779067cf50429e65501e5d63d9c937b16f83646ef956a0555bd6037361ae6cb320750f7f3aa6f1dab40cd81096a8cd438c63652d7904cd247ca6778405e8b13424fe776ce4c2f94a95edcfd052da08b587ede70cb83121587d689e43751de9d35d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffc1e60ee8bf4e7a2b0ac01bdea9205b163384463e22f016ac2a60aecbe2b65feef1aee1675f52df61dbb41e92b579e5b34d3cf34806825cb0174215d52fe8985cd42f53a9f450ce47b661db541447790229ccef7bd9eb87a70c8f390078920c16f1f72ff22c89aaf4af5810df821390f74da39a30be34ce8f329474bd4dad7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h398f226f43c74e6a1b5c29d4279f65dd02096e97f5c878c154e7c060602220fdbd5e0041f8778306c706eef9097dd8372534410eb211e8dab52059cc9f1146107a3b59260e9bfe6b1c5d4222db5fdac287cd7419157a90939cacbf33235ccc27f3cbe9dd01f4e953e0298a37ae7d71a62f389d97ed52b3fa0f5c2bfac20b11e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6f35e871abe4268011b3da2bd4d0929ef486cd7e6c5ac719aa7683ee6bfd226b83f72a1a1f569aa6ec04245ceea4d98b016bd13ba3e4e4d5936073ae8f93a76c8103727ba800fd83a8b5779fbbb712f9d3eaedeee8efb9e9f0f1acd0962fc93ac5f0d5524af277d1cf4b26c9dae1beb3a7a88a36e0fc94265f22f93d3ed4bfd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd039eceb60159c65202395356a0b414fa8b596e7417b04f6be38b9fa4faf44f35dcaec2cff1ab620ac04c4c6644bd2f1d85938508f4fac16763174169ba86143b3d2b4d3840a405f567bd2fcbe43d8439feea656d5e4af5a021993c5c13b23eb04b67e4b053dd302f6b04997e402ad103d33cd774365ac248fbe999e60f0d59b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6b44a0e4da4aca8405f24f0b86dc17276f2117493d492383e50674fcb63a645bfbe5a6e602529ee987d16ec8f8d55c7e8ab605ce8a02800f8ec2a530ca60c62cb0c87f365d50a48e9372c7e84c90c4345ec175572c8f7c1bed18baba60e918fee6b2c646349a57e4e7975ce943cb1d76f95ee9f3cd16ee529daed52d5c60c85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51018390d8dd8e95f9debd50ddd468957c24a9165ee72e391e64a76097684d5726b8f541dbbcb6bffe3ec026ed48e4c8035705d4d6cdcbc9dd445c182d24ef46250d257aa720532ee86556070552a22914f01bf5221f88a0c21239377f3d3949ba0a5093ac1169cefb88f0a2c0f2b8c48e752201e143ca3e901c42696019f83c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e76ed5dd805c996689425de7b757b72120dc1141b37fd613b01ed4bdd1389337b536f3d944eaad53d41780d1dcdf08b00ad8bfe5683f4437473bc1564fd6043164418472b68650a6794fa38a24c5d76f8f28caf98944a8ddada09db1de57c535c5a924a881e905970f451f640f1da9e23a2bf040e0d9c1c267ef819477e48fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52a6559fb809650be4eea3e570b5b713fd94b37bb1cb41d8daa3a81a623b795df09ffa62f9e983e41ebc875faaac6ed6d8e1081317cd71fa237f9fa23f99c0797b7e18c899a85794171ec6ad1aaa28153397398f9a45142cdf7e7aff643e49ef956683bab667cfaba6b6dc1175d905d8d758cb753b9233919ea6a13ac70e5d80;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a9add2d3775db51b8f699be245f08a1be713bb6dfcc95d1ac98d67ddf42a14eb26d388ff97a823d0965b0e503c3196d378da69efa1d1015453b119428f7d4196f30f9e4e4836b8f72676860e8c92145bba8fa01b7a90f02c229ac7ca8b20e1fb99ae64684d8ff14fe5227fcf8ad2dc170bcac6ff001e8bf64ac9f1d358b96f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h744830c4e5a72ce9a4f1e2888fafb10cc3c011346eba15a0f0137a1d2e475e6d523cf904e848d3aab381e09aa3fea3891413e015d29085f125339f604b59a360e5ab2264b12df52489f63f0889102cf6fcc1ce3e6bfd7e2bcda74017f5f4686df44407bedf6927d98be05e88843c639e6de3eb4dc9b3674381a60a982045693d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d155743c29ced858713bb042905f86246d6a31db607972cae28b773539c9eb961e77f6977dbe4308db5385d4b841fec70a0dfb36ed503120e5a4352bf27907220a78d7ebb8f8fd9dfcd3d02f5c6efa52d62f856002342a18846a77a83ad43bce1b02c64073bdb8f102fce299d6b11648207cb2448dd4543b857aa88e8ac122d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b9f982815f52cf829013913175ce89c510565ad5615ecafa683abf68013a59144150e89f39a8500e8f84178725585268a4ffbafa6a0df72061e490b2c5dca49e621dd2c65190e0361b942e84925a2b1f46741bf28aeea2566559ce4d91cac680459aa661942698d6bd29610b1857cb052f4fca3d7c90cf0837e27c902ddcca7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb32c80c48c29de05a1e8b75547105fb4b3419514c7604cd9359d18ec56d97bd462729efcadcb3200ee4f582442635275540d531c4620c2ef27cf4d9a084feeba7d55a0c97860c725af1de516ffcdf174091afef379ca36325f44acf2335e11a3862e2715aa02c68771ce1dc0e61843cde39673922b59e9e3b9e41706d00a73fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fa7abed38089007182ea455779dce7a88fdd8b4e3091ee153c738b7b9d2e66754657e1f72c0a85e452820918815173489c0482cb958e78cfbd683354b51ae3329f5e26776f87943dce201269ebad375d964924f0d69968944da2127e1e81421fc4f1bdc7488e1e1157c7c6fe79703504f347f8af3667b3870ae4eb3d2514845;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2c9ff78d3ae1b97afaf092af37d859589b9eb46a853e345a939b9cbef5ba92bfbd7bbec278e014231da7dd7e1d433ddbd9bc40c1a4f29e873c70ab7343db2f061bee92821b168fc895bde0826e997c8df6d702e494ed9c7d074215a8249c50cba5b1ca05cc9c3b1f38248a896543565196d429f612897689bdad79616f498e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h410218a3c5bdd9a2b41e55a406c645fe237b093fa8304fbee666680b6593eae67188bacb39a8d1096b4af19af9b765df1804978b31ec7db52ec6d9f3615913e40200bbf61da9a249d7a02c37537cf964fefe594d33f60efd6925e52bf2076419d7d797d3fb549c43c5726688f704c5166881fb1ddef62c89e09d39ce5e142a30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h473ffb12c75681cbf2026f3f7b5194685785d8c2327480644b361ebc7ec376c8cb243716ab0c69c5a90519d3c7bab0bc2c506ea9882d37f94f1e435257f7f58c6368009421fd5c5c91802284554c437f00ec4908688b949d8464ee880e3594508139f0a172daa26aaf7d36e739fd61fb620a5167f293900ca8a255724f8d9f87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2953c71333eef4906ed06d49f65d2a7260c8eddd9d3a0a52655ec0d9b6c1aa4082bdeff095cb1bb6f9bb3c3ba9e19ef42c541f6e988089ada6376f1b7abcaae9ec29a00e575705127e1dd356e24b90da23a1aa9d7319034dffc4528297f70ecd867742140f2f50b266a805361558c5e555726653997ffe3a71b65ed0439479d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b6560abc370b5ca6b776ac2e96b52f7916c9a23fc04c17c8ecefb7ee8b674f537f746481038d83e3125bf3a9fda44908a067faf2d5c0c0192ad6cc7ddff0435036a93f822101280a464a8a6df623395aa115bf9fab7d300346ff22b39a84a5e834542835e882bc58edd0358e806fdf51666f85e2596ba185245f2cda84c91cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd684002b9471d15075659c4e08df1dfcb7856636ca66d558a426de6306b16ebf913ddff74795620dc1f2455540244fa7dc7c3cbfca73815b880159c9dfa59cb61503956a164ebdfd3978fb542b629383a3c04b0ba5de4a36dd003534d76359fc778251a4f61441bd3a081c79fd720473b89c470a7ae402b167ef7d18035d95b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdca63f76031a2090239b37073ac4931c7a73030186b0a8ea07a75e3c4933d3de50e535820d7f04fb37f3c21c029557acd4b22ff9b2b0c974f9309e36ec1556bde99613e856600dfd00b14f6c0d7327dd2e2e0ed435a49ed339367aaba06e3a0aee0e2302bd562a1c46f96f3ce7a7e797d88ae6cce16a7e06b2c287a95676a96b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h256adb55863c67ef694c932b397fbf48fcb3c313edc300d067626074fcb3c8605c321b8996a5bdd669c9e7bdd91ee429eecc76a4452d5e855d5adca7a126ec8e38d42ee9697aea7d855c235c53dc3bde9cb1c0904a19604846b1ebb4e20797bb3ba2c83d4f3370584fa2eb602fda698315d598cb87f31de77a7760444cb98396;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0d5865c5a840fa6d8c8adb69dceab609df13ce68d327bbea0b6fcccf91a5750729f857e695bf1047ce9d74506b7c3eac3f73223a131104af7201e8d9c22ea859653bb89b102b961937405a3a60f9111f80b1525bd222e144ab65b5fc18bc136a1d0d55d64ee13c23e14d2368c59e32333e48913289c050ac5f9ed1dde4b21b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82456db8c85d6a2fb9369fe93e0c03e549dbc4d711a2183ea69d43af9c3684e71c22d1c1b540bfbfd819a3a0d338c15cf0a5c4218a3c9dd142399d50e9615b214b0767a40e071053e7dfe739b4e1c88f34b6336beef88d43249f3303e1a21f6576a1b0b2d5d0a2b8dab6fc6916ec63495a88422cfbf8432ab42f2a7f5775cf7b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d5c1a33707ac0904995add72e28e82d0dbefff175ab04cb1deb626ccc895869fc470775cd24ff6e890df048685240907e72a9a535e7ac4b84f7c7bf6ddbc40404d31b1c5e3a13f7b09ea0b5745c5d2fd9883c31d72ef86217cf11f0c39583a7a4f15caa1cfa3b9318e30e47bc6f6afbdb05ba81ca89e0c9e415ca010034c847;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd35b60ffe62be6d32a8bd75eea425ab307bc5fe3aaa7de8a0989d4be1ae7a1c8248f348ef3b28e812a93689c920203366f70efef0604e25723b7b3f9de26de2971dbdfab27b7c3eca68d35a61dbd8968d66adb384c08e4c07808610dd5b4fba73ca7157880ddf8929d47540669e21b6533d995d9e727007289da46a88123883e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb19d2d40d962b67a49c5f01b3fe8cd172c85f5a53354216994599604fb72af9a03be633380f418cdda7da9f740f2cc1cbc05bb6ed9e9ef00d2c0a37c815cba0cc26ec1c809874b82d448d3f6691699a78ca69e718db5c618b13c617e128e5326a8cc575e5912a5a07018b7826bf74f680a7b274cee7460a5cb8a0b658e61d2a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd733630155bfd1a6eca3c9aca9d4c1b0988fc26e5e05f59c67b9dd2284c23590fbb967292cadd7153c1dbc25b97a0ae8eff18863cde712f4934e193c858e383d49e77ac4b5f06622a5bc0db31aad96cd92791e31d2f117f74f8956913a5b3fc344b545d6ec0a9423dda49d323b9185fd302c988b1d0601d7697d7d3783ce2aa1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h927273f19edb40d03dde04d41bc739b0f8e19c5274d8c496ceacf355bdefd3efd8565aba74e0654d229e5f15a789ceea9a73b062ca20f1c434e323cca978b9699e7024184fb5704889f9322d915baa28721461aece1c1ef6b0c9a4beabeec707dad61dd58c17d80d1449a14863899e9d01b1bb2902c620db1b94997e1b330eb9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb81eda2a028439c308d218a71d4f2230f06d5e1582a4094fa9ffa390268c55c178b91c856833632536a13b0cae6fe9f637e59925f002adc7b7325b7004df5ac23a1714e3d905588bb7458ef6225bf54adf0b8fc133b852703078b9534b0e813dbfd181dafb895234ad2dc4631948298a939a462b910feaee33fe50f03c2b807c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59b3094acf384bf297352fa986848f3a3d96633c703d4cf99d3c8ef519e576fc28a89907fb2ac55e8856e6c5d46f81572b3acbfceb23148e0404fe5ad2cdcc50b75b4811f90ec807550bed08452f1d10ced207e8e10cd589c13e0d83b9981fb801806b9e224e601f9831fe38959bba660a6d7673aad3267d03a7bc2a47d99a9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h543ee25edb841b731900e535d6f8527ca42663380970d1d28c7f2991fff5a6ec80282cd993f01b4410a2fef57a48837f0d809f386696c9afb544d7c34b8af7a321f7841b7da6e66626f94aecd3acb44bfdb787b693f3c0aed53e2c1dbe3c83cfdc429fb5b280065a12441fceb553978ec65afd6478c027411608d6957a3f8659;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fe1b5c3d9d6580992a3d210214c54793e0c7081aa8d5e44b52864b34b4ac82d2db72353153ea78bfb6701263103ff3e954e13a67fde027d84d4a3d9925061a6e1143df99d3fa0945126a3a683fe126a2e472df7b17c4398f6c611909f2199e8a7eba59781b00f510a0c5609fd4d8d1b5627c1e34b8414b0c87f2de386ce9170;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ff02247c53f758611d9c852875b37026b37eea27c0fd868f963a82041468cec4a49fdd1ea781b35305967ba9b4fea6010889b1dd0799393cb3849b8fc0cf86afd5762730e245fd2589849cf3a8c2df57814fe6d8f33c11dc330076710918b63618641e1ebae307dfba5cbc7d3396f0b5174fa83945a8573a0dfeb0d7f30022b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d4caefe93d44e035fc694b74f63a2fe6271fd91b9bb4ec8db6f90eb47152662c59c91ff2c1407d9d0938ed414aba67ec676a2cf0506954567d73663f5d24fc1a6f8a6fce21015df7265e1bafd240265fe74f376fdc94a391336dcb444b6fdc8730441f4f2206c54cac0d80e33f58ab83a9c862dc80974a45236e85307f65c06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96b4897a72134c8ee9b20f09c0d66c738ef0bbd3700809d2455563e9e9243d6c7f15f279bc20734ebff50d2a072a8cd4a29e3d9f11fc228d3f2c8127f4f35323fb4385b11ca8b507e14ef7c1d3096b01805cb7dab43fcb39dba9b25a04f2a4ef64d5d91856c2f4f991a8963904cd2df99e58c7e5fed762d4ec9bbaeec7c84b2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heac8be5b907b51ae3eb110e1e5f92107bbc1d7b272fb36fd23af02c5844bb121a9c7ebffff9e82541b213d056283c6ef8cef7d1a06f9e91d6574553d35bcf897dad438b28c7cff09d805bef6903606b204d6de68b99d6d53431596a56a15e528bd662b41c388374926083e4e9de50aab8219f88eb4b1e1acdd0cf02557acb43f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e5cbfdc44227345759a7fbdd472918f5fab1144b3ec147ffd9ecc24f5df4efc1cf91412e37ea239670320438bef481efd8f6124eed45cf3bde12fa2f19d48c4e567db0b4397ba8354d0f8856f964882a7cd61bb21a344bd37300df3f54eea72d82c49c7618d007e0eb2cafe4cc29690bd7c63e777055f61c23a0b9b8f5cc4eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f8095f1df868ac26a569cedb19922d7f57536efc84bc99c9e41ad5f301457526e899b61ca9a3f73a65b1291b496f97aaca00225a08ff02ba96df7b08f3d58ed5591795847c69cd6897ccede8b0aa0cd89a7ecd14bf0b84256be50df64197a8ddc03072a267276183e3bfc11677b140db68fae010e8bd095dffbb79d25f0399c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6563db6a16cd4efe9d2023324bc3002509d1b165c136b657ca9c190732e92eed52ee1079b80056368856e90bd88b29e21503e3f3716c9e7778ac71c08fe65773dee645e720113ca80a8509164aa982b832a4d891aea9ebee1038d05344d7f0bf6bb688c2b26f662be21c575ee468561d788b2991519ecc756b0ae7c3993af927;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30945a0e37030e4d105d5738694c9f49916e9b679ed1dca37fa7fdd48672f3f626e5de9b95d203cb9658e14437fe259e8c08ff0b74d6d3cfb8a7d346fb7352e2ccd8f8d903dcba0adae159f2ae97a845d02061f7e955451cc4adf8805a55c637260773032cbf513ced52fef873081d5cc0520f501d455e75ca3f31c21b25ef39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb81a8006665eaf6d94cc2d3248b495e16da1d94fc39b0a1fa147b003908d8183a780272522b11ac48b18350126c6b8f04eb7281732cab6ed3903940e5a355ea66265dfb86deec3b62f53c29463aaf4ca897ce467478eeecdbdb9b920fd39a607d683713ef5cf0e523bf01bf03b6b43a479864c0c31e018ace2a43150ea8f530e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda62b9c879816b10741b98253275a6fb83ca4240c7850be877b7ce655abb171464b54068a3a66e05383dc2ec8c3949ee9c31e66f1d863514d4fd66bacfbaca52466a2ba045cdfa41d1e5a263267622de9f4d6f21ee351030fe0911fe5e873ead068d681fa566bfdd35e872fb8cfb3a294c4c53e6e97914f5c1760683504fe35d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h703b4693fd7d59bfd439015827dcc59f569ef03b98d5c6a47fc18d2bd45f3823b720f26bafe4cdd9dad0555232d1187d4c315b277241a39bd8bb4b8396661a5bd3d17cd57c7b3e263fdbc8d148ebdf7dd15c56f0af52e337d78a62366d43843467c5969d85abe12b3185afda7ea4aba05c5cce23d0e816f9b31c9e42539840cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38c981d9036103b55f9f626fda3f8e955716d50c5ddabc7e3a82eb34c7fc8b4674f202bee276682b832056ab2f6e662af06870e62a0ec6d674588826ee13c5a339c394e5bf5cced47a229d91b55206ec7e5ca4c17c2600eb2417b04f54febcb746988bb66cb79aff01faf2c4807f23dd964496456676436a596d6b570c837112;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccd16e0f455ca687cc0b0fb453162a6d6ce0164cc1ffdf48665588de9df89fb79b22556b6946b106435a54665ec00c156201a04cbc34ad46c1d0d360252e2094ba06f449af0e60cf0469771509f5eee0c71cab3cc87d8e8dae10f07f6e01c64f7eee262f64ea999d4eb16c5034f8efaea386f8332b5ea9159f935b53bab5afbd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15556a805d5b3301ece1681dccab4c7cdd651b4c23f90f67aace7ecda20410e96bb834b2a69fa84be44825fba3f7ac70af6d46f90ba647af48761a4fa344408da4adf689cd1d2378a43256479ff4ecfc6e02873ada11c46731ca8fb34fe88ad740275b702382bd2921798805120ad325a6ebe0473a6672133ab2a37f56f2830e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h889230d1e048567e7585ddb7d0f303846ce95cb5a8f060dd3c36a13bee17ad580a289c77253f9800c884971320a22c260b03592f3bbf30cfd8209d6f050599b716bd6e5964d86100b2fbaf233047fd08832c063a6e3cfb863251d3b4134c22bd226b4e795340c3bfed054c811a26dad40cdfc71f1264b8bc58722a9be28b2003;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9cb9df09365ccedcb6242bdf196c9cbd6bbb2f24060c2ba266c783a0b746a06a340c7ce15eca4df16304842eeb04157d48c61f259d5a0ee5e9ed523768eee3e58cdb1f72951eeb819a7dd83bd1c87fd5d7536d8830d5bf2afec457a825f83c8267678b05a0c4d30bbbcc42e1b2e5954a9872051c59e08f1fa647a800a3a02a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedd7e8ff28b7ce756ced4a22d6ca119f4950e0c87a4c4e2283219eeb16a19791b2cdf53f3ea4a63638a24854301a59591a24098b0d9963a58eb169404ae08cd7b67210710d23850e3757c64dd53d2ad51b91209293f4ffdfe577887a700864cbd0099df938626b6d474938be703f726ec40c2efa57a65e23814d3fe7a0f74e1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6af05ed38bee42aede2c6154a5c952581fee5d3f8e4e1ddfdff55415ad77c59b73fe0e9ef4d6735db8c4669b4642b491f4da534027c6b94a388ce0558fd8328a1f30783b835f8f693ae960161db9b89c6ec2c9cbefa04f88a57dcb5e00787688eb5e4a9f9559ce8bcf4e3b83cc70bfd4725d244a05e21d571358bc63bd26f34e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e60b04e436e1ac49ab389c9c0399cf2598f4166c7a114102b3d47579f7811eba5b9b8b30186407577b23442ab2db648cd372ff0db5753ebc3940c03f60046edad38b9f519a6de706fcda9dd3a577c0cf5941b213ab3788c6b8078f97ccc18bb256cf3fdd774361cd86c3ffd954b2c3a0f9afd019284cd798bd6144bb5e279d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f47516dc74687444941579a1953388a54608fac3290713f5ab7b77ae715cae171fc177837ec2445f33baacf67f5f5d4e17113babc4077312cda68c06d95c4377223e0ec756ff7af45ec9c0149e0370207c8b8cdd1c442f8d589d3bafe913b32341dc7b3d92b98a2597bf095a79a606a5b4f707f019d5ce7d9b383893dab31f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe0a4d14565e96450eeecfce791473d8ef429e9d2e39817cef3f8fc3336f22636c9a311d3e5fb0cd9e1f22b70eed9b061915b1e119403037c0b719d7a3e4be424cf882df263a1b91f2565ba029cb9be5ecc2c20b4336f77363c1554e23fedeaf7c66b6b0611d8bd022a8464c866f7f94d0a865e2f62ca883f173f4ef04f77a94;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbb2e6eefa32989d098680fbc7d76412bee657d629e325fe4b1f810ea53a9fce84de31d3225283f06d19fc55a77bb46083df92643daba4c3f672bda0501cf9dfe3bb6c5dcf730d88506df38c668a69d05d9eaeae2d278d86172383a74ee8cc71a3ebcfbb325f3816ad06a9e842f71469da9e71761fed0e7a4ec47ffe142fb157;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc43b14b14944f863d7be881eb7cbdfed0e2cee286cf76019771ede3fe57a59078851f77dbe76b0eb626c6e14999759c1cf8ea3d0d8818ca17158cfdeafe4d9fcc19149f714e06035f420c7238906622915965c8e92fc26e112649329614b2550e183c97041d780ba28bf1efd1c8c30fe26933c4c160df734bb9135df29a8a504;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h164a6ed6a60080e6dc9653f80d47b73cb54d3717041a65e741e7d2ab2327c7352c6a7f570a24eb57aa45d50c35994b15959da9f369a298dd54bb7de04c71b58f054b5143a8c3879c7ce94c1423fb342f6e9edbb7bb5d4f596071aa86af49de20b9bd531fd9623011112fc40142f314003558c721ba7d99039957845784141ebb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ab01e85bf3265ede1d0d8d91243f7fedbc31a06fe39fe97cc1031f80537dac022d77f003e5dc3232dfa36ce757c6da07fc71f4d45f389e0d340a3dd66e2ab202666628ed5051207e1417a5488b622d7eab1da29cbf5d273c219252aa323a6ffebdb1130e3c9fec235aabb10ba40b0ada85d2386650b5c807dd1bfb959060b15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7946e34007b88e81da62fd5bd36b030a7a0a20ca8936cd1576d59eebcb7535d767ef3d737a5b6b94aecc21bf99955596ee3edf96cb8f92a1d7fb9aed06064ce5723ca6073b39359bc1fe5c052b9a781493e9ea1bc00f3a188be893ce768cfeb22d130752b1340c234bf2540c3f122c0d6a2316f5fb640eb8579e111d483986fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h915cdb2a7b1e469b5a0bb6ea41a21de89659ae00f4cf77d3023dbc0ccc61973ff5eac92cd07f64b854ef76e1738d037f7dd12e0298fe4762f67565488a435b02b14244cea28c071646288f5fe655b2fc0736a4a7a361841728abf91582f64ad5a46490babb354f55e799d2140a63597730dccd445550b2471932e9dc27ef59ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1bcebf843a11e5c75e774745a1300147fa92031e894619fb5b83059cf4889e25037a6285ca4e922ab786cc778c917575ca83290d24127d1bdb3df72392f5f49daf3e060f27ba908183df14962a060f7c2a9ed30c6828bd9cfa42a394f82843d3ecae11e563d1511321461c015d12ac4cc8eed3e0c7bd834fca115bb13b8e9b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he14cae7d4440974bc5d5038638fae940528c9a4f6a23ff6f04cac6e93088f2d8a4f5dc598d6dd0c69a8a6910a621e0994cd42d2ad336fd48b260b2550402dfd2c3bc0e09872bd3738f08f48da4c614f87dfa57393d5dbd7024b9a4728fa74899864cfd08f2357c33e1188eabc70f05ff5b7f0509fb64607be0bb0290862eaa95;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc47084bfa2320b23d8c4d4248b02e36b3e091aa491f2cf3aec8abc0bd1cd52aecf17080b9395620cd63a80eb9787afa08235e13c43339369b39bfbd73aa3a3be18435f4ee136fdcc121e4e559b1501cd0a5ed62340624216a01cf391092a60768f3f03a3f5304b29fe94778d54eedd0c4e9e44640f6be7a4723717fc2d73696;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h844edeb8e2af4224176cd4d82fe00cc2396415ca69f9c432126899d3694098eedcd716ff25e3d5e74eef3fb3d8cbb1231c5ba4217fdbfe8ba0914128c0daba7f4e21411a1587f56163bc386f11da8bc9355a82b8a9dd34ae030ae1a34ff132308621f00d50e988d1f0b43e3986c4ab51ccc78cc9b5bd9adbab71389b630b0819;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5a736c3e41fc13a9b0204b512b2839fd458859d37ec30458e57ab8c8e5d3a077fe1d52f0abd1bb82d706b7168d9477f8f13dfeade0894a83f54c2a4fdc76a2e78d4bb7d61f206d29d3b35759eb1a562d94fe238c73613327b1951b4046df36d02290cc4e036d12926c6e8aab5562f559ca8cd0e90274fa4346eb07c7a80966e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78edae1b4b50ab17716b092bd78db5b4a810f01e4520c23db3c8e695bca660e97227a11d96ac060c2312fdd7fbd411b3e781a3f45557a168332cd18e1287b756d9f2c12c12686810109c36a023f890d357c6b57fe2a2966e2351e66e02de3f727804136e0bdad4f64daf67a0f7bba523300d341a47ccef3bffccf1e031cb1db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fef060d928a8621af5f63b3428cb0ea3a6f53e587bad16fac5272ffaa5cfc0d3dd7c8a47d6cbd0e6f688171c13c8309a6295c370228bcb35bba6105c28c486dc26787e9e5af6add051c397ae33ee6bf5f4e4325b763ba7eac4ee1c180e826877a6c7922905d0fe028d1ccbceb506345ce3ddc2687fb3d15cd7e1a86d963c276;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb02121d69d470f00af7336d080f27426da0b65ada76c4f0e4a9463ad197fb156754c5abbbe0a346d5c0fb2e2bdd21b51dca06e957267e9f34bade0aa24bd02af69f0c2c1ae381cf54a7c9fac62495af6e1b302f1097b5846aebd4c2bc959b68cde9b2d6d6583bc2ac5b31559e8867a97c289aa3636dc7839140fcb536b333e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5087d32cd8d54633be870dc565ffa868c89fd5a101f5096d657c8f7006ac27370723cf114cf93aaa4e044f4bfb2b64e49d50a936fe51540b4cfc8c218327c5ba5a0dcd1604e56337373cd1617ed4e557060817c82df69a1cd8b2d9219542cb9265564d69c3b730ba9765c3db5992a16c9dcef8fafb4ee58dcb193ebcf911d39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbc7cdd99ee414e834241074988e2c8a6b30ea27de999875fa31dab714cbd005a8ee09f7f31d9dc3a9f89aa231cba327ad96cf674ad2aef2aabc1795916867ea5d7fcfbc9ed1a78ac12b6d67bc692a98c50c0331ee64aa0c0f324ebac10e07872607ac758ed865d780ecdc76d48ed94552ed42285d1206e277e89ccf9ad8c830;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc17fc511ba4812859d63f993fe24cc131590f638867b756c5e141374c70efb6a2eb87cf157cc117b5f3929b83ef2d6809a1348bed48a97d4d5adff33406bde614cee91a57501b6b71c26b22d25445b125293586b206867873386fa8f2d9a7ff03afdda26b54e3d3feda535c2c46045d4a238ffe0088b05c15506107af0a93d85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38f31911b41b391e93f6df66056ce1f5e27d20689a6b2f9212b59f5d2c188de4d12f7ce13049cc31721c42b5a72b62d700ce845b7fa5ca616db50d4a1b55007bf99b254e7da9c40c7ee197a8de607f657bb91330339cee3022fd4d4f24b0c516cbb52581327c4dbff8516c9458b7acb3a80eb0aca938e6d0279b6ce5f2d7ecd3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed3d9da3aebc8213fd3e9fcd4e7a43893950cdfa70d10cd9e4f117ea174011b77cd4bf3b47dfee5557790ad8dc60b68cb9a6787f56f3eae20a4b24075f840e8b8877d57d5c72e96e23f4b32a13f52543560dc6c92a4fb1af33011224622c1d81bfc1723e4308a9070567494ed48e233e76251a471bdb0a65cafb06e89a93b6ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1df50075aefab63dac8abb00e7c53d7942a110f9ba4436cc175f139ca0ff7ee07a6fb2b66a9042389ae4fa09d6eb61a94261b52c74de029b2a6045e3f5ea3d0bd49419d129ae5340a568fd678115a9ce10d766374442303e0a2861348ada891d2349a9ae47a2152592efda1b928b5161f8d56942eb291fe157069d02efb8b59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf9ba9dd6e6dfe7fcb73deb85e35fafebc82ed7bfc736ac533bdda652207614f2944b004fab49479d58dda3f36fbabc8e423ae3295eaca7da3c480836223667ceac3e8d148c23d388369ca4d002b6e5c1105de5fe47a6ae94c5f433a8b6e7a871a7aa16fffa0cb59bc3404da2b5b9fa61bfc7be41378c20752f21e1db787f114;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b07e4a953eacc80d974fbb50fa05615f840d62bc6ef775df610f0beaa9a97d3693daf656d0c06e5373b5b54347efc767abd09ae22bf793b1ac3af8ad2fc68af986746e407e472330a2e69e8cf087da83920c2e82f7098c1f9635d5ff92e94c94cb0f2dbaeee7dfa3d7bb7207ad649bd2f07546f9eb6b62d7a29cbd24019f2a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde393ac571d6906effab0740c9b3b3d52ea28376fd31c771220a1532579bf0dc09b032fd7f9c770a4e2a4969102a5fa0a334ea22ec5ca0dfe68f6330199f8fd04387b1691fd18af6846664b97fa90b67a07f8d8ef5d7d215ac65a190044386df6047dca011271d2603779a99dbeae8a74654e68ead495aacc00fbb5014187b93;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e1dac5ffa34902e703938e0398f3564a0bc5444305d04bb4cacba94c0c55ee09101e085c75474ef52148cb908e5653b52b9ed1b45602a26424bf1fafe844c26d2f50562773ebd2680234176203e6fac62f88385b62a1c542ae4f9446f1c6ee686b24bdd6019bb25a304f75715d25147b000d956427afc7633d4bc9804ba34c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72f278633e3008a46c8b805bddb195812fea4af941ec35c15097014971b72e3dab0c7bda85eda0aa47ffac48dd1e4b6a92abf2306dd77de82d597656bf42263bf71833d58e1ae411b79171e00b1212aeec33eed0f70ca58cbd07c65d321e961298a34d3a56411583882acbc91a057d6d60b43b88f262fee6ccc9fb4531aa264c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c79a504443807f54f61a61ec9a58edb5238489c6140e86c82c8b6d967aea91751c79d365b3f3cfbe979fcba61b4fb9a370d90d9cbdc624e2a02660058ace87f07b51c7bf483bb24f25db8c4589da47df5fd3d52ff784c5c3077ea8aa3624eb2379e261a9988245a348449e3dd0403ca82c028061babbbb6adcef063def6d64a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ed7386c871c2abecd87cf9013fa900a1268be458bb0c31f8aae69ffeec16254de62dff359acb836f8e1281cbd134d253f7e5fa86933e32399cb11ff47e73df0a80f9a6d9ed6f3de6008c5c5670fddacf3ea69c3fb4bab06567897e8c7e5c73583bd80c7597f21fc28bc2ed42bea329efc4681131a4b048db8b52e469fc94355;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h403bfd7cdc4b12fde8d93c4ea95b63eabeaa5eb9cf997e6e1e54365f9686a468bf856d8aa64f5bb8c63e90de126dd7b38993b9298d989bf660b9f9e7c1795c1a323313bf9165b73d27d12a8072c69c5ea5f3039e4ed59938f6d5541e4d74f9dab160815452a7e6126762abea54723dd358b4251e12f745f53eec548b96d24494;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f70ed4fbe54f38d90f3e131ead83bbb6346d95b56209ac37b8d71f76e283b3e78842fdfc3f814b701f6b8d7262af9b9918ca5431373d1a28323e66648da17749419bc57178c04dcb0dc91cde56587b2e1c8ea8b3978e5a9f59a7f5a42bd6f52dfca932489dfff53bdb7ed6293d442dd983b88766e8b70a228108b149ba48d2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa63b06710b9c64afae256e5d5d53b9c0c0116e2dcf7a663c4501b60f0465e6e501d138ae7e0b8b62bfd831ef969fec04365673c36aa7f9a68f6cdfa1826372eb382d77c9efd493a1897fcd82e4a4d39401d8f8a2819d2da69bb1235a3d91bc191432232dcba1f7e2825b7a24f7c2c59e53fdbe0e70162caf6c5853a4b2f8dbc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf123a39287e42cd6fe021def87df27323661eec259ee4e9f292629fc93eacd888ff652ef3fca6436c75bf411a4a61f4d6143f5b684c9df0ddfe4f799ab40e7ae9e72ff62b10b8836c3dcb780c795f5030438471fdf8ce2abd7d70073019d0ab6d73d5d19f2316065473fe275f3f47b91acfb081aebe50fb1713418651a35fadf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87114e46b402189421c14f8967229e705debd92a0cf91126c5001f1f40cdf02f66811ed7b9b2bddd5583c9d3a222bc5277f94909e776868c34c1a03bfe54051fd683279cd1417a0e6af0d9ac3fb3ecef8f482164fbfc3b1bbf66ef6534ecfa64c0a82decf9face2c729ca93e764b4da8ad5b3c5477172551a64dc79eac286dd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5bea5d162a81030b5b418e5666532059de4767a4dc55089dbd7ac3ca8db0480db5dd573beff0c8c7169a52b118efee470fd4ad21ab32b8d277187bb7c597b4be43237a6cd4d8cbf0cf44f42a6454b2c0d15c843020b08b66d431505448a99c8d9eea04722a7f8943bb55ab6a8c711d33bba4566ef746d1f665b19bd69389b7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9101d36b2f631c0170e845adfe3812178d456d922ad881bf22872030ed1807a64734f8420937c7952640531495e30775202567f967c494f7005d905b2c6a0f5de7e4dbf87c42d272734a31a6692c99594ef85b0a7d36cabd1aa3a1bec9d72b8280c2872f394b09ac744880d31f3825636b26fa20ec5f15ec25101b8d27d16756;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62698566bf69db30ac9bdfaa034b5c8ef6d89c8f02f6b36401f25ccad53feb56875037232599d0ee319acaf218067868441997418a3efbd1a009f0a7e7823e6d927f1944b8eb2c8680bd7c6104b2907aea2aba52e77517c0abba62992dd0da2d49bb08265c5593b880f0bebfb187261ed85ecbcb16e2bdbb2236d82d170c9e98;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb90df6aa284b0c48625dbe6c9c44281c4ccaf0fc13fb121ae04b47effef008b702e2d8bb0c2386347685ef0d9b1818d4e448960ae3108a228d5d6b87001f8e5d1e87edaa436945b3703d32cc5bf6d5825afdfb4cc241ca87958670edab78c49d6681aa1e606ad428ed5bc916ba6bd2f3b975afe7052804eaec77ef96c61d0fc2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb23cb13306de3d404c5c83263f0f80a7d3ee82273ef3a2e9014fad9d296e55612453646df8964ffb1bb7b2bdedb81d8e37fc1ed2a5802dbdde5a66099fdbc23cbf0dcfc4367c45cc74a4546bf1909a3e70775397050c242d23f5c12969f34c8233c757b37d30b50898c8f710f122dfec0a0b69df4b2d1df6f8d97af98de75ab6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cfe87e42b003b972b080e722eb7d321539f53a42b040619e9fa1ad5a28bebcaf637bb8ceef7c002b2dd783badd9f9909d7ff32ed59728838c6e793f71fea6db6e05aa3dc9ffde39d53c02807cd7bca227392cdb6daeafd535fe64463cf860b441b8cb797d76e82e17b1fd760061251ae5456de14919438ad73fe810c4dd9042;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h720f963cfb4d000751b3dd7af1bf60be766064eb1b0773a9c268a63ca397019a38425a96799eb1084b811ced36775d7f9c1360e8fce533486947118c5b936f505a2e6076772fb84fe4bab473de73e0def247142851ccf4f7c6688f425f8983fdeac3075d757e7f84fb980bf3e17ab84cbf7b84e17a6878d3d49d142f3702ff2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3802aef978217ce2dab67f550242cb123447c553970dfe6eb019fd51f883fff73f512b85897f57f9dbc46ce1a5fc303ab5ecac737acfcff4caa78a0c91d4cdac39ea2b3cf010a8b9f8036f58656f29752c4f59728239bb910428e1e9df6f8cb411fa76b9788de6eed9c2b1866cdb91638ed77a65a4b256ed74ed1fd2c6618c7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde844abe261fa090653bc0fa6d7401203375ca79e5604ddc6f767586e68a6c0b6d32d701e4a1e572892e2b77e5fc4bf7d7fe18d74c19aacf91661c3fc93a528f8bbc4f25201913c34d6712c41c895fc2b5d1384c8bc7b3ba27a1451b0ea8a5519834ab6918c17d930f4a4108b70acd462a3bb2daf7b424b37591542b5d29ea8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8203e5d4291b139f367e7aab8561a732debd333058be2b2c6162db9b79daf8c5eac5129073ea18126edb8a1e9310c149e8eb2a14192c6d9331bc0848fd36eb562f7a2b900f804726aa814a11d629f9afee3d99464bdbff989a2508a8f704bcecaeaf62fe4038309b54d9065e12ce34d7becf0c540d6a1be052673428de572f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83b2164d3fd7f1da6fb586beaba1fd2811499c8ffa9dd675f9f172ba8730996d7007a95847a0e9ba93f2b241691601dbaf7f042b427226ba2de573cdaf3fed619e40c01b937e75b19c7c31e7e91dcfa0b637f3e6a51d8c1ec564af75ea60513fb4a069e63f2074a382219c944a3d159ec05209006097a344c506b5d5932a1243;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h292681981426b2096fd7035c1db998ddd507dc215a6f08824bce7468532d6d9d1fda36c401c1a8e4e4017282c69277496cedd76f193d5479f89c459b8cf4da1500c320a31e26f5285b1b36a160bae6f43ec556998805f43a151846ad6ffba5ebbe21767b29d9b6a195c9fc89a11ec0adec0695bb401f72cb40916e95ab7c9af5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9381ab5cc71e9d1ae5b5c906cd7be82d57a5a6fa04fef4391de80ccf477c7823805b46834418307f1cb28e3bb7c142d7e08b293e747ea2eca0562ac4c4f68ed5214e78d0e30755d4113f228473c1a93068a349162da95822770bbea39d097a40c37072e614a562c9fa4038a4f3e5d97ff690e4b8a27a0dc4f6fce2a9dcd54760;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5aa921e702012db1ccfe0c4abac5c08c6a3e7cbd98ddcadbbe657821a4bfd947b286a1f9ab30401405e8be2be6480ef8b6b01a36e2bd7a6f74b1513e431200d59f02f93a1466c014fab196330a9d64f5fcfe9ab28bcf2ae98538c3403b6a3e7d39f0b93b5471b87656880f77933316a1fe66e3bd68fc03c0186eb6494f0e728c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h516724b7aedb39d3cab122829175fc442a54c18efcfa02b3b40f4367dd8903d18024b474607955c5c5917fbcd9a1c37e9d0f5fd96eed2a64c8a57cf1c7a7bd5b63d6f95df0e803f3607f21f3091c66e53c39ed7f08b98e0f2be954755dc021750722132ac78fb56d2ef0e4c1e43f72fb3695faec76f305044e6618afd911a78e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24f3c6b82f76b225add5b607fad6551fc4259ba5a358dd32a22a2ad79c1f0b3b80abc92d5d23bb238b5ca6f2130506d2a3de804da2750f972ddd45ea3acf869ee6e7e6618673c610188338bd7b8ae12e5262e1ce509234714ff86171a5accbce61edeb6a1edddc0e07e5dc9dc7ba1d534cab2bcf5e1ac1c8dd4bd2c0c416cad2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9fac937c7b82946268746ae9dc57ab33f88a380c09e9f4192a7b09a00c890ba3ccfd24e92a7a70c440b6899721516644c636a38e62980d590c5630eabb2bbf28d6452933d9ba7bbc6118b1338d333b99b3652c48ee88b0fa9a0adcb8865d074dbe577cb4f6e0ba4a261cf5a721dd77af44982091581f3eb6ec3e8dc1f622fc5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bc613a1e6b1e798da5dfa22344a8e7a1cacf51507c6e49a5f1e2f22d562199199fa5b92a178a8f7db65eb52746b5d863d0ca9b1f43ee6e67861e30abeea51b5ae5bb29c099e6be1d7e086314c056845b2ed25a43aa37eba1a8d4291f0b62ef1e2522a9ff8abfa248489e45af3a3ff74999344eec6b5bb65074c48f9f67b7688;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cc708ed0e20d83ab98e2a9645001361a28d8c0a8d43b64371d9d8126a1539fe02ae60b1d669eb1afdefa51fc84a7bcef2b287fd2394d2228ca7173e2aeded22b1a3cd8a308db990741575058be193f26c82a54df66a1f34e046daa9e5a41e79b9e8a974db5a9c5a8ad64d2e21ebbad1ea4b859e492eb858d116f65dd5dc0052;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h482475514ec371ab1ba191006c0eb6fc05382c76abdd47b16f087fae1d8bb01a0cb55d0645e1ce41536a186d2d95d6a90ee49c07f94d5dff2042e08edb72533b863856ab3616536b93a9ba9c41c94d1a4e74d40b0a795bdcfe9d35a5764a17584cbc6942bb56f3b6b05cccbd4bee1e7812e0d1ecd35b40bc07b64413bef9f58a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf21066ac5fc02705cbc9464631fa2f66c5a9a0035b0a0b034894549145efbe449dbd2b78e40f3d18c1cd8811e7a7cb7ecb9d488a07985a8a998b623f5be025d96706a06bb434a89e4da05e8e2e99c1cb35d313ea7e54068170d299d5570122124a815a9d6df7b40ba23ae7456daccdfb8de84ad4db5b834cb4c34e038aee2387;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f6a329f1657263acbb86d06728b3809cf387ec61d13cd58c07f8399983fc85f7f3fb9ed0b4f10580e9b11c31f04490d10883590e9f51d5a61a0df01dc70fade67eac8a38e07a9cd76b6c1905b9e1c551a4ecd024456c4b7c5053793deb55c080db9ce10f316346b6a130edc30a1b79e94e6e1aecd91bf5fb2ab9e1d398ea7e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc13516b36dca524a258985346e71e20c1caea4922b70734729e819866d0be0ed639e4c26ebeb29b96c849d89bcdda42d850bfe393089f7180400c8f6016de7a170a570bd648ede14f1238408f43a6c7db2221a6d349d22d9846ac3d637521b51f4041e03228043769d69546de0971dec06455e8cacf53df586ee712c9eab67dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58946c266e13f7f237065b7a51233f7517b4dabda880d5848c7c8d66d6a1de052247849f02c1d1633fc494bbdc1af866a67343278bf0a1d5a692ef7751978bd5988e4fb07ed6f482cc2b46d4b55fbb5c597b76823d26801e0bd27a3c563b10e8660ec5a0b47be3d2e7e6ca3367b646a400a5eba01b3083e1449d2808e7941a9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff8275aa99c74716c2a6917d447bf40edc584263e77085518d053d2e966f5417a5af768488dd585e4fffe124521ca17f5c28d688c380cd56bc1bc2fcc89cc9bd25ad7b84a364d5af07d16a0c3326d32c00cf22021a36537cdb5ac1d1e97465c84579ddd9a4d6f6e840701f1eec9555b2abd6943f9cf0cd7676a0d92d677af240;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b2c6be8f682be196edba9d48733bbe224e47c2a47ff6b5d1eae5da9f42883a6ebfe51f1e96447b127d45b6d014a0f3eb0cf93edb0c9572bd32317a2f25e4766301197c04aeb067bc44c66655dafe3e9ac87d4a7edb4775f7c4b96ec105c1a0d394a953db7432293b14fe901f1729ca7446ed2ca116f005db408573bfece5ede;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1785817a2697da07d7edc2d3db1a754e94cd2738b24662fd4da3d6d8c348ea4fa1d275192f29afcb46c8e96168933c43a509b8f431f3269f72248569fc96b0a4c2d1d89344beaa8c1d542e486e15428d02c84937865d1ebb1ca4f7ba28297fe64e6c888934f914d935add8e560ea60c820f1ab75fe8be6d17669ce4b024642b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd205b05ad906cec0598ba003a91a8ab38e57183ccaf883dc33bcea36664baa859374de44e34e598ead4b4620819a13e4bc96a87ccce142cb1c1456ab9c5848f30e5e2565d688c813401b984c3335da75c489b15a3269d75f72cb4e14dd7348b66665ba366da35523920e056051b2c66eaba115ee8aa7e82555503c60a3f281ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4abeb6ef4b2454bf55416c31b58241a8b2040a03167ffbbe23a8c5644cc818abe28b791197ac5231fc9c2e922fd4126bb29c1a36374b2e22667cac11c0336284928477e9a5d65306b6e3610860c65e1c1da038ba66725580c3daf1f885042bcbd5de73600c9e344faf052b12079a8ded3734466bd849444f32d6ba5b5b346c04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb1fabf13765c8f087dce7be8f94842991580f8353ba0149f11e06f5e3a137e96bdd0076cbe4facda211a45be783a29d8d70e461245ec50f1a47f5900e4592acd4f188de284718cbcf6ebbef23ca080fbef1b0e1f86a1040a318f0e600a6dce49422a5f21a5eeeaae0d22bd41855cde4f1bbd5be89363e560e8c3768ad780e3d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6955a51be16a5a01dbe5e60b337fe317cc93c15ea206073b7f02c272ae0b7838a734898222abfb02af531f59d886b15dbaf27f9a956d921f730912d3b33d87aafc32624ec670ad8be4118d807a27869d0327328b7a338303bfaf09b08e3297cd53acb083ed0cf3d49c4370cd1a9b0776fa6382bef755e5aa5898ab647f0da3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c9964cfc16e0eb85dc62960a849e3721022c19000a6ac5665c02f708cb3079685435455451ac3ec076b24f7691b71bf2c27c4a093f464d200f47ce1666db157eb213895620bbd057f8ea41e3b9e5c2bc839f1996cfc974bd42cc5bbb5895329a5a7954182fdd8f05cb0fe690b9b005dc688746c30ffd163dedf9d4ef0ef1e7a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h334496a9b913406bda1c7f808fbed4139fdef3f4e207b102b3e96e7feebff1633e87b811159214f7dc29b2fed1379b475703aac0ae227b29bdac85391717629173acb40011da5005e78873a9a5840e532f60f3883f22942f46962d56ae27abb0868500b06862182d38a3e3cdbaae2b116de6b3c428da10e4c9ba058924821944;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h926e970335ff3fe483ac03c42848e3396ac31677605c14ab8bbc6f960583ce177ee2dbe48493211b0fb6f21f16de1bf79c4dd0fe3062d8a87fd1cff3f32efdf67fc4e8af320a0eb3f6167d0244a215d7b7b84bb5cbd1a12279b61d9f0309a8fadd8b67416f91b937dc65599678de596c8166dcf792e0c7b17e18c2a32dd98741;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5688d693f0a11ad4bae3b3d67af9ef810a925dc490ed50e766ff59104f6779480c499c150083d1d2a3817abef03f97ff0eca5362f614d83850aed78594897d9b9397e2bec82f714944097aef7713765dbb7246da153669a6ffa067d32e8da752d476a12131bf19db2479717dcfce06e193e221e432d579acec674fa1dc845e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h241c0013f22336c2c7ee99a964be77b10dd93a4df763fe49dc095c201569acfd385940339dde96b274a3987c7f31624cb5486e8da3310f46dc76f31b8f42bdcbdab9b7298faa469a8fd41cfa25c0599efc26c189e307d8ac09a164a8ea15ded33bbb04d983e98825af32b65502c122a25fc2735fc16717a8904fd2d478e58930;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46866694953b55f5e17cc91d34d2ee57a5204c7d6979818c174610c72a48ae83444ac84109d7dbb1927e0eca88535128ea4e87c315b940bf7ecd04781474b755522d01c3daf1d37c6b2d5ed2cc319c83bb1ff660cecfd653a66668f2e1a32e829ed09dd3affe048bd23ab7afe7cd83f77a6f03e601823556a4820f9e82f70e67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8001eac26f0a393a664f15030fc0f85bdfefd8224a90d50fa504c9cc968cd2137d599143ad1fe553205f06ca5ebd079c0f83866633b254132e8dccf8a116fb3c1e002bee3b0a7cddef18e34c3d2aa6d1cb35a489306304935030e2c48a519e5aeb72194469ceda49ba99f5c0b274907fd9a1c805ef4e818fc0c4e63aefd8429;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7781615ac8967fc62f9900cc90714b37c677b3ed1ca72a39f45fde32b99544637048d81e6e00287ef9d825a3178f313f1c5db03150410ff85bd430c0c5260672fc103c1bc78851b743195fb1e4d9f8fbe271c2b7778fe8a04d5199446ca877b732a6e8b68d7d2e28fe5d63c4a67eaa8c33a063a21be445b0073fd014513e3bbf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf15e6d1638fccf6f59066ca775bc06ec03d40f1041c7643ed6741271bbaa54795aec2b5307762c65e89ecddb153b964b81bc438ba39d9e004c7155b895130529745ad1bb75254cc6ddcdc0855c362d1e0b8d156cfab58697a99c97ab60eef7028d7c0ab8e0479230f056b85ccec28c339692cbf87807655527ad470e8fe6ca8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae5afb679e80641aa5ee07f7c0e32f7b6f8792341fd58110ae0da8d7862a21f9af7ed1399a7f39f24a4d60da6352f90947cae993ca75958ea634571feb697c174efa644efe9a0b3fe9494a11ba941c4ff3600f96790a06e7d503c618702189547d2226e292af69dd1f6d421b8f60089a4e89815ce0887e1ef37757f67a9fb71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95b896724e77a09732f13ba4da9e0b2bf94c2d8845c0637f0d37ae702e59e40cc8615c21c3a3ed0180d8baf6342e3fac856936b0dfb51fb8953f368b7a9cbc2fa434bbb4592f891bd7ed5e7904c28876c431b50ce5808207ac5f9e27bd2e904ecbcd16f03df3c78b8ea3a4aabeeb673b36e7835c58e51e06395eb4d917d3b0e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd602c4b229f1ba28cf7f32f82b89c64cfc4fdf1cea5cba42d06a8dbbc097274b3c29671cd8ea3c8bedc236eaabffce84f11877d52171827677347af7143dbaeb6ff48c78a381efd9f17d62330e894e2ff940853440aa37f3eb6a8325510cc8aa9ca210ec74f85961c9797a211eab29d889c99d1acc13fe46b65904330f427010;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44b5cff5db336e043a1f600efa97cff2fac774c9d8d7ae42c85b00706d3d4d108ef416d63eb98fd56e4d825f88e5f49d5606411db0682e68903b2597385deb9ef6cbb1528dec015333c474cd31bcc02402f21bcfd6a49be2955b0eff588596e81ca8aed9660e42edcda6c2b1ac09612cf27e2736f0f82050650360ce5e29cbfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88fcbd6a411ffca2bf14fe0f001e727971e039a9d272c849a21aa7e2b3102fa1a68a9bb091a074212223d5951ee6016b62261079f3c5387b9d1c00b3adf0672fc1beb16ae64f1c07d8d1a28897558d661bffb34e21b465c4ed9c39a3aa73a5112170cfb326263dad602c75aed524d5737af0dd5d9b4f79edbe9dc510d7c75a49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5afc5dca142897122633a358197e483d5a85f4c04f9a12a8f2a0a09b96ee25e770d459174b9c2c749868b2a6a6f24c43a4619a57f97e0628ff358baf5a60569556aa1be28cb7558bd43e0fd7418238aa4643e9e70d140e71853103f46f0c71460371e306e7d0793cfab26aaf8f1529fa6b58a90576f379142a58a2dc49979bca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1355f5ccbacaadf4e8d63e1c495edd44e14cd5636121252cf62bb94a90e6e3a32635332b70329a3312cdaa97c4d91beed0b9efb9712bee6c43bf6b880057eb94b90decdf1325f857cd73d3d4d6c99658415cc7bca118695fa55ebfc6844ef9efaca24ec00ecd6c88ca498fca2c379e357be2efc4466d272e239203779f9cdcf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd30636f39ea4d6145482674d9ad2e271dd6bfed5d67de8aa081b4070b10db4156c4b5fa742e19f12dd6015a4960a9548c06bb0fc3a250ffb06e63cb07dbbb9e1a8636fee6eea644120e47fbb4c52356038eada75044e1b2ab7d0e194d539da8f3d677283965b0fb49f3d71ffe2323d354393091a94cf2c347134a36556dad542;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98958049cde1b5e03d4c6cf29b7307708c43c7ef88ddaa2cfc90d1a768c203c74469a3cd7c8d74cfc7c40d7de6bb206664598f1240598d28c74b251172602ab61c0c999a131b9e861b09f55c321e11402acd2557ff8031cac8bd1688ad442542feb63a2fffac1297edef52647fd708c9ba4ad8ce20b84d3757b431857ac2b03a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2f0320c6d56793a9a6fc11e8fda04d80356260959e1deef923b70ff9cbdf598e6a4fad23804d6543db3aa3d119e5ee80a0445372e9755ae5c812af4cea6ba1054e2c3b6986aa29065dc70c2a057bff30522d407f18aa968e13c121cc8c050cb09b1051ef2fea5da4908e4fedb156105176fff3c30eb94a68041222d30c8ed49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a0798dd80795fdad630bf72c7b6d8b385ad748bd9742bc78a80e0aa8e3b6dfad9e5bd41e7efe18806037946749ca221f69211a6856bc0b7dc25523c7794346155a5fb786cae830bf5fd652251ac804e00356cf8e8b900472115a18cbe64268f8d24e4b6a6e674711d71581a57316b9bee28f12a418a25ae3fdb76a9afa5ad9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd43a37c6070747599d579e70039b335671688345db674e064c224b493bf8cf96848be5cb8d40c82d1eda555c9c1c999a277b5b435de145e0696b0d48a10389e722120b94214aa7ec1880dc75887fa5efb79fc895cb5293a9ac8874d73be42e2a7b104ef76a36880c18127711633626bad8e83088817ac0f1c9954ce847a93b85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4ffb62b05ba4c149597216e448387f263cad3590cf8e29a0e5ac30c650ef53a013824a4eb788d09fad0bf4ed0f1567e614851d60ac91dfe696c33be2c4221b4ce477ebad1e6b969ecc9f6080cf6ab38d57e770427e60060fc2008bf5d32654606b1c6cd7ddee2df7bc018e82536f10cf4984a36d2712470557a7022d7b9f80e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha56b85ea8314df90c9bc7189f4b0b5d034747a60b065f330933bee8f518aa627abd6db6a47db13427759a92deaa94470a9d72532384e82778ae16bb63b8495728f993b44c8f8a38eca1e64e9dc65242fbccd14a245403a2bddede729f06fee48fcc9fa39a04de22331e98395cb3aa33c43479e9d51083ae803b63d1e4146c141;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h759d173a2b294fcf2414b8599043e9a8238e4d95378c494bec7d9592b6290a1b899799d4655d7f984cdddb16a9541920570f4c8f18b6bd7527d88d36f78455e89196f187139f2ee2c5bb7b2808a2329f8e4e66a41a0fedf15e95dd1f718a7a5a131fc60d0b7a1733cb2f805440c2706052d6f1d6538a0ff35a3f586ef7fb377;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43f10a7875d43e7592e4792abca487b3f87d314e62406b961c086b18a8f4bfe66d0e215beee115f416fae1445386d96b9e84991b34f59c5cb55753c178561d240f97a88bedb7b5cc6f15a75a401f6327cac6eedae6c9f531f39abdf2c0446c92220bb617a2747df5b8520fd148fd4005eed274a33cd100244298c6abe78b4909;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h264946f6afc6dbf6832b592fd1a2ace042792c1e13451ae86aaf5d4ac3654e6a267da06acbe1281f5764b0fed4317ca81d4d24540e8056e6fa53e233fe3fd1bb1f9b648ead78bed4654894b5d36313ff8cd252a002d0a264fe2d89e87dec1dee00602f406a5a035ae142e31a2a0f4f002f477d240bde97d9e5a87f2af81bae61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb00ef10650e56fd378193124359299f6720de65c93dd7e4031231d058cb3e8f5cea705d7e1a27c8b265c659d354e4f3bf235320c1d0d140c75fb9342dc266f7b9308391824a41b8efaef848fc4ceaf4e9e80b9fe678f464a8c292217ac6a681b84ab8eafa1c281e9b720ffdb429ca5651da7bc035a7bdd51df0ce3fcbfefbb73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h125e3138a62d47662af39681e621cd165c21edbde4355d4243e18c75ed9fc4548cd76192e53b556d67f697ce4e0c3e54da12e231b082a0a7b456e1145905fd1e42683456205ffd331a17e4e2bafacbff492e204e0b47049b1711b8812ec4372e2bfe09e85fdce0f58943c2e32e383b548e7d39a5fe8264fd0f1f8f2c0cc19665;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2500e22861e8560748144e099c53ae45ae0a1a78d73db026ab60ff3c9c0748708d588b11c260eaa7c03d9cee0dff6b17a84630be447d56c3903d46078aa679ffe0d4d221745d39f2bd30a3f501fb75f38ccd6d80cc040b96ea9ca1a5f7fa23c00ceeed697a3ee0ac9d143f419ed060794e456ebc4397246a6bd1d97d6c203ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h614d497611bbfc836021efa2f92ca42d8e7742069b2e207e1cf0e372ea427c2137618c927fa04f3edb0777e275dd0b79fa3ecf1f73e1d55c1c93cd447b3475207714e8cc3ed747eddefea7be96d20ae2cef20548b9edf6b736b3cc10beb9cf7a69b55ea81b77355786bd193a1d7ed961d22c10a2ebf35519c3fae3f4b94b300b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cedf7f0eb601e0e1cf6b45e3ecc92df0e3a4aeb9b16f3b8ef5c7553e39f96243b64d46568aa14b564fe069f3110c7078fcb90b03ca84b7ac760e21c92b56727d5f63c232a441b9d970c3f6efbe8703f5a30dba221308920a5070d5cd52dbae8c99c274f5350e8702813ae5f28328235f1b842e4cafc52e83efbc65f3ffa40b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e5145fa487113843ea61d45a79c2278357183da76dbc281a02b348f7d92463bbd2c49b597f575b65393abac5e4fb331031e5649a12f6dd56cc409173b9d7fd1f2e1ed5e4060db85cbadf3b55e08cac93ff75b3c754773a920992ca9b9dc07f3af384fc915652f2a302284b87aa0fc5ce72d7f9cd990493171c50e6fba964b23;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha14b423de07c2366deec37d5ec931d0697d5474d3f1318bc7f6ef8c127754f0b0b049c2b244cff90cc0d5935c63a62942a8ff5bfee5d4174448d028cd855812f7e0c87e12bf85a1f42361fcb7e4e7d0ad35269747bb0e5f7d9166afe758685433220b5cd2dc9ceb52f485e30d715d61c2cf91f69992659fd99a601be85706499;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35cf068fc452086d66e9070c0868003698cc5852a2627df51f7d1965a20750e26e86af40a6cd2762a6921d90f1a6e73f69a4d3e85b001921a88bc5a4f6253799c4ab5475b27f889dc7f534a166718a730a195af6304c9f2eccad6affd8597f40ad20cf1204284a03e08b6c9f1902150bafbfe0b4bf6ebf20ace814b5185be7aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31348ad4f8a7cfe65a7819dc045770f1c95fb95c9c4d0ce2833813a0755366ef3c840229a4e0818b127c1b5182f754db7dff5ef38c6382d1a47139d5ee50d8b294fe000a44016870939b9311f363b9e187ad50e3813b9f70639503bb11dfb6afbf40efb1a15b7c309e638bb28a661e2f76502b2f13410bcd968f2898f27b8ca3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69dadca8d006f45cd768db1cd3246d70d7211b1e87e0199a5acae6172b6cddc79062bfcd720607ae555ef7f7c50fdd6b1ed41e20ba224341cb0ca6aa7da272b4031726c383704eac91e3741a0a38b9438495ad5a2d321aa4cf231ec4d1d0413b24f79d8dbd0daaf762768acef89fbf045671caa571d410a14b7b230cc65dc6e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4765a7d09237de4cb39147111f51a8b2fd11176aa8c6561519259beabc20c5a3b0c06b0a7ec0b44f30350f87e8ebb7ef70f75132dcd3e1c443be1f31fddc2f3cae2aa9c710a37d7c20008d63b6832b9529a3a61fe0196a078eacbd6c4d4dcd9598e49371d9db083bebd3fec208e1cc6d99a06dee98cab24540a2bc5683c38e1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a9ef8fa96545c25ca234529fbc54fd6c4583a7807d18df0491159e234bbc80e3b376060108207d7815728b4d0c152ba58ecf742a451f02021cf4f83a7cab7edb299e75215124096db3dd694922d33480cb269f03e553ece12181f6556568e6a765618dbf85b54cdf6be3c896d9a1075056a4f205e66a2a05b7708595c953d55;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23a10f8813aad34c3c8e7d0c549d710997c682465a9832fc68a30cb5ceae7db8e3995b5261c06d795f1caf5e3696a59d69d1f1df5b8d155595b0fcd23444c6180c8494f3c8a89897dd6514dbbadcc01435bc26262ee4bccf2ecc83c2cf94dcadcbe06820157b2cfa8eec6a021768d5899ab634dec185447e92622392aaebb625;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70d6b0fb80c74871f6d214822b6bfdc3ebc9833931b8e6939c4046bdafd33f1239df1bbff157e0ea94b29420ea70b4d2915ee5d244e980746c492e1dc04b51bae3502792809bdbf8abecef3bb38ed9589dd8df56d3984d21c5d0640db3cc8df1541b36978ef34360d73a9b8eb9f8b178dfadc16823b4262c9ab87a18e66008e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h847a43ce2bd9526937c3bb840da7d093c7beb54f800fe294086bf1eb0a0e6edf20e96c56958e4ab285f82328656d0c7f9693466662c2a63ce9d65fac5ea394908629863258965adcd5e5e97cfcf456ad21cac918911a53e5ccea4fee1ef35bf5583de97a785f584475dc9f59499e99eba94aab632834bb9fa50b27871ea8f08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7961cbd70d668ae3758695b306db4c6c77a55a45e94cade0d911e82508f416d46ef61955f9ef8d598676cf91e110731a7758b2585e71dc3f755b770eeecfc087507c3e55f49e558b324c0f8e6f84ebe989cfcade7c0558617dd1e717227167147debca860354a7505c5c471a8aeba3dd214f395b3a1a006c1001b9fadcfe4823;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b1b7b691037b9efeb3fde8debe19aa6fef40606456c8d4e69e4b4b61858e93247c3880818d6cbc0753d54fd4ca4b6c8997774e223aee4ba1243bba72ea5b01b79f9a38052960924a214c1629f314816f8b218eeb3e4a9aa3ffb6990767776927280435ca7232a73430bc922b974966d1f1c332d3168b88f902cb5723f0497e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97feaae16e1ef87aab56c8172d1f27aea2bed73c11020d7c5edcc42e385bf8b8ebbd43f94c0504942d52462f787f4231aed6f60618b9561b6a99ff519297b8fa2d0e6eb8c778a7875aba80e4ed33712b03991b6510d28d823e19e12c52cb826eb48826ad48af8c1c8d2c6752e551a5482fa8edff75a7a7666a9190f75d0f7e57;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8710be777cda034dde88ecb79f5617abf6aec593234e34dc791ae10669798adb4756844095fce13a2d4ea3a60d3d93578c3d63d7e2af18a1dbb2cffa5fa3b1d499077806f64c7cc9cad5ceaeed449424397b3632ccd65c51512c15b18f6a96acab4aa70e941e46b9f1a01de1e302a663bc0f9c52374aef93eda4cc7a932d0980;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6df3a448c5dd9e9c7c6f6e7db7567df161fc730d7b20dddc629d4dbbe3f2e6b1716e011c9f898d3c8e0bcb6786e72cc68a11514a62dc368de2ec80f24dde2f907a9fa9ddc452eafea1236474a54a7850961e6cb59b3302f886f2cc37294a4b1b9abc3fefa9c5a2459b959f6593dd50b83f19149986ce7d2965d55000bc9eae3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cdab08c649d46ffece8f6e7ed8013d5f966b48047b4ab4df6886adfe08ce6700b7bfe1ae3370dd299528b9ea0300699c1e5fe1febb564083978713022c4ecb17cb7bf1e8f5d3ca19bff7ba231e7a5e50ff91730eef96fc56152b2b008620455427058b4504a504e9b3e65c97ff4aa58876fa442323a9891bb06f1ba1ec45b08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf070571cb228fdbeae160fc95d7ad8f74c5db6cf982c6a3dd9009209ffb458bfafdcd363cb298ac219cc874bb6ed1b353b695ffde5d4e5b56e25fe4fecc71fc32d25d17954d5e96d4cdb3f6e4bff0b5a6b55ce4ddb6aa672414668a88d87125801bda420e83da54f8e36a3f0d88dc233a01f10ffeae2fc0f7a908aafcda6548;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc44235eff122e6b81df56cbc251ae50343ca96164af55deb3c5dc91e0f980ebc5c579a1251085fcc4c44134bddb0ffa3a202c99ea109c9966d68bc8c58d5c879d5e9f7f8c5f2d4bc8a0d169af302f7d95ce491c8d4f635553690fcd5d0ae7bb9e69fb7fcbdca184ffeb6cf3a6004e3e05e7106bbead9bce914638af56c957be5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf55a9591afca4aadc49fd7e3fd8ba6aa4bdea0e3d071c35407346391545076126d8805e9b468e34cbec458fed4b3a8bdd008166106cc8aae263d23a2df7b04e477b70ab7b082e0a9b0c4e9fa1bff0d7a97e493f06e063b9659cafe9aedccd77048183a625025edd96824d91aa60974d890efa3c98cae0322793fc82d8160db3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce6887d45bf97a77ebfb2e1c8f9577e8fcc87b31e951f135249917adad49a0bb2a1f39ed0f4e3971d8e647779ee8b4f6a620b58e4e148d0427592c66a54f341ec287cd6c028319b8372df582da34403c98869246b688e1af8d1f2e1dec70ebf800bf5da7925e988162e3b473270d4e58ec037af94987594401e0496d22d2cafe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dde0043ea712fd9964c4ec1838f201501732245e0658f77ffe08f0ed50539ef61bce198ba8be34390ed08bd2d8ad281d18d6e917d5143301bfd9a6da44cd6300f244c0975e05c0e2b8176c43f8af0432495b9d0fb0a9b3771c3ed98fcc19a579b0401e702cdbabd597165e1c9a9dc14a983e09d28452e9713cb96854f9344c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb18e4e5e134a3e99c7c575e9ef4084ba88408582dd5f9ab23e441cd2653c0d5fc079a52c9fe540b7ae7abf8c819bc8b9c138cdf529fa34cfa4ab40d20ebe5c0386a4d91bc05cab56e133854c556035e5b12e42d337c69328ae1ae21008a8874f66423fcff4efdb0b661ca224cc38e4c598050205d9601f9ff37628fcf367e26c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f2eb261ee35161de97520138af19599659dc9817fe1e126a39bd198e5e23f94939fd5566c357ed3102c0010f427fe17fb8e5c805c01e2be9b9fdeef23260ec1f905374da1ece50a11360536b1709f83128af1b57b6517f27e5f0afbe37b9b01734bf55970521e23946d977bec0b4aba3d929852c1623ede1d3fb7d985ca346f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a02aada0170f1e4fe3ae309d9020092713c66feacd00cd0bde034502006e36024a6905221889564cdf722047955d4722194bc16688815f446c467ededf056d5c96a304a7963529dd353322ec30d5e15ae9dec80f61ec511e736691a1ef8b4a301907b8315e4fea1b385cc28472b5cd561e701dcabfeda095491ecf5dd8875f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9a1eb2edf5d9f7783ec72ea3c06e2a44a56344f2d3f671be58fcfd62820764b5ea49b512e88a8208fa77fe0b21ef1e413b9485d2f0900292ed67e2f6ee085b39b5995add724f9747a0128b389fff8a9e74c936d47f06d6502b919d4c11455ed3d49a29a448020d45569b40479e1ed6f103f89c9bb05bd015d9a56bdd23dbb1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb442df51e30179bf694d2b8d34cca0c0bb43f61fe669d246ee152a4ee8414defde4e0a5e3e73b6e79a1aae38caa50fc6c33650ecdbd1116935265ae8fdcbdf2bae5c95bf54dc12a3ac0350537ecf07bfa71cc01b9a625fa91c3b43e99e534f9f6c5edd2170b0993c6f7b7fb8abec2120b191eee44f377395b523800769faa6a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2f38d2a65b82abff74499269cc352a85536aee87baf1fc5a91e71e87743f188608b2684ed705955c47e30a42606ddba6681c4533f1aa49290dcaf180bc366795a3356f67acfbb1e488e4510639ae5018d76446c9d6c9546b58b77bc9c22082418bbeb71a84cdf2a2d19c1ffc5836cd121f370b990f2c4d0fc685e7fca8c8815;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8384e65fe1acb2b9b626dc3fda125d8339bc0f1ae17b6f8295143469036eeff32929143fdcf08894714269a4f9b7216f867d2faa849e7e4387cc8af37df66d45b37684b1f8cc5c50baf1f19ce97f04ea4bc1d6b0748413f333f740f8c1b8f8fdee360b9119cd125f7346a5d96a629d22e99254bfcb292ac997e2375fac733c2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2aa3d4bdb0fa417af46b456c5af165be11900f1101e1400578dc19db1e2c6e9d23f96322d4c12a47613cf0b795ceeccbe016047b09cd11b1ce34e62d2b9a92f6dc24e5e91c7534f63cf69399e9a39d992e05b5142a515dd1d8e173531e015b8fef55c10d00e804f0bc097a692ea0ff8d2ef016093c8d73c99fd3f92456bea78;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99d9986aef1d1f09bff954d5ef74ab69cb95c6d097985358ec1d88db5a94dfd951eb269c0e387c4dbc9150a50ba54bfb7cb2fb46be333f2e395545898746aa2bb44a0c59b7d473268ed914cfa32d4c16892cbd1cd88320c0562ba5d5ccc60a5498b43a58df256556f373ff3f9a318a28072b34eea05055c5d0f02e8552466644;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb144dbb9bcf919042f4994b86caf0bc356457dfa5f618069942ae653d3f45ae86c62ca5ea5f915f3ca3abb013c1fbf9395af041344b61f75f2e27ef0d9906ad59e607870d21c8ac0453f1d144a5308315eadab52b47f29146dea10bf24d198d255178cf6951dbecc1143f122359254d371ce09c78a8871309eca337d4eae9eb7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c6ccfb80d4fd981266544fa4e8c183d137003e3b23e215839037823a17b52316c42c8c8af0f2b1e13474117ddcef0ee27a7417359bb8da568c0ebf5ac4874718887b99beb42220ed6d2202558db274008928612e3ced8770312552d0382699f0f4a3113a345043d41aea540bcf399c4de95587df5cfdf5fd235a7080aa43246;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6381e144ea806dc787edefddc0892603dd30714930768549ef5d8bd4ee96ee58feed965a39884f72cc846c3ac1ef7294bcfbf8f181c9a89fdc71c729f92b747431d9c416a21d655ee902f0872494a09db393defde40cd1ca4077f4f612864e48ecb4c04444fa3a181f4086f12c1e41ca52cc05a808be999224836445e753a0e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b5b1791df15abd177944bcb87d8f57486562aeb28c42395d524841989b0bccf63e47bc081ab284c821de48dfd3c0db3a8aa8c6cea3ffd42c3e98166d79615b7d7eac89430d716eb24913ab68382c83ad7117540677daa3bf5e5e3c8594c0e774ad1810ad363c9b39f6aad5ebab785d4ed8bc191ed17821297a03da6ecc781ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff96747aee8be8a754a19c140bfdd63b8311f6a3e96bf14b1c749708f57871ff13252b49008b5965d31ecaece812c8cf1c9f187a6f370a4474d079375c25c37d7fae95be1ce43ab6b6c2426b732d5e1f89cd712f18de3209a25a522460f4ef332fac0974ee8f10665b3581c577dee5d8921e54754528daae959facab64642029;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85d2f6736d4d72570f1d4aa72be90b0734129c0239a5c64a47589752de00e016f2bd0755ec35a8786258b1b2ba87f2814f50c6825f72d81bc50ce2443eebd919971fb4212e2ce8e41347b13d8728ba43c0c3702ac8a4badaacfe9c7a7b8b0cfab59836c33589d2668df323f2adb40f8c6e0ef7b6c5ecfbfcd61d57f67379dd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37cc98973b6550e74045ad9abc16bed8fbdd8fd25f4861c6aa58655ed930039964369777c22e4478cc9e2bfb1174a92955143d12119c52ed1710470b010236cf5e0f8699bbee899145730498aa50e0271afa3c9617f15de4d8a11cc25f35e1371f03e00de8c5a89c2793116dc56c219ab0a7120a20b06b09f7d07c73fd6f9f5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cfb22847ba8d90571f92bb6630c194ad990d92dc475dba73cbd591db37f9d07822629e450f2fe0eaba8e21d275a7b824de8d0b0195ab4188df0cdbfb0272bb5c10bfcb15b49a487daf382870774cdbb3a1f938c734b3da552e9c0d452295b7ef9f04493ad13fe99a39acef1b12b84d50c94a3e1fc846ec56694ff596cbc4f04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c0401a848766375eabce563f30603f66f74742a8df7c3758fea16e40a66e2a5e87c88d9cd1cd298a3843c4532be830590eca71e4f94e8b8b96097732c85f56bd76864e6222626309895a53189f5fa2b492128248a0d1c5a74b67032d3a39437daf46e7d1d2cd7be06f119fa87e89d63ba3589766730feba886363d492334c21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3345106da7196cef3abc629188669ca59500a43fd92bdf35746bd6a3c6e92a3b0ec7f935f8729b68a38580798e561c75255501bde09780a5018a7adf237990c5ad16b88b73d998a0f9fa701d93c0e568b243fd7e371b7cce0295724cbb9165e2faaa77b110e4441a53fad0f76ec24160bd8f7916db45705e8b8d288522618c8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h744d61a87887705f798f4bffa799f064d4b0e72695a67b38b757b6aeee16e891b90d3ae8e9f4e50009f569d098f58a2301e9add3d97254e0da42035fd8e9d613f76bd821a5b84394e5f2e57e157ce538d6f1cbcd1f6f1ade62e029d29b47be31d147551902891e2cbee88cdce1f6ac5cf0f58a85fbd19a5c5425862e2677e490;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3446b54b21712e9d2a4bb707fa0e86b68c09aee964f31b52f67edf0595924b8dbc64941817a4c04ab7b034d7e468a3e821420d5825287e1525df1ed9b902e383e021f9dbb3fb01afab9b2b906cd99a88704cdbfcbc92cb9f12bdaa2636e079d14f6a51de342118cd93d97c3acd601c56e6c7d87533f82e0856ecbfafd3ef8767;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90ecabaebb73943cb26c3f5e938f440a56e6dc4445fc228a0d670a123b660c39b7cef843fe2235582c50fd250590fc6088a5c142947a2700fb98029e2b2ccf70a0397f4998418c2868623d16a9ce3d6004039491c0a105d54865ad36df509690c29de7313552d28794bcd0d53bdb795896f4407a79f21119b15204b6af6d3f64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25dce8dd6c682b5461a9ab840f720fd31d1ad2222ff02579cfa1d369027c794a0817f1038a099f2c027c62b222b92d5d7565b23e3acb0b9faec02fd1ca6cc47cc119d9067fff0874659e76d8f9d4920a94ffd2f75ae9d6d4cdbc9999b3e906c65f69bb3149f799606deb913eb798afc9de0ec574aac8cd69e80177c6b4dc60b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8051e87e5919333b351e723daec749d2b0187a680e45e4bff967f5b5ab3f7defc0fd17b49e4588e4b031c46ce95cf7d3521d2f8c884e8356aa8d07554647bbd3b4daabfae303a9e1485f7b29dc6d177d76a7a9f99beffa90c6d2e700a3bf68ae1ad48e635920dde6f72f84819e863763d1c6baa642b002ac2168578e2f090f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h138f078ed17fb75d06704dd5af5b97b3e2ceb63285472e4c6e3116afc4d32386d12b978c75280bf2cfc8b0ff0877a8aa42a9adf938f121c3523c14a5ed15e91475e2d6c186972b5525c5d415548bea755407f291ea6b5ef7870d82476543f7e85e07d36f6c16709d8df9cf1e654c7db88f5a3d69b6d1875dcc875b7876293028;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bad151a2d88181c9f486d34851faa5b9058e6fe9188596d642e10e26d459024a3e99690c37d347d8060d8b5e729fc6f03a033012b05c1ee7fab01aaeea1acc7a49b7775e8e570865430d5471f0e20b1d594af30e8f6f847dfd163dcaf0c68c8df157edeb5fb76d3e1c44aae9bd8ac9c96338aaf51b6bff42675ff0520c151ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7de91a6096b04bee5b3c42363af8f78cbd5c3b8708374cd8ad9355e3a06f42594593b55466e6e91b7323ae22887d4dc09ce9198545fcfd4a0b349cf1506c0fcf2ad0e0be0876da3db3091717a9e3c8087723752c1a5778adba845c06474d93e4afd0ec6442dcaab3d986c8120cb3eb813f0af81184244d4994c53a40bcb549ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f4bda9c09ec5c40c73ae33da5f19e497a5a8ef0a788690491c345ec640a8ab15037d3f2282bd7d25a3262857eccf32849afc8262837069b39b5ebab728fb7156681555715d0c3c0477d1995fddcd8ef9555f17bb2ecb39b4e766286b541f8c60149b126f3c71b3a58b00afa340a18052ffb7a557ee2566b161fea1d77a830fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45a31b84cad51139e56a9b4c49b2f04fd132c73312083583b0e10543f80a7e7067c5490536744d48cd955459e23db6c34bc280710eddf003eb4722ad0293e747bc251fe3474258b0c93b955dd9fb025812efeb4cc59dc1cc1a85f8a7ff239334ab92137407046f29c2e0aea91feb4664546cdaac05d8346d7a24e34795a681dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdd1e88ff109da8b91f1103d92e20e0284d48ccd0c3d43c4cb575b17e84f5c516e4eef2dc0d2a5827c754061a79f8ba8abab731a2f41252f0bf76c174dbada39d3cc542c984ef40943babb23a17d14959b0bd0e386095e0c7114acb416c3e1002888055c945eeb560dc5b0ab14fc4a0f37aa9d2398a6c65feeb4f60354292707;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6830e0df6f52a00e79f1bd40b00f653159802f67004427a91b4fd7f77874ce76fb036823173d37aec6564b2f26c6fa9abf088140241c15aef2fde790b1187d0144c6790a09315d788696b5367a62c20f812db2418780722c46e8d808ed0ae8d41aef6070d2abacc5d5a06efa2537e48d744a94321a38945c9031f076abf2055;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d659ff497bdd7c4555a222e6062a47edf132907a3b9b91eb84f21b6023a1fdb2e48cb9645d239af47346d554684369cf6631dff77b02a1027d98e6ee1262c3d8c7426e26f1092b2d080de45b9b06ca45f9ea95a45997f6e8b92185a42f686cfd7d8822f8fd2fd573ec89a3e27168fc23b63cf4b4ba152726fdba73b2541198f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ad03e7669aae01a4b7206420a7322173a17a7117c1aa33b2651e28bab8bed532b6bd594d2e8357e1ecfc8416a2aa468c80d142c91cf366611f08e0b07d42a50a5ba81371afb3c71cecefb12c0ab83ca24dff84e65037f1d1fd661f38a9246fdbcd85ed112837df8af9e1f4367c753d79e58387120eb6afc01bba68c1d7bbb38;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3993e3046b5a1d75140bde2fcc87658f79daa3597b62ddbfc1952a48df022839d14e8d56942437b1f558ccbba1afc420b4e343b9cef14bd2bdefee84c071743cf6542ccc40375efa28d3b7ae8c150ffdcb3d1c5af416386cce2d6911e276a371e846564da589c4aa577ed0e5a68f7e5d537d944976ae8ad74fd4992ec691d6f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h501eedacfa63aa69ca15ff619a18053e8b3436f10ac1bb4217c863950a57b4b55c8e7a75643871c42bebd612e78fa4a0785a21c7acedb6da3c4ddd0bbe42d6b91a56d25b1c60515c0f3d37603144162aeb96e794c79bddcb9b418aff9cf9240f4b910246819bbfd307d40659b62b89833f94b932b7dbf638ecddef10efc8ed8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb54e2743d830e6a47bade959b0cd773ec24fdf66297102ca5f838f44bc9691ecbdd9928c0d1d844c291ea4b0a80d8548c907bfc564650bc3fa60f84f83fb572e8c9eecfb30f980b0b0a8989ef8279cb20f15d0c195ecc59cc00ecb4fd9908137d5563fb444299c3eb9172cd3ba5dc2903e296570fdfb34dc0316f23dd100a028;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda9a584fe9ef1291a8b924ea4e2546cd797d6db03e97b454398a1f4084cbc8d3d48897c1de11089442423bfa9eca74ea1a96927bebc133afd8ddb9d612aa9d493233d9ea8c427b1408b5b35d9ed3964c1bfac9f7cc87843ecddcbdc4994ec3fe16a5d2debfd166d3d3a61098eb87e05dd129b0e064c642c4668a9953c2b0bf6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57f8ed656c673db21fe161cc5adcfcfc368cf45c82ff778cabe266ce7d44daf9a20fe15e85a224eb157e6ec474d13df0b5dcf3c6ce0f46894c2834e4b855e8d9f79dd44e90e1cae188f1ca82dfcd86b631aaa390b61df7b48deace71730586040c9af2f02391df1f3f2644e7f419088b66099c20a66d8d3430c3496dfa918bb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44b74fd9947dbce465edae59de447b908d75b5ad2fc75fcaf428173f899033d06b39c006a041ac726ab31959b8ba1f5cab05b03f46178d7473866597e9bb423d94737e41c446d43275878daa695bfa4e929b2d4a1cf597879649fdd94d05fdf5e64d5656517908c52691409aad612227629972733fea7662a5756b7d1edb64b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bfcc32e0c75221d8ba296574fe006accd24852fd16b1434ef624da8b46bfa8f27a4372a76fab8a1cd3a96de5a4f94e3911e0cc7b3854b8977c14d99e8af960f50f105f15e069181504443f86062c4f93863b47878c2ee0e425ec623f08cd84234b57412b97a3e2ca9a0faeef29e608afd294d634081926077c6a166444d385b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e6f33a075066a681d714b46a050077955740b436320d273c9d7401e55e107d02d0aa70496a135341d5c1bc2ac3943083fc4ada5d4e9dfca6b4368fde17569b1f92c17e8ba93837f99459799b6ee5386a67ec47c2a847b65384093f51827afe6552f2309745e04c07cceb792096e4de17bf48b17cdef63ff4f96956f22cb3b5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbc4d169f952939739ddeb0d0af712a4c210537c91b7ee7fff3539d445302bab9d6b8e8c50b60e23fb1c414762c6dcc5d2c206d5f9ee29276a98325cd82410ab0849eaac8cceac118b7d61edde3c912b47eb82da08b4c3dfbfe0289d368ac690496009ff3a890b9e73e3dccc4d946fcf1315bb573dce447087476450265de3b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c3aa11717f5ddc84bd581da1015053bae188dae67a7a6b1b30c1caa13d5463fb5ad7913063339910eb3d18adbdb6796c92fe403d043611aba107feb197242c996ddba3790a6e6f6ed7c0340b418fe7bd7c758d04c7dfaedd2640c74f75e4b4a3f4df2f0d6c66a32a22677f0d6bb3070c3096ad34dbc85f99e740c4f33ab53f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf39d193d21c36fdcfff9af7dd69edf9b9d1409dd3531fd2514d6bef5bbed0b92356d033b7e499d459a71389ac6025d7ecc20cceb2f1e5218e265ea59d79dec48d780b684dd7ac6c61dca81856b43dc3b3382d13febd9a018c66334228ac215b2e16372d33ddf0af40512a4b363692a5c3c8f4e82358d048bff6a3e9c913f5400;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h580a23f1df58d4614abd95ac0eb743aebf4b05a0174af255a2be2f3c76fd40be7805e0461c797323a31893e6b9fa3f165e9e4aab067388cc11678498b02446f18651c6d3374f4978e1b6acfda54db8de1985950a9e97740df8ddd1e412dbbc65d34d9d87c1b3da736e9b58ce53fdbb2f83822bafe20e8bca055022b15713914e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12d58d7bf29782ce219b83e44cddd0cc212d358a9f643ba3697cd86ac5b729ea1668bd781d1c5952474f9538ea495bfa941703ac8ebacaebb2e36317b32811dc283cafa73c45ad525dcc3ff410a5b9f13dc859190e1b66d84a1dcacb7539d7a2558f2cea8f3e68b4000e790d4b975765c783d422429ce92303edd813a7218a0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58b254808eab746dfcc4335dceb3127361d346a2cfd1197400b8dc278e040d7dc2ca95274c188f2948eee1887412990265b80f85cf297db5b02fdb09b193255f4c41f4f0fd908a8caa20da26992a24cfc56c037922bfc4db00981771ba72ccbfcc32a0bd4fdb83aba4619e89608570d4dfee6d336727027cbe7935ec6fabc11b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce6651f0767c65f1023740a3bf56621c83389680e211cdd6ab2390afe48fc24025b90b943246f242eeb71cb4904266d13645cea1b15d82d6eb1a87f3f48b729e4cd8a4dcd91e0ec2471d1371c7aa0a343ad06faa09eea23e4837ae7dbfddf6c1fb606c4eca5f8a9bcb21c3af7d4578f4fbb9e34806445ed881635c63976e1aba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab73223f6b80fe92dbf947e0d87471171fe208a35af5f0c350a1c4b46fd5d115d8b85eef90a98f53a90cdfa164c23ff2872a05655af155ce038e584275ee0462c8a35b6469a9788ee7872954b64f4d30bb9fc54fdde430d2cb3300a1c8eed586d416635e1794f69b8c778a94452a36a07250649fff5d1438469dce457939b6c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97557cc382b4da9b35abac4013a8ed0c8d5a290819c79fcfc44690e66f6b63df2e36c613fff57aec5a5e07aac00e21cfe29f4b1e6a2aa03e1bf1cb5ca1f30c49780bca705ed21bde9987827819eebddee75c260a53c8ce8609261c636b19ac2e63ab1b2aa29c3c5900b0b1aba1305e67e4e75c51a4600fed658f6407740457c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66c684e389c55192ce4ae063abe61cc853d86559dcc2c7518a62f3d1343b871b05c6553e761fa51c75a038c9fe5f64925e7ac9635f2705fe7aa40bd89d202473bb0df148eb9f46d99958fac95575fe07594005952f271d82f4f1c10febf99beac469d12b770b4759a3221f93136308221f451292ce05affe26eaf3cfe9153f89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e21333d88bb63c65bf4eb07ae92dc5895d2a622412afabdc95573b6cb80bbaa599e1d0c46e374de70942fc060046b882af2314537cb3fdb0ddc72204e78d23eba816f3c8a436c86f94b3fa3ca6186a7f67598eafba1d66febcfc7cda6625d341b8c313acab2dce2c9a11b2fdd484cfa1fae4ac8fd1756ebedfc385f2da07155;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb48d88a7f99ff7974c26079e381d4d0b1a9b01aab680886da975787dd60c478d9398405fe31c0fae01a871368f43fa164d181ed1991da7c4397801c2989c6bbb12d4a6f41194212e307a7ac1db2641a0cdbd809300f2524a37672bd33002075bc4fbcc0532dae565d85be8d5d1aca992cee8c6571f7ea2245dae3a78cd316b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78a276b9506493ad540ed7e28a2d83128bb43dc26dd208108d12f466ffac8385c139b3a9902452fd24fdefc18a80412c44571268f8ccec7c5a6fc77f99ecb24a02d4c9c356bd3fb3205dc0debccf027adf4261c12f12787242570f8d51d6f31f7d7164bd82bcee46c11e8d4421ba762f3a228ce29ca2e3190a6d4aa85647151b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2671322b41c8daeff2dd640ccc2dc43aee7dbfae9ffb6487135dac7bc153b52f02db27485c771bf5952aadd965fbe09962e1d3351263626c643fb159478b0069d2c43b78c0ee47ca0780acbc73d61840bd52a1412829a12b98bc95ac62c9d28615c93108f4f9cb26684772a1275fd7ed488395d775c5f9c5cb21dd5d8c225d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h160a4035183bc040e7132a779b97b9feeb4ecb79e317830e7a95fc693e2e3d588643ed64516f9ea51d2308ef19bda55beee1f21062941a1417a8d65fdaec06b1c346189dca109a526c33d15ab26705646aa9d0c6ff04866a5b8d938c94559128751c7ce84ed6d5417b4948cef5b310118f19118772e20f98c90251c6d7a23233;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc26f389d0369df98b588d82b407827716af3c99003fcc5d7e308ec1c41908af0315cda80ea1cb6f20afd876e5dc561206e0ec17c77cc892c8742bc4002fac14b6450f91ccb3539d51fada4c8b56b2b5d341148558baab8f52d63eda7cc98383f84795a67234940973f5442c448999f88919abb7eafa94c71f2ebc16ce216ca81;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6829e6d304db43589af4decb5f68cd1e67501e201b134aa32d5f03f8e5b2c95e141e99257c6fe6f9d577b7b0e35aaaec8a89915f432062f3ec631f9493d80a075afdf978d8cf742a886ee1f32b3894f7f35dfd99c3054a9a4aa43f1a76a7c29549bc68da74e387e4d4c39793587168d80e83e013d8e511c740d9a40de0f8c28c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf4a969a430d442470bd79ad8ee196369fea065019964ee1fbf7e48c3a8a84a1a0edadea9cff4c53dee30b14452376dddb5062e905a695136f851ac837098f759b16ddbec92d36454f56f36cb09e407e6d864da5a8480b9911b5664fac14e197fd886b5b8b9e4edfff667090fb671c1c2afce6ea3d7e0fcf7e44b92dbf863e5f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h838bc427b663fd076ed92ef44d6a1a246836ce7520300d09c55e702ac09c4e498ef373c2df199ebbc2a9c2e9a37adf410c2ea1e7a4140c531a20933dc9e89fa623620868e89f94bdc17da2286942e2299c6045be11f09895fd76746fe7deb16ed49741573f0b16498fba69adf7c13da2831f375adafba7905612c5874e7b7097;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h921b9d60bc9c112269ee133f51318bb7a3e5b455176abf9639205af0ee099d6b7e2694af307e14b93721fb7c0401595a1209acc2cc8a4b392b046236d90db8c8145d8d01893ae253f0851497a26bd382d0136d7c1bc34f872dc78ef21fd36a03ecc219f21d572a4a46b73af31beefa88cec21e615f1a87a365cef319715e7134;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4cf5c5512256b1d757577a30b0aaadfe834511a23325c76430fb9d3390414b57a9d23f80e7c5acbf0e596b91fac3cf4ea14517aa266b5538accd0704d8154749ff968d79b3d0c547504c595d73b8f9c4128c6ebdb3672e6c858e8e554c1363260ccaf2c912277012f5c93c7752714bf7967e1277d1dbfde5ca633063c9e6633;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc473930a495ad028abdc51bc0a769d06bfebf9072f78c77c6c83d77dfd0c0bf5e88ab6dbebbcd8cfbefc6e28e2f293fc9a1fa392e9890f7234cce0dde7f2fd3c69e4eba428e47f3a44c55d5c96ac66eca475a42dbf6d8e2d63fc15ab1aff341943eb60fd239480ce52e7ff044fcc895a3e3d545a23b17b89029950bfc1a027e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87b043d5726422780ab3a7142d15155b4333f4297eebcf0f200ebd501c6fcd7182633e50b86b857d47593260c8db408883f9b643f14d1e7d2208e1e3b0429867aa5be49fa95a3d7ad26439db0cfeacd85a7efcfbe73e07916d35af815b570e441fb3d2ec1c142be1f1abdd6f1693476ab8698db075120e26e86f358a2538afef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8dcf21e9e37cff46a659375ef6698232d2274a5095086f92611f020d3ca87d221d512c084bac3e1d0e8edfe30cfd309dec8ff33849f9792435d6b98ab8fdbeb0fa89b12db000e4d4054cc2a177889bae3727baad025cf5935b20a3639ea1f8952fca093d98424ebdb21c65f0e03528b2deb20199c4be9df7c71612bc16920e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha48fdd9d2b7d13bd031d9312e8ca690650acae6c411a9f666cdfbe2fdd69421c434f550fc77c5d40d0eb06fffa988dfff6ea94d0f608a73e96277b87a28f90608efdd245d3c4432d62df791b72f3ccd71a9c96f5a64a230b01b2258f112d716ba359cd63c1e37c54003e2130bbfed47947f983f531edd1b7caa4e8466bb3e44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h992dcfdfe878822b3bfdcc0b15defb0a10f4892825860c721badb0f80e7f00e3ed21d2ee8d902dee7857614ed0edd2524806191d96a45cd04df5bcda6369a345af5d59035d7c209885e0c142992b0e462828000c6ad6ec5a14bb48732427ff5f60b42848a8af0d3ab1526ab74dc4adfeead036117f3b8a4f7f83f4073c7aaed0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8de0f73f0fc3dc129cd6d53e9be1b3ef7ebd64e034d0ee6b222f5804446cd0dcbeb2b570268089bff2677669056c996751b59d9c040256d639d198d694dd85ca10b262290bd15f91c0c5e5ab8169b795b7960ccac1697129f8cad444604d95d4abb4ff91a7eace7e3547f1889da827abc6fbb6cc3c556627dc1c06fa00172bf7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h466aa3d1338ed6c37775083c49a9af2ff904a5d06ddb327b36ba2d33b68887ea1b22aa5fd434629dfe14825eccb920897490cd77715155d786c0a0ec39be27c131fea212c075b5181db4c04bf384ee96497f926d33d3a74f545e2e825c527437f5ee2caa5555f8a8217df5ad2e86d20fd225d73d9fe48a9c56cea977e857eee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h766d04634beae6d0b41b11902218be5af8dba9af5fef9659f697c5380316a930812d753fbde6f69941e624becb1ca0fa6511c6efd0bb901e9cac4c32af35e91eda6d305f5c10482b494a0adbf98dd88ce7dfdfee4fbb1dfab32f90865ad0f875652b6d90da63924e47b923870968383a0b6e7088ec8f6319b50264151354cd09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf988255e61c8b7748aa92fd7176803b2a235b28c3e22cf6e906ac46337cd0a5dc98a98387b6fdc79629089f35c30bf433e73c2004a5a79ea83193fd3ef7a392ccf88cd95573a7ed39d407fadaf3ba6738fa838797ef77b85e7a1a208e581e4fcc52ebf998e139cb34650d9ee80e295406eb8bbd2aacdf1412c09d0490db37f58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac5ab423d20bf13ef356e1b53b09b2395dc0d73e06bc4953836c0c9a3cbb892d7a5d2e2be07041b516c4182db38786b11ef96127962c3fc09f5704ef7a3ce9e972747db9bd736ba49fc1329607d62d7d637383539912a56e9e683734637244c3b5925f0804559c35ca900f44151e9cbd257420b68746ef9d6abd6a2c189ed9b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he31b444ff4cb55ca57ee748f25cbff0d21db3abfc4aa3b38af9a58e3920ab17d9babaaaad3a241b8ffe8076761a0d481ecb52e40e6a89a6e9136625284b23a9a9965b4ab833de28dfc6f9a95a096481ae01067f9ec4d8c98f5635671a022e7372ad67bbd8dd6e576620c2c156463e1c997415c4470ba136faac96616863b0e3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbea2c22b4aeed541a37ac70ca8b354e80f2231f07333e4ca2ea3c51d15c1f6a48caaee632def155db1b830012d7b7021f519fd531b83c0db830228cfe6f918a3fedef657b94eeeadcdec7fe4b483794c0beb04436e04dcf6e3ae31da689d375cb49b859b49cf2e135425a60f7c3f9f99527819de3894b12709f8584eb262c77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h957d8b8c152adbafcb682ece69787c6f2b514bba1a4800364e8287f7cb522de4281913bf28c524d85dc3065008e6835f2fae5bb240f29bf7cf28d29047f004a49699dc177c41540caf0f63905d5bdd09c417484c7bc85213d6cb707169cfb4639696d4224c7f068db4c51ed1ca6f473398cb0dc98b098bddd4ff7d800645d1a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h253ec6bcdd51ff9252972d5cdfcd6ea8293ecb852cf8cb44e3b2e0cd18f99fb072e0ae7d8493519f7830222a10854492d24934324143a5d675b27226253f3ce2650245c99f59d7d04a5d8bfec0beda88e2ee90c711f57a3c0e3775341825b5420e34cc41a7c1fe63106003eb59d09d71570ac82f0faf88702781ec90744cc96e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5802060930399c6a3a8807841fb5b35c217cea8e3453bef6f427bc49de380b60fb45fa99a4049fbd945c478348d8f99710de88738fb02e098053aeee7918fd22738d1af08797baf028eb6dc6ed7d9f61a377079523f50675f5cd9ab48db980b0c0f26eea3d18bb1d2e675af72bb016b4996dfa196d68c40fa54bfab4998ee68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c94e255521af45f92ca136b74302998455bf6c3edb089b4209c8d5073abee0cceb6850757760bb68767d27a658ceddb1a301a20be0b40655221713791db3cf4accc2d1c8fe02fae27b401d2bdc1d51ab028495e4569d5ab2328f5a2f31940a4cc659179aa196a54fafe430a6c64806deee28f2d930fd97f2d23e25ea49510cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7fae314f950d08761d2731f97bf8550bdf0caa4259757355f41c9dc319cfd77a13c880d8072d306652ebc5c2a911f52f3bf54274ac2735abe6951e99f153c76dd8b399bbc2ba8675c86cd20e5cf2001abd446dd6f28d0b315cf2f255ff8a21cfb9bd81792c153eb3943d38beb89483a13871c61c16d2c142131da733108727e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd25942c19f766f4cf804d621355f3d3751a2f43f47ea87728a3c70b28ea77281399ba7219b328b6fb94cc20461bf6760b1c1cfc7f5fb798e082b11f2d922eaad888dd8c9341536c61c1a35d92bf83e5d9063855b19b31377860a5e28ae11e0ccab3c512e78d614c55f745066b678c8b5a17844aad2fc3136a33587ff3f421d05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15333a90673914b10d4397f4c28f34f1b91823d433ddada0d1c467cc52297f2bd2e3bc096f3fe5b91ad254ad004ecd8f86cd6cd3f8f044e2468a0925f80e24a4ff25eb86944f8981f7260e6c3b0fa0716e740d0fc7eef46201b51cabb79d63be0f0370bcd2502ea8d6e05858c6772039a698c2cc5f91cf470ca53d591336840c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50132c5f342520a9fe9bd807765a7642a45298b3ab0c9925532fc75344bf776fd62a8c3f389384b44e9240230154e67addd4945e593f8bfd10f5b8242ac4b43a17634baff518a907dea89a5faabb51469e6ddc9b66c56f7dcc605a5e57dec4130b7cc9000fd186c13b6b2c11bf06907c3ef74481d1c200ea69a72d30082698f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h459e2efd4e50b1a5d9119cfa56511bea674929e3fed9e6eb8b17df8d7ce458c83b32633596d9eabec53aa105c5d351ce4776808dd0db06c1b4fffef7cbad54c0db6e5d8797305fe48def52291451d50a6a3d666efa1b8acdc30bcb595b98da039106c5dd3a364372053ae61fa26a22e1bb0af7f86d2ac0756804fbed886668dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab1c69016c20b79f9ba75f39c2934adff2f9b85ebd68d39fe14f7a990dba64f2e75a3d7135667a0f731d42f8823b84041e775d81905d8f46bb272e4425a7299fe21fa100aac68926342a5963d9b4c99439b4173bc2e19042f3038c47bfd708c821c959b88d81c40c95b22b8de8ae4c559b1b3287c1c7b72a159eb7135cefa1b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6ea4d1ad50301727b49ff5a8bf9902db72065004e33b1be06189bca3b9ef361ceae73729080f8a8aca24dad0e3cbafe08ce1d3315b7b43b8ffbff2c4939c68567cef298f3b2fe73f22d03276b8c005995d40a8fa586ceb6bffb3062704f3cce8fe6abc9382c6ca3dc2929634a0d65365a9fd6b049da539bd2b09dc47e493aea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6c6e3349fdc1e4d4a46f29bdf0b16d896c5f39a3d59225c1ae1f4ec486574e9e49a4dad089b1834735c8b1f56070bcf57cc312db5261344c156a108486a58ac30c0074bd74f1322e069366fc6f25ca1d9c7834b0852ba9ffe2bf3c23ca0dd1a78b5ac1312a2284d01cfde29c7239c00a565f460d6facacb21a8a0d19c4a6924;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87db7c87224696014b921de0739369f7f137117c0f0c1215eca00fc930c119653ee8d4700d65afa75e8b3b6998050b3f698db9fc677909fc9bc29ab0167746e90f5936fdd843a2bd87ab8b71759270b8a80640c4e101b49df7ddf9a52f9a33469fe6c8fc3104adc82d99de0cbc5950aca7b310fb9e9e8199abfeec4a97c6dcd1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcea818e9afd2930ac445f33ec9cba0ef636f5b1c36b11c25650367838264edaf7133c8ec996cf1a82ac7a7b144c3ff48d1ddf74920a9993c153f29cc6c731e738a9aa9b9dc930def3cde77824106495f665a223b8ada69e758268fe9a73fc8b98c3be46bdf130c859a758a9daf3bde37585df204d9e4bfd8d54686079e031389;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h273b6176a2cbce59f5d9ba233f47299a0b6834e4fd4015a09c4efbb6f01bb718470b5a156da3be509acb8abf37994322fdf1f50d7b564ac0cdff8d6b250106d2e24d3ad8f850ef8c6df0948a65f35a20ffac85ad396a7b5f6255bdd1ee39e997ca0df20455e92a6c743dc8df158021a77ec8b8691d3c6e9910137d39a9145c07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfeadf3f0fc002924c1843b61afb4b8769af4605c2d12906d6e97ce9acbb5f4d126e4212df3c7181b56d0e183fae898fdfa4e601045fd05dd102352adf13f7cd49ee5ff795778528c268817253f7fc3077c4d37f05b03ff5bd892db863f1b239610e0d18dbc8b57d13c49fec6d0da99c318e0ea45ce8d7eea09e4c29b1779bc0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe34919738b60980909b399f85cd1dddade514210903008146e8584595ba1a66e8a42f7aba3e639f31db67d65840309b771e33b89c56d0ecc0592051dcfb042f731065e615ac8df9e981a3b5e72db03fdf02b61546a8627bd93bf7eaf159773f619e088283c659846863671f681288976e00d0ecda14cded815f3a4b55570575;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dea9d09602e9c3a99702e351053762f4d4bba984a1a0896b64431089960aeab79fa7cd140bfd55294e52bc74f3016f855f244736c2a2ed1493a202b7e1d9dcb64f2d9da77a173580c65fe19f596dfd4780491c78d6c3c51713eb7b19c6141b2e676ded87ae74d4ff39653dafc2b8b2a3b1d9db886ab4f12c8956723c3d7eca8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57734c94cf100804dd8d36fba8b456c00ad9eda99e44091eb304fc1508f9fb3d454ac7a341c0afdb75ae30d6de7529698c8018505eede30727b0a2954ebf9c5229eca88324bda3e6a167d43f76f5b586e80a0cbd06c6f343e5329e5703bfd85bc18ba4a4567ea5aaed11f3a0cb24004ebdec0a72d6190fba710fd3e7c367c3d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8b4eff883ff31c3a1700fc4d57778bff9470962918330f97247572a76038b0527ef1fae5ff40b91a1e79ebae5ce3b39822f02d0bfaf6b7db56dfbbeb56a86e887ba3befbd1f0fdcd6136e01d77719e6945cf8bc3f0b4022e53a971da882a81e053e4d0d67ab9347dd0ee06cb280a42195447e83863fceb5ed16a05c83a6f77e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fd8905204b8d8bca4805fb96451a9ddd99a393fb7ee2f08f40dfd8267d4ea337c2f4cb105b5745f580b9b7ec8873955b021907d05467f4e3c2483286f6a3962df56ced4aaad6bd180009363c7a4cb175ba98e467390b316b76717e484cd3577320e0f272d48f8a5967e57e2ff17a7b1cbfa0dde0f16fa85187aa3585ca185b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4751c6336c4d0662e2de81c5f69ce90d1523d18a608818b49c5735b02fc2c4e0ffae0b42e378419efdcad357b2a7ab94ea883861dba9c88bb3cf3626f573badedd4a9a4ae0262b54362d2c2cdfe271b3536381c1890feea77738d97fb6d76ff462ca8f30c5f63bf212e2734475917d92f809f203ffa7c2d4c6beddcde6c04425;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7b37d288287f65f9f9ac3112748b99f063f9d745bc3fd1fcf07d07cc6ceb09eace29289e3eb6bb4342ca27a841e0e5a49455ac4b9bf5db415e8cc77796928fecdd9e01d967240bad433a4ab16e0f236982fcbaf3da614e662e9ba51fb87defed9860212d7c26d6df7a4d30d702aefe62d6fa10da6f5166614ddc5a548dbee2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc395814051eb3430a0f7cb3a4fd8f832e9de2839106069ec083d481d0c7cef8778514a055dec498225e5caaf9cf2c58b404fba2793fe45ee5a53519babee26a4ba40bfd4744ba65d5b03113ee53e7ed411b62f5d8ad94e6733ce8074fc3eed39dc0dbe4338430ef89738e52b81a3ee62cc1ba7ceaa99a4811e0e31245822ec7f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41eee5abbda3534c62a7e53b9f907c7ec848ec76ecdd940a1fa5b3baeeed7d59ad42e6bb17efb940d4377c86527e7df03e4ed1eae6861b7be6d7dc9a7e1c139b4ea4a5fde0cc297d2f2e930ead53a915ff4ed787ee200d4c339f53a64b197d137e73335cef1372436d3f96fce4fd8f519cf1a8f543298ae370ba7934ee55b500;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc14808aef7d37ec4b63427e1e638e57f6448795502ffe17c7bc4265f9fe9dcf89c5cca6d3affa3fbeff97ca92eae3fbf245586abaae4cbbd4e8ba64f888a2d9a8ff8cc05b70f4393461ece7de0d80087c6f27427ae9799907f3d30193708becc31a36063d5db581658ec915be3ded7f9afe8890eef7efc29a811f2f021c126a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h236a1da10915dfe1caf1c6ec33c408d34b58d8d6687d867719eef5599442f7c3e1c36f27c3ea4a35d60caf015e061c61cb7b204fb0f5c8b26bf4bd15dbc9df63311d6e2d3f9f8ec9e99d4a89e980f10cf79c4fd488fa27d1e763e49c5b6158ac4923ea46fcce4914d06aca6a15b6edcff2e019f9ca31fea2d2c1d05ed4e78b5c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9305ccaab91396424c0ebe5000d4b4193ffb7c914a96aa0d55124156b9578466780c3fcae000e7e3d85635dcb84ac2a38439187df9b08ea797db082d21856ed3804676d1a12cbbbf6eaede0a52a65d429933d8cd978a1837e3de3d9bae14a7407356157e1e826a607285b39085c2c898f6fff321c595a50ee8b95a1d602beadf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfb4509aa1606588814ef9e882a2171fd551792c4cdf370fcc9a4ff7d06e00244c2f55f24787d6c0a6b92a23f12e722bee128e14d0a1407c02ddbb383e9091cf76764a98bba9bda3f70c364a22c04bed69155521ea479acbab0ec078f75183cf991a3c36fd4526e1f1ffe8e8bd1cb277a74f6c171660ff92a6da74f18e06883e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac50b18208a406801e08339ca1b7850e43e95d7d97373194759d3c2041d07e5ff53777e94717e82f67361f82f25a77bedb26ee029fbc022dfdd557250d6e440cf0e6be0b15672f06d8103cb1c6f0a1cfbedc0107761ddca2985e37c2f887fda1e41b5bc7c89ef55b6431bce00aa24e80e8be575118493f0a88baee7516304039;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc847906b01f4cd5fb4e1bd5668ecccc0c17903dcd74f10afad0ab385f912f84c4aa3fd6be93bbcc09071c45c30718e2bc41e254a90a306bb9b1dbf958a52dd0f4567474ca5ccb5ca23c22c48069e935f85278b4b70229f68a4ce8c602d5eb44c5d613e50eb8f813d53fbf7a9e2da5a8101d628485bec610037947482f8dfa0d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h757b3024d777790d4a03c2154958d94a1db8fef642f8ddcd757d9ec3dd02385a0c2f3e5275100f2051330e73b9ca36a3ada9c257351b60bf7fa89b8008b6cd21302f6e3e5050a219d4ccb5a09035218c335243febdf43adedbb87fcba57a8da64ee8479c7addc4a8d4008bad4ac5105aebf1211aa50f463bf69b14c823637133;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52147d51efe8dd450459d1238ad86ec8be9b9a00ec0c501d8fd21ca09b28caa981616308b89304b8615848d9422aa2fd6a5d87f54e2ce11e2a8aaa3a7bedd1dd73c81fcbb009bed5ca55e1220b6acd60df71993f3197bb7ed2cfa6eeb9db3477cf66bd1b3e9cce9397afcea0903cc3b40601f0ebacd2aebce8a78a6a84b7d65f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a98a86f31263a792469f70fc0d1627d08c07cb445e89d98d732371c29c37f753c0ea9c10cfbffc07d5edf2dcbd7622b2874d2a5afba30c79c66a5adc421cf5fe9ef3f0b4d85b6dd7f56ee878e507049cf1bdc2558df0f489292dc450fde1cadbed102860783956bbe2cc2806b4da2de7d251157c161caf14769f780c6e53e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc95c88b501232eb276116033bd572cacc1b0a93ad17df717cd2518b08ebd5111c64e4c3c00553b1f11783f153bd988ea2cb6d10c9cc2c6f339ce89a1036bf03a60f6aa7d6ae9fbc0bdca25e02cca596d480bb28b2adff64f775d8be9110f8401009b7f92128e293f4c527b80c0005009f0d2a8f27cc8d34b1e234a167436ece5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ea9253ded09d0d65baa644d9338619bbe9ff2d15c7412595eb29d79cb58cba47e8cf5c335f693931d21d4194cc07ffa9a20f64986356821ca45e549b0e7ced3ae15d33f6b1d5e5b41e62dfaec3fb8dba2da12330a56d7641ec458b42553432445c05ccec51c7b1e65965a22d0841dd247e9c5685f05c717d689b1e9e7b33a9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e34db2123c9289baffe815348a48321e98fe64539d652e07675d38d3e5833b418551673d1ce3656e222b8b2ea3347b124e21cf6fa97c41555cca332d658933c9711fc12ec1eb9fc37e60684bacb414b1a32c9cbda922d46fce1d0a400cd20d7dbc97c39ff4353ed1db4f4d7aa128783cf4c81b92fc3a88102aba60a33478d12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33052e970495975d860ef76058a1c5f3e64a584329cbcd40551955dbbbe98d6a9a3cc56ad27b6e41a9c34e259c3c89ce3c89c02cd2f37420ff580307f4afd3d8031ee3d2dcb9bf72cf4eda8da890e05b9a3c52e7f92742a7b4e51894f4168d322bcc0ca5a4158d8516b683aa2bba7c649203469548a1be402b8127fd95a26fce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d2703138e3af5284c967fcfcf3717efad5c0a87102aad51c7686c70c6e3645a23062bab57099ddf5249c00a7a575bf4aae5e82a2aa16f3b7105e78ce14b543719bc37cfa48f67ca11eb1faf505193017c44e793249284f3cff1a9a316af031ab80da571b78fc0ff93931e0e8c4e8dd53b0fb506f48d252e5de7452fc03787d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8de23322d2ae899fb259d330b713b8f734983c73b73ef5cdbeb5bd2a111c3606810207125e467187dbaa1919b6d153546bc779d77bf07749cf413c2117f050146fe6892000cfe87b2b95b5e5b9da266bd154f2f8ce61203465ef147553be2634d1dc7d3fee6b6d3c3d1e71206071f78b575c1c35fe6631e9a081b7afdd0edda;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf9a47ab9a6750f600647bfb04145e647464d141c5413f28d6789bcc1a19357ae5431c379e6361fa87a4671357694afc26416b9ec81507ae10bdb17c667e887974e3e6d96c2274310cb3f80d2baf974c702f4b977bfede18abbb1fcf1f8fc82f2ad4c53a4c23115a9b72ef29d703fb208d73bd137d53db06d0ac43fa51baa5b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1128d472d5f2c8133526bd795f45b0f8c2c8c2e5a33c94566828783f1739a52f0768f643f3761fcbc2597122a844833caaa879fbe028f91324ce1611580b62cf1770081a3fa7a4d5336ba677c8c0fbf22c4b407ce809b20e594181d33c0a54cc9e1e98e69fbcf14fff7a9e6d1aae742dfac51bbc1d8d109e1656b2cec7f34d0e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63e1ccbc59662b65bd825cf885b433cb5a238e45773b1067fac6217b11a52357572f330e690d714442fff5d89249fa40e100cb5ef912fef20844723c6917a1e42a6c2cb4ac3b1ac4cb2fb13e0e7a98aaafe0e74e695afcee385b8c5c38d63b37185c3b8ddbfe13facca14b6884da85b43c7ce783b250a0ff722a110652d02bfd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1630247a9515c3f43f3702c7ef5f85bb2afdcbd882c4e69b26cd57f2a5fd9d2e6779e2e2f7651a2f647bb63f6cad1c7b799a20cf0727a27dad17acef072e2dcebad840f07aaafdb45c3b75f567c76a0971a8db9428fa9d66d035c1c9f19e305439e6e1a7ed62f2ac9020372f59b9354daf6f80b58610292b40226d71bfc9a64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ba56792f374461fec0ac88eb1181ba7072710e5a2437976dcd65212c865c9b948d5dc65422b3de835827d2565b71c24c905075b3c7e6b4f2b278dc35a146c153f286f709b4819f2096afa32bfcd7ab5743bddab10a4c96bdd1c9d61e5daea70a9f708d786569f5d954e533bc7b9221b8d9b359b180bbdfd007b89c365bceb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71ae4b6edb22baea9791b5a635a341f5384d14f09a6bc00968fba67461b27c62d527671eb21052d18844504a5ff6c274a9e972b662e786945bd8065c8f8ed87b9e18f92812a0398d9e25049b6496b45f96ae0aa02605195322e5c0cac482848707a3ac00b4b8559a5ac7ec0750082dfce3b5908c0880548dd39e9a3f27f55636;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4969a52a6c4e457132b18c7f680e3ba6a65a930272d2fa15a4d7797635f368396b888c862180e2e9fc2d438cee85c8ddb794322f02c1f9717a6cd0c8fa5f014e7099ebecd44bbeff83fff3693ec9188777e173c1089efe110bd2fadae3693a464bd4a68802af5a2f3ef5d36a40266df2ef86db0a415631a67897aa3d13283788;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dd183b72a8c20d913aa7572c1e1d59600f8897f50d444bf412737ba6d787a942d8fe5b9bcd4f250828aa618e2c2d3af0a5046f85baecfdb9fab6fd5ba8f85035e764f3118b499b54cae58967a5ae6395d20aacfee67437ea1828a18e8c1af9bfafeb26de42d47481ee083783938f63cb347563b5584f256888db5a51f05b26f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf120e25e9c0afca89bc907722a06b0712705ebaac538dbcd8a0c9bec3ce65ef1ae4b1b86d88919ef2428c8ca33a214dda57cb3b3f4166841696bfd69adbf2a8ea98ff773ef9639b83997c343887f0b8e86ada61f6af6bda49c0e1502fbff5e27f82d0137e4a677e8a7712e974ed4a4d420971649ac9b40e6f426d8120249487;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5cbe67b45a5c78dfc894cb7f80de747e3f36130d5ea8e9b2108479407ff6e62c7402f5d82b18e353b9729d2d7d68c116ab2f35ddc7d480112860571d3ef476151364824a1ef7bf4614aa1a64ba9d5810565aa3207ab1a1904bebb6c988a612c09583edb284f3b01917319705d1d630b9faff050f7820542cc008b55a34d8843;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a88a8715227249ccecb4853b26ccd8f037b36810777ff85228fd54a9111a33797324095116d4c2864c1aa54e07d902d3bd0734a634018614ec44d288bef68dbee555ea1046f570464b655380395f9dee130f7e613f0ed90c514350cf72a0df48c07a5644ab7efd79e5ef093e47c1c62a5ab6e2d6f2d521da2b5449b8edd7383;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11ae118da7594037b7a8f62e408fed2893eb669d7c280945bae918caee9bd27a94d28299c6806cf0090a2d6f3f40c22e3a84f3f00b634d9240bd5fca656f8eebf9c17cab06b4672433a00c2607f75fca495531f6f2922bd97a89b8a73df4adbb211081c07357eb5ec4d434bb6e6b1736a56511dd7353acfe403a7463fb516772;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e5c70575eec18e1a6558684fe43135124d88f4f9866102328427e8c5cf81fb982ed185e6429e48869d5507cf1d91c7cc316bbd3ec21431c364ffe027ef93da00b2c87c3e87d88a9966657afa8581fc794b76d4a44d5f220dd1be35399a88713e2d6112cb09c384037fd084356d927db269a1e33f8c528da9f14475ed0d0516f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5964fe3d6d658d84323ff80421e5bc0c29413b0846c3ba7d0b6ba19a949db274513fb7a12c09d79a021013c83c19bbf25efb3b459d62654160afa6a28381771f099037f5bd1f1ce9e0504658e3ae6b07271a2a25e02419c4c0e8a926aaa70ce601bdb88067119908a697205c29a229457d4437c0ddc4db51d76de74d38074a03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7260c3da0552d870c41272be7522c33accf3131294e8786104bdd1c373b499ddf5ed1be7e7a633f1c6f65ddc30cd95ea81dc69c71faeaf56c75c99e5f458d9c242839ac7741a3b29f805624d4d331dc30171c7762348b96c3147952c95905034e0d2669bbf43258e683526275f6c3f3e7e34d29bdb482ac8f05b1d3c1c92a18e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd0bc2dc84aea3415b41a40711a3c833ba949fddba468b970bc13424921b6d1f5ced2176146a047674ab74350e33e062b3fff5064c5e42c85f864993a3767cd5a3c94bbb919cdac8f72ea99bbee72e79a5a3a61441aeb398592ade1ac8693ccc4345cbbd0bd8580b39bff74497d14d792c7ca4bb2a3576147f1efd9d7118e1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba16d25988bb9cc43ea24805b9bb277bc33ef29908bcda82f2aff814f96ffc160fe36f7795f8baa04e940436e01c1148e6c118d8e88ad4c627b677bfbcf79ae1ead63ac50ec0ad8072da988fa44f59d1c3399d4cf33c2a342bf3669cf0ea270ac1300d190531b15da4f40bd25e589d6a21c890e8c1e1383a512419404ccbdc05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h733af1523ba4915b1ff653006fd1a43424dc7d2383e78477247c9f35dddd955f307e487fa2362d4d7a59f3702413b2b6825cc7d04a49879943411dc4167657e23ca1fd94a329b125e19275c128cf08fdb79e7dff36c70c5aac4270cad20568295ddde1d22528d1ddd0df692233f54ef5a9bfa48a5592095189da9869201e010c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44d97a7f38951919fabb0a3a2899756dd749a020d2eecbc2cee82d0c4b0bb4a7c098349b8951845b05aacbcdca590d6183a73db50f7571bbd8edd21de82d329a6ba31146671950d1cae9fb71005fde055bd3aa3b1cf26b08f2affa0ee2711856b2a8a77d3b0cfd4c83005d649be48def885a92c9e85ae077001c6c5ef2d03723;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc4f6e152f861fe075b78620052fa054d1a74f1521b5ffdc4f29a287e545665272b4c65641e25fda243efcd883bee8f772f4cb785e595fe6468fa9be4a4371bb9b444780415a5c0c35152b5d1713faab1c09df6d63db0fd6414e5ebc9263b60b254c561e19042a1cf84f82e4205541226ef0c222091aada500d6a2eb37d62003;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cf2200aa8bb614caff1c9bdf2a8251a1e23a2c1aca24ec7bdd7ee31701e33faa1b2b910cf8ca5bfc12bda59fe02d8458f09184ca40292dde971c79f9d54e51d3b167fb12a2b2de9836053a8db0a6cd1242ce893560150141c93299e6b0e0cf1297807fd5c43f2300dbd13843a7ecaca1ff9245033cdc0012c07e462a2834b34;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5628cfb03b9d97585bcc851b4dd8932aee9507e07ef6358f0630c4a3074165971c3ff1767eb3acbe4e729fa3abac4a03c46fa0b9fc57cdde8c3b794245692536c6bc4caefabf75d054b5adfdbf097e0eb45bc49afa985dd5750a0d8b24b9486e4dca425464bc415e5fdd01c5e8c6a4fb77e2eb4c1117ce5a754677117df2c0e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedcaea817c2d711e7a0591f69775c10071f0418bac78acfe4f790c0726fbb87c10ccef2afdecd37a43cd7f3d5bc9bd95a04573034bd2011e4e621ffabe56a1d2735a74a49809088d31cd00c5a1d055832dbf375e8db925df8c52ce5ad8ea0ac82e723b076ce19859252c3e778b42720e109697ec6d1c1824fc26bf88f87c4d63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4827d476137de6e04d85de69f5902ac566c62985afa6348fe07859d646e857df4a9c703ee25f4b8082abc50ebae81b99906583dc91e8a1940e37aefc3738f7e59b677ba1976468e591c59621e4f6ac2923a837339bb34fa8472619f736f2776c3f649e87e3e06e7e971562a4797efb624c4e5ca0cd0a3b306c3daa0da182ccc8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c8ee6dbfb4b19b1c24a6a911a581e5d2eb00bbbcfa15d18968b5ff72d50b414dd0cded4f60fd748cb17f7be2ce02a5dd77112ee014e424ade4506bb896a5d33035ea6c8cec5043b54b1b076b775a8ff91aca9ec2368c0275ae60fa693e72d24397b919a6af86a7585106b49d1da4cec8de2084cdd2d42c40e7250ab55ebdc1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h839485cbd55728adc96b4abf65f3c5f06e9cd17ef9dcbc283cab9d2433909ef77bebef19b3e39fcd2581dfc878b866ebc7cdd8bc2c900ff938643b96a3b9ff79b221e0ff5a8030f6eb165112feb3177d0397a3ad3700f3d1df319f4d96a8e2c467d985ca9e28a70d0f1868e9d6d4ce66a0d18a28ba8a8d45b8756dfb2d938ba0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0c1e7ee4a4a23cfea371f2ff0b33730262e150ce5f144f64811e43f78441db2f8c0d2d22829c618a6d56e1d74551dbaf9e6b7c207ab90f908f2fc502be99efc00574ed33dd2608ba93b7c5a69d7edba3eb04a556bcbb028df4b16bb4132d913d10f661ef35ded1313517b5c21e59e73b37f69be04521eff96071a70bb19922;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c3dd2b9db7a67854bec9b9792ca05818a1bdc928404c49f525c91208bf6cc7b1e8d10d78151d4b996ad94b8f8b871861bae887c761baab9a865fb6c1b4ee8118fa153d38bfbdf05bdcb9cf48f034ae0ae9d2d5607616e5fb4c230a5a2025a533ff12be0f11df6e5d1e49b6c7843046cfbe4207d22fec486e32160c1998cdcf8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdda766af0efb115fde9e4d3bd4cf73cdb677c8c8850cc0be5b3d26cfba56f93b2940bc3efdef873e8a1faf40b6f3adc7ae6dcd12afd633f932867000a8abc97445ba38bbf93209af45d50e8557c53fd9807c6a578806d4c0cf9f2298f1a452c2fe8e7d83e486cac62228fb8727afa0d3a7ff73591f274f052db316b3a24f4002;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d7a1110d989f6ec0ac298fd4eb0d6558db2ea6475dab05f854f04093613492825ab96f0d3f379a69657527334c7c99501963516e34933ae7b68977f12dba7eaa607ca7491ed18db3ee7bc0ed98c946170afafbae7e2fa3ceae2e39a9ac22f7e97ce2ec347118bd4d1f2eb9d320405ba272c28f06f289beffbe0c46b90990674;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4307414f6c5e2f1ec8fdecb6f4f0726b8fb26d0af3bc8f826d7b9464776171b1565483f03ff74312ad4c48db82bbc36310f0174ccb69f835771eb8748cd5659dd46989c6b86b42ec176da01cbab313812a132bd27c870be6e7a0107898de78826766f4032506b56f9f430e1b4450161888c69505513b9e8b698b912fd6840bab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h888c188fcd40afa375316d1d453cdaee0616925b4c3e21564d1d906a370f862d779dddefb3cebc9085ecdc9941ae5da99fd214806dcd7fca74d737bc634a918b1622d60ec1ddd191c24f58a7b08b1e989a7aef96784556f0089fbb7ce451c523c622ee15990f82d51cd84fe51b57fa20b87ae6f896314bbcf9ab15dbc5f64ed6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78fc53eae4965bb73147a11e71feae32926976d7f1253d0c290707a958c3ec29600eb7eca3575e680373fe60093f3478e7f3c26f811c88952fc42ec12ff052ff0ef8f3cba9a5760470a65772a32d8c58223fa8a4262e725b42cd534260382e3660a1361ef59ce2291c146256f0ed9263f6aa3293e2db5fe859f515675b1a317b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16d31c16022a9e94eabe39d2d26cc3fdff5bbdede523e630128502a035b65e9f6020a66cd54a0d47b1b92b3e96eb46732a1278a3b9bd526ccebc1b1326da8389fd9b26464f42dc735ae3b657507dc00a8933e85fb571baef9e59047c68fe784aea19c99a73247130c19ba5f03a8a81b968d79c447f955e2749c03ffd48c4d8b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59e460ab8ce89cf494da6e8f12147be77b7df49e0b5850a4876f5d677e4be7bc840185f47a7baf3f3917f2322291064bfc3093589d94dca1fb63596a35adb0c3f687655ff8bbea6ee69e5de461fc04c211a809ed4ecc2d3caaf6c8e89180878a3aee50aafc0cabfe2dcbfc1740ba6e01fb6ae4c6b4193321c105d8db97f2bea8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5af1d47f3d335d50dfc085f49c85aae3a955fbc49e47d73aa397136afd2d36f05a1e75c617a0e5ed3493cca6983df5a9dffc4b25e76c439ac0925cc1a54a388ed6ea91afba1f18e6d0f863fba5ac7dbb06b607bc482aa93909148325abd9321599493b3e44c48e84a1e7d28fdea67c049f825eadd290adf676cbd264a37a5235;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccce3cf5bc7572011d11bd65bdf6624e5e4a9c3072fb56e62a57c13e2342e5cca6d87b1f36b6eb040b802130c6c02c7d532e5c8a2c9e27baf886b369d45264efb0c8f32c6b9d8efd1b70df9fb89abecc9a4498dbb32cf8190455febe087e5032998af0ef6eeceb342bc5d0c22894b917c3020b247c3377cc7fb08b431bef115a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9a5facd1d6124b305557bd566398e008e181056ce0ea0f833d867700b183821bf361d760c8add755751260667f71c1e7d88c0835b7b0ef29cee2b854510004e2b5e3783e176ca5afa039207321928dbf0311f0033c79ec7eef1a0a255a9ca3a4c489d638583805d2670e9c0f1306924d7a05adbd9fb08805a73f4eb0c2446d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14f0e6a14286a3cf1f45d9b3873e390e2d46c86b05a821b183480b4879328ad8e791ad54958c3fa6a6c7348e13c8fdb2c89f1be1788eac307d8a6f0612709cd119bddb41464983bafd963975c3439b9ed2ac7fddb7b3dad73c2fa2763ccd5e33fcef82423ada0f2cb9dc2d851a608b48e4ee0f39024967dfb61fe04420e99146;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52938a6400820ae0d441296e90c1002a013e5d25443903fa3fe0ccee1a0697163720c17cf382c8f87c906a22183977b131006d3f38a176ad22b36265d3703beb05cf51c1d2057a1e742ba84f0ee37633267b77529ce583a3547d39e376ea1547507008cda56d1e51a9d8b5c154791ec1b55de659210dd8cb18a1dac3d7418fce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'head833aa8ffbe2ec3fe8e193bb66782408018e7fec9d55c8c478bef2fdcb560286ceede52f81ac6a85747d0162075be784c708925f33b757eddff56b2b12a0759f5940366ddfe5778324ae6cf4afccc4e5a8f9950d25bc31233495a9af06ddae93337a01ffd91e88ab15601981c5cbdf85d22a513b744a670980b017fb423168;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc867094115c3c7c03bedaeaf96c9eb1d8b85f52aeb60db0f8b46a5923b2deed36c07311d5fbccf11fb6868df9b6e0e384a67662d97934fd0ececf53c5df5b85c8b649aec2acbd3f48a43c7f0a1fc55974af2129893ee3fa0122ebb81f86df5c1b92b41b8d1ab7f619f9622f5bb15795745f653c3151f265faec618ea055c6fbd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99694c5e03dca187fde723e3dbcb7f243a124dca559e7ab1c76d4e0b7f081cd2ccc1ebaa6cee9e1e7d21e2136bdc19fd117baa0afb3e6ed14963ef5de68692572477d510345ae31275b7bfee75c36fb15f279f3f36ad21a490a3fa172c04453177b0bf4b8b875d48b3561f55b79795b23ace21921adc04dc6eb15a175ea44d0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5462e5209a4b1b95b3447f0c5225f7a60bef5136e1bbd7b103f1403b1e640d11f116d23ee75fb26e1a9f801771db640e28c9dbb7176b9489a3dd17ae66c9fc7998f373360135418c455f90c2edfc4d8d107bb949c9fa588cdf41d82d713db4c6c1750c5475067b47ec1d770b143c59cb04291f7ef07484a260a8e31933c8d680;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24ca9d478dc78d8f17b82c52f1902234cb6b24fd9ca7c0ee089bfd2232e632eb9d6ad94f647a18b35ab035805dfe5d5e99d4205f5c2644ed9ad4b1ab623d9a432794eca4f22afb551b674d931b01063db815f76c8102df7b28ea85956b0b0f27f10b1cb25cbb8fd6a3444e8dbaaa45ec27b9ce01f0bdccaba43cdc6e691d493d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2223eae1224c6a294d140457651af714900e7c6c1bf8eb68f4584623c32a8b290baf3e041a057bf0d7325155a68fc7a37fcac7501bba3622a6cef2ff0113c6e3947b7119597ca6e5f36fa1477cf68b62d158ca20b113233687e37be116aee364f6b7b1c4c69c4835248df2dc13257264a611a35a91991ebd587ca8ac20e467b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2a87967c5d150e71134d42893486f187d03e445ec7790ff0b3113324d171fa50acba214204d48adbf9b8f38842df5c8c179db0b2d27041ff763cd08ea65e50cc68980a9ab894b3b181181c20eddaf4bca4e0564ac3bdcf609152afc699876f34aaff0f5e0d3d817984b9db26eb56d1cb8c8aa7d5ce7ce2273d196dcd62dd15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce5f11c1b8a66e138d39374fa741b36b62694b88a566ffd0b0f68ab09287589ebb878534d0506ae72108e5902172315a8bdd38d1729cec0a53f422ecf89819f81bdcc312661c4e9348abee9e498b56dda6e856bf329783e9191a4efb90f6f7730e33f17e25bfe83d643941e63383a43f0c215507e4bef3e7810e78df6f1a521b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed089da31bae7bc6e96239c527d61158c06a5178db02632cecc2c7c90b1a9ba8669380cf166267ee51faff01fe51732a1eb66c4abba6f68813d44fa988a3aea51c6f33d2c444d006796e8367061fa6fa26a48e923a9e0d198d7874bc00a9d0c1e00d5460d03ca842645e2fff8882e1b52d914c3a9779345beb313e60001c9bdc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33b4f4d0533ec91488bfdc1a1b552d92f2d5af057813380cef053ccfa9601a1adb684a39f5e75b0481f96b6a582b58d4693be7ba3e74939ae603f5ec7a72e0662102ab6efbafe0907dea3330dca9b77c309d5bd367cd07ee561d627fc13623b8daecf9f3554108a235dbd4764d4fc276a8e79892fe10ddf5bc9b3d94cc489440;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73cb77bf65ccf2a1089427d36f19f53329d909d8e7e65b744ec4f312c0b017179cce87084840fb2be315e7f4d1b1358c94ec2ac57677a987091950c90a59c036297e379e169e9debce92c9daac8f45ab1549230b53efb01cce20a91ce9b42a1578ce4d37ebb1778a3e4bfe75d74feed503e9fb26ba05335e131f82418f9cb2eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92090a1db11b19ada22706bc0424e04417f85dc0e469b5197042bd5abb7edeeefc81ac806375e73c8a546adc9499c9310e6bb9893e17ba0e081c20b39dc87a89c7b5b624d43936a6ea4bb0ba2d71a96379bb62a1a2c974a73c603bdc2c7bf3de4ee9feb81ff1bb7aefb7d1467a403a840cfe348bf61332648e5af074be3855f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7cec15fc4b9922eefc022370478cf969d7d23d90da66f9e46e3b17daf4d31943199af84f4276cdd1509442a3634fcd559ebb708c7150c192da1305c6cf5366a3d4a72e3602912f2e8374f4f0673bf9068eeb6ad2d34f6f7aa5604c8eae067173d497fdb1938ffdf9d7e09ee5a432a8ddc7279a2fb5aa2bc94c9dc71cd3d5a78;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c0ecf5030a8e7c1e6cf7203c164871336dfb404caa09e3329fe6e77e2ccf083baa246e7b1b971981bb5ea5c3413d5fe90f82b7625e8090b8e5c53add2f18251c5b210894e295b0055533b3688ea50915a867e7f85fa000514ecb22ac42f106acd1c190c7cee57d3513ba14d38c38a7b6751bdf3a77f2c5b2b7643b30c719b27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaf4e9c176d7eed669e1b8cc2d5da6b447149867fb24b7496411fd8652388ba639ad6f5445281238dd7bf11fbff476b81e2dbf86d43b45d3cad7ce6fb95653970a8f178590cdf9af1563fd2b6ee05a3b161971da7ac9e2a843772e96670dd2206728db28731570bd960f88b2f043f168f765c87adbf2e6cc38b950d4ab9828c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hada465672dd6e06bd7541b664217e4a0179765795f36f99f2b21cf5fcaa7c11c176e5092615687454eb227749bccaffcd1362b07732968e1662cf6ee247983dbc1f22e49361ad8af37ebb0f54ccc3b36c2ba32df3719ac4edc4ca5b6900d00375e0797e53ea2fec712d93475af8b4760fdbc56977a356d0610d1c6879d1cdf00;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1391ff0922a9ac536be1d576d12e662e4fe0e3694ffbad232c065dcf999c5e0f8eb132dd038aaa172b5f2f814785dbded93ac752cf2ba0e6b1245b2d015ed346cb53023ea1eee988d37d334daea5ec6db3beda9d00cb7e17488819e7a0fde9dc0135ce60e6ecca7157b667b5a36e17d389a0ac95d01895de90f87ff99fe8a9f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had6ee2cb24ddee3dbb7a4d7d799b2e1160cfc97bc3c273fdcd3b04e2d870256378370a7d73ba75f26c56ddcfcab26a605be02cbf91692139b3cfcc3ee380c47179c6fc5e2c0780ff918a91d7c6968b01b168a576e64049de985e602c12be8178ab59a97b05015b191d31f207c78807f3a64556888482692bee43815c5173423c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7e0171757f9de03bcb1738c1be23b77e8f062ef4ed4158484a8384235140ab763fc34856987c130133bba3e8ec91f5e59428b73da0e1f9c426834f7a66b30238128031daba2085ed3df3064b00c95bb11cd228bc7fb1a94ad9e8f59f8c5540ce3002020a1758b328c14e157acc3d8890c24c6f673108bd11242cbc642a8d242;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf61e429be2a6dc377d1204d7144e85921d36fadc22636f6e3bd302438b3cd26a6ad2a790ed312f2cf8abfc8d36f00dafa6b5bd77275e3944f86c300aa6c7facfd1450fac5a83a9a250fabb07499a325208c585e5eb9762b6b7cd0d1364ac40ff0989334b0f14bf5ee9fa2b39d6c2c20947c9b6b4808b98c3f7b6c766e347186d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8aea8d0474317141f807b98c58ec0fe11d9296b44c6f56a5bcc5e35942b881cd33c573148450f78e4bf500950fa21468b69f75cce8a29f46d43f589f043cfb2fd74846940fd141cd12bd13192413af97f7d26e024ddd48b8825bc8351d543d87e94ea58b2a210f4b2e3ae6056473d1337fcb6456f06d6abe6410facf1961a159;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9406b4bbe752abcc2c6fd5bd485bbe29f018227d3bcd587c86022ae3fd9f16cdc2dd5f54964ad98000a21ace038fb202bf0c4f87eba41f623e83438933ea77c610ac4800c89cd1d762f3294c29c64dc46cb255ffaccffaeeddeb4636fcaf92cf71bbeba796b52744b727617714f9e47ab44d819a637c538207e0a432e8015a7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27cce7a7622fbb283b96f702199bdc836824e2602f77dcd92f3a480416c3582aad65faf1b39b1675f70d8b515b021e029b748c1eb915556cc1e1b5cf8a076e3d4cd8610b7c4a753f821589dd8bbf06485b8d8d12e3505615847c05b6ddd493ca8d4e02e759002c871a47482346fd14d5a188117dac49b69db8a6de6673cceda5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2aed6a7d7da03c1bdc4471d1e5258c9bc98fe02f900f50a896981518bd871a6dc4c412802a116fde99bc5194afd6718b19ee8240f2508ecc6b7869366f81ad00f6214837fb34026a3544d6ba50d69640a9dec96a696ada9392285202dcb696f2bbd9985d757c27746d7a0d25b1680d66078e1c816acf1d58d0a5ca12000b7b8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb29fcda1283bf68437459b2b6704d9314a4a3e30423022313d66b4f11d8c0391f21653d041a007ba3adce3e606a13a0537a0ad22cce38db71ab5212efadd4e50ca433cd6d7c3b48219887df0c545d2434cb679d8a96929ab9f2c6b272c5689fbdb1a7db5c45eff5dc0cb293fe4ea03529a18c24c6e720701eae9945a0aebe02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h758ebd9c5cec6147befa048c8f20b070fabe113c082d40457551b2638fc099712a5e32a000f21077c75bf6a2a41f89a9c5b4be6160ff73241e85b33e7c96324025d0f6e9b55f73ae8f903dbeaa6fd7f41facdd2f38d62c813950d18f49bc687de22ad58e554f22b96cdf58c8627177295d8c459e37af4aa640b15cb2d3bd6365;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67949ffa7048d85f12add36e74c9633cee00140dd15b642d6216dcb198d509daded08b7d7d6894d6ead2be201cbd2000ebdbdaf5797caccd817c88cda507418031a23181bbc1dfa4f756be84a0b184033d6840d61467e2ac171c77e35ed523c0a202cb272c7073fe37c1894559596360e587f7d489d94cb801b8ee25cc594f04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebb73a5d9430132e1db02c1b42d368a2165f55b9b95d751fdf57063e4e379ada2116299748200806998c6c15420e436a6145ed454430bb0541acbedeb7f7d630acf548dee848107169cc3032ecef4f4d16eaa591591fb14b323167015ebc8305dcfcbf73fbb948e8a948dee7f8ea0750bf2dbb3f139342f0dda564cdcc1e337b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he237089b13e169436735fd87943cfe3701267d9e978a1cac728cc98cc548c414cc367a0661ffd52f0fd0e7d51f57b28853eb619dbe82bceddf21398ee9461522e6e30c10ca1ac8ae6714a1bcacaca5538329d09051487e0d8dc4425d66145aae5fb4cba8a3930032272c4975eebc166b6cf2b616b81e59279428d9f9902c5978;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd598a39c7b1cbaf462e085f3a44b1265a0b367c572f7eda77670b42876b72331f67cfbaddcf7ba2ca4017803fe7b6027c787ef64d7966a638036a304afe935ddc1392bb7b3474cfd1c34615a9a2dabb794b267db37b3de49cd2c1e03a2aa024c9ea8a915a343f64361af3b21b9ffa8cd47841240783ffbc46f8fbb50a83c5d24;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9288e4e27ba97b653e434aede3eee12826721365eb5c924c0d5fa6e0fc1ff3cb2ae56a235c9aa5234459675300e2c771aadf117b52a30f996a1c72104f1d5d0712535c269a3405ccede12562f15867047ee4a73da89578322d10f7ad8f0a792677c1aed2079308eb60b94991a75472044f32983a3ed1465c72e73375a941900;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25f4c06e2980c56a6c1ae318f19860b6f9a57931e3427cf2368a22a02cbeacb01c06f40a8ea5e99bcc91d6d5fed6025066381667ebf41540cb78de0aa3f521f748ef64f22c522da4b3faf299ca51e2732a9182990d7963eab83bd822cffb3daa1591847957c131f622e9e9fb55ed79c7ffc90a7083d3b9d35bfbe1246f04c472;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a4e919e269990f360951140a259f1d8386e6c8198ef89081a37dd80fb1267a9736f088173c0387319b5b3aa0f2f959803a4a1eff09c6ae907c1610632756b95e8bd8a9a25b076b1fb8eca04f7534d47439c675a2079eb62317773f9f4d9d2d379bdfab5398d8e4f02b0a47c86843fddb1eed9edfac5915dce1a99a319433046;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1dedb0adf3003b7a4a4a6ae3a3af55a72f78fd86a55d0194eecbbfb30545a560d38e4d835a99e625cff98013a8e53a34b10e0661fb0c73e23b1d5a329144716762d182bbf777778966892150e4e377f0730ba3126d7b62ae4fcf4277a34e212a81252e52251fc74b340ab7009f1e787149749024a659ec883958f3132167ba9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9aa4f4953c9b89aa6d6704e0f4d3a24257c821f82eb712107afb0fb8a5fd478c3951cbd6970c67c843f331c6f23959009ac13026ec6b1eff400cbdd23e768510907647197d544f2ad1f3c5a92c7a8bc7cb2eff1594894c05977e14aa4f3848d4c41d538af0f6e4afb0abb9e8e3f457b5149f86d45649bc589bd043823381f127;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h610cb000ac2502e3ae6a0380d596a986ae5c0f8c5653777a9c74573da7e164efdd38c6bab814563b7810bf122f33ffb457ab4adb19a264ed185205cf9682a4515f06162e5b2b588317a48748d1cf5e37211b8ab483b13397afaf2b59b0e22ace28073eab7c50df364a9e7425c457599f209995e9177731e047640319b28eb305;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e9b5e8245008e68de89d4a47c365d15424cd621b66d47b900265075ac4a02c90348e40842a00f3ce77f8dc073f018914000e0c8ec61277eaa3af4babf6e9516bac25c79d3b26626d0ce8b4aeead3351824aaaa922a9c44b0e9f39a43f102d6904492acd35a7d24f958961eb70c61f14898c247275d27e2df0b5b18b0a83e646;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he00e22c71581dabf5343a16f568a581a90aad2b42a4c96c5676cb97cffabf9fc077381bcf2f63b1828f28671db0fb6ef08be0e51c7c8642b0a668ca8d04444a917e045221770afbc2575a98491c5b5cae20032a0f35a1f19d99b70b00275d90a885d0fcc2c650cc024d1b2a9e021082cac8c24e568b0b53e2ceba76ae349440c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38740a3f3c9311e25be6a727b490328d633dcc19ae95588cfddd0ec53dd7fb0fbbaf8e425309ab41dd3d533f84b61163042a5ec79fba0fc60846db4b649816bc120a62a793eb4efcd7c0044ace8e850ced1c1bfa4492736c3e704837dc97524308f9cee91c89891adeb5a099a0e89049e3ded5f2f73b12180a5c3fa992ef5bf9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h987b058ba4ba20929ab7d6540f6b2e1eeb92d0952e3442bd78706ffc6d6753bcde09d03bf07950f386eac2ddc70a0c2d5ddf585920cb9a63a238c24585733c14b42b58e807ee6828bf4142562a32c035be80983360f5957b46fd2e04626d562ff71d30f7bb4d490b62b80c27033699e762c4cbd85b1cb9734a8b5a2045506b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74e05a9576b9b89e4ed6ce6a37904b53ea6fd740c927a0f52cf30ae9b26765fb85f372271b4f79f94294675df26d9f3cdea9ddbb62cce9bea86759a2c2ab4d9436b5c9203a1048cbc5cac9509b02db44b8713adfb5bdbb9fa5bc9c492e7427c7de12f36406d2e76e772c2f6f7df922b26e67ec1f54c8706b4f7453116093a0fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f1ddabb9cb676125e42756af175d88f99da13bed9abe59dcd88f9dd50217c3ef4afa75247c2eb70adc48d4f5fa3a4950ee9b60ba05de28175d8e63050254f9f18979a6717cd8ad9041e41362c6034d9c1cfc348de0bd996a718cb1bf220d8b9b3f342a395cde3aeb9c3821dcf37a927d9f65db5ba6e4f52a1fa966a053a0e26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52b252488fe9b2f9c029769d62e1411f80e1994fb3b63dee140c8a5663d5f4aa2d2e31b45b65ed3773a6ee1d4615e971d2d79148b1507b8ef58f3bd4744cb88aaff1f5a66fdfe4f85bca3171603904517142d2d704a0f9c6bf4a50293f2e98893e44abf611a0b40fea15052ca2d42145502d47ecabc4ee654d64a59bb297898f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b34b82cea990d43af1eda3b39bba4e42961559067561836524aadda933f174ca44d3da631c860ebf1f51facf22a501141d675ba869bbae34bac4651413a97cfa74970d97f42f43e54aa227ab963ece7d887d96df544dd0422419480a9554f9d407c8cca3a8ae3f4dd0ac0151dba39b0d4f7597080ed1e0a4f1d869bba75ba5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bfd5817122f187524a074d6cc59632408ebb4180ec21f6ad487150c4ac7e9216eb4e3bb4539ede2d24bb9817765014dd8172eba94509df6390ff298c099b921b21ad794ec7405befbe2c0b8091659b69fe6366ef268c532ffd4a46442c884f675827f3dfc2bd00dbb33987161039aa8981ff143da3d1943def7b6380b23f873;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6a194e987c12d877285733b2cc482e94ef22d1ce1dc4934b60661f410f7d5f2f753573e3f75dfaf44f87f9af5ce2b9189e420aeabdc8ade0dbf8a2a179a0fc0a77822593c4e80aebf890a192a0f8d0279e9ec991442922016d330039c6d99d5134a57b7e24a040060cab7cde79477da4782226cc2e1a63da841c0b16a374df4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d548fbdb2b7e03887eb2c62720ce7ed20467c0b88ad7f018fa137f420fef0590a76d98845d98ba40ad86432dba6cf52069f7a354c49d74b31fcbe3dc06d9b43898d98fd197dc2ef6b161f937fec8ba50430ddf8200c869bd02305a7aa433f62b1811e0f154af0022e7ae91659b125f860988baf4b7e8df181242497f76aa54f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63ac2302adf53fb5d0e129ee063e65631538b0035f9f89d40d587ab41b54992208810f6a91fec55b51c7bd7b295d54fbbe782fba0539bc3ff368352623da42a8d0fc421efbcd09ba00f1c637c6c0036979d15fe24f7adf14ce88c7b5247e99bd1077180b0bb418dfcfce0bdf2f433f30afea1b3643f5b38f66e94f2b2bee72d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf36f9f01c76249429779579d58f2f198a34c564a0673b308fba37c1d383115090abe36adb40958dca5949149b27fcea4f2048e7fd12cae71fd7affc2b55c32129dd58e4d161c6cf3e06a8972d5a05c03486bd686fe6004a63b155f635789c0f4d542daade39b8ef2c404baea45ff44824e61b356d4bf17e8ecbd124a1801fd8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6406946251ebf8c4e2b126564f9cb9355e4aeace7a42816e3fb262d9f00999c9c06e8d5e4a5d0bf536b46c2f5436eed5931dcee0acf47b99c8f9c41e2848bdab7caca0ca395bba6c3f0170c164b4655cad4edf9316d1150f9b2671c1f12f32d332df8e56659a111a315448fb927635e301c2f4982e9a5ec46035660be265799;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea3ac69f9b4daa5e1430d38cedb23bc246e6a93b802fa042853e3b897ccc6a048960eb63655ea35b028fdd87bbf3a75984673fe797b7490844be0de622fdd10d9bb28350bbdc285ccac46ceef21b9f949542f2a4b54d1b5771dc0e59550fb08a272ea6a1fb349ed867e2a335b773ad333acf2ab0a7e315e0ca405f4908b2f475;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4bdb66ea67b8cd8421c219dceae0109f6277d263bd9514a0d4ae694a9b8c442677f1cf6e3993f1a75e376d57f8bb23bd596d114c25b3cb892c03c0769cec7af24cd01c0171c104a817fbf1cc8ebbf05269da3f008124ebd050bcbfc45e555e4c1db51cf5d1b882d0dbd0def24baebaecb81d6bb8d1d1d1b7d71969880a62b29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bb70eeb3d2425c1797fa0d1056f08f66f67fe328045a09953ff2295d01b17d5b7847df0ea37182e252e9896cd8ce88c870d33947780d8d68826625349d9a49f70900fcfe1c7ab172f862c6bf39c0e306c5b04273c275212d9b646b60947cb7087cbadc4b475535ae842b277a4c72ba1142b849ab0d76f53afa016e6d75d5143;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf45f8609cc49378d358e23e270e72501ffc99cf36206381d3dd6c54146551143455acc5aab36733c55bd26a339100e1ea1dc5f2f3f7edce8772dc79fb55cbc4c1680bfaa9371c1f6edc93f0820313d5c7bf7093d362cc0b7a347f81cff92fb445e2962f522093b64ef054f83f3b40c81f7f001047ae4b43dc777bf65241abc84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87b5e1ad51afe654c1113aeec4a18f4458d9b7b476185c73a16778f253b44ea90f018abb3ec25eecdca8a2c53992098662bb6b73a521729d9e0c69db4b7e12e391da4e691bc2f90d1acca022d7c52163cf5749a60ffaf1652858c418fe4dffbc99f14723dd71d69235f7a1b8d415b459fc994d0ddd4b48255e545e76bc3ccd77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf783ee6cfb42f11bb98267198fdd33ccdd6155967bb712ccde08b831c5e2f67f8b7458ef07d9fe9b82677f516b30742abe83552246714c3109defd56c506b10445e44d015349db7bdf87287f1ec4a0c170995add0929d5af87574a39079e554932d49d2496d0efdc377ee79dc54dc835bed5dfc267b48ffee6afd660467c16e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ec9b994ab3732198d49eb026681f024013cc2058bfb425f10d5086cb4d75fcbff820633aaf10e41864fb1d2375395f92b29d13f74818f0a4db6fc6170b4095d7df8fcbc1eb8a688e64266921168b4732f308070ee14547d246371b66dc09824a142498a567039133f68a2da09be61cb43feaa76065f0c85e92ffc8b18df8bd5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ae75244778b3ec537a65b85b6aa8b36c40bdf40305c2b4504c135b931a8c9239c860321c6111f54ce977381cd6d93b78ba99d25faa95214db82a4886cc78f986cafb6bfc1710f955ed77ce58afdd7c572412b54dc4d8da0f8c50d1c7b91f750aef2c8c4835053f4a8ce7d0215888c0fdf1bce819771419b688b5e58f074ef63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bf1c6916ebf44da9c2feaef88e71c58b18f94ecc75b891f0fd5a9a09e5da5a05315beb116856d3ea78bfd63ea38a38e97953c15119d4167f53e77dbe9be8dcab06ee19240e6da8a95f40ba98b388df502b5266beb61854e06c84086096feb0e9072e1694d9da7f5cbaeb735ac7e9a021b4c99fa4805a48d6a2d6078a7b2e04a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21ee14c677f7956ea231b1ad15d7fff0b8bd86c5fb3ca9a062886ae1192249ad553c47d95ea8f9127e956ae68041584f6377cdaf6ffa038f25e58a879d2b4b0c2534e4ad9fe35766a1d5b070cd579b0c86688992245a427421f8c88119855d60e254684244f8b7bbf4a8131d413194ac41340bd633f7be8eaeada7d4b7e2d834;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4be8c8cf75309fd29a33390fc6f498087a315eeeb769206966dd161a4f1afd3b7453145b92727c521589c72db20a1b5e910ba1b0d737f8a3c7f3d8d2bdf4a2d0dff894ebabc76baa6a087d75856cbab38fd366b198b183c3c2c355907f247e5a90f6f91bf9d77f34736d71804ab964e2f0b4eb6e9477a4b5ef7414a295a59542;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ec67903a0ff40f8edad720bb90b959bc72f0f3f81c05f3d1a9dbc19cbf1b5860df29f054b375c60b366a45439c7ae5c4eba515fcb03d954b1628ea83872722171fe5c6a81726fea60423602aaad1bf974487a5c8f26a74bafb2648d2e0df04a854478ece9dddb4328e291d4d76b32d73bb85a51a84506753fb6f25d950cd83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f6a92e807881ec6931eb32fc14bc1ab5a09234076920f1c1a55f955a52812be04029f51e4b27351ce4b299ca30284ce953b3668e8c8677e545536ee2efb36162fabe2261c16a1ca074b5b9e82edede2f073d6a7c9b2b24bd539a6dcae575d67c8a9e65ff06ac7c972cd45b682bb6f5944a77918f59df322dc0676ca5431b946;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9bba8c9d8e7bd1d91618c12b8f947c0f29734426a2edb938ba25e1d440f4d74ad970e5e6fe17370b5293de2fe0db5c02c6aa7dd7461a92ca18996dddd966393a13fd515e16b4a6f751d2f01597ef39ca1461365e3a3a2bea1e326ff3977814888978e92d60f3509edc1d0e52f6bd17387452f52654b6e5ba190ac3d87b5e274;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he45a5aade69e8da966d04b77dc12f7ccf999398997c7acdbdad0c985fdcfe8e98e3e51f983056bfbb06d14a61edbd688dab5eb4cba141a30490875d6a79a23555bd5b65cf4eed943a563245464d492b3263b09906ba47abd7e6deb8c5841051bbd9af80c31987d4df32a3778071c2efd20d10efb8f7678601db923221fb6352b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37624884506a648ba45fd985e1da9855da4147011236d50d3e2293ab6fec26d6f9476f0ad9f565f1ba21beb646a232be1aa56a9ee1f924253ffb7c632e157e7203cc6a64731df50f68a3d3707f8657eddb779e8386219c3cbb332b8ad50923e0f45b8279ff757315e41587f1e1694e603acb90fc545bc1c885d060947ae00308;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb30296b422fda0516f3a6a9821a66d0b6fe8d62807642803f44d42ebd0efc25330a91d2cda074fc7082e6b8c22076091ea32c71a8b023087b7a1606d1aef1a673999d6a7f8dd8cf93f2186d5693c1b3a539f0a9d8cfb676a3a63ace192c71c45330aa04bf5faccafc69969290448dac15541d58348a64ae347d67a1ea2a426da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59e72ab7e4d591e857847ed12efa41c9b574a406f3b86cd3a75ea8d8103521ab237bd4e8b18cb1c2502fed84745a2715bbf74402c7dab17397449a022a6dbb64c8a4024bb6e89ffa2d8d013d8bfaf01956626ae934357a0f04cc49957045ae7b1439f65caaba2a57e409acc67c49a54482ab1b5290578fabbf2b25cc7c40bd5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h649cb9f393ec8fdb69be78f1dda71a845c8448b319c76f0ae04ea73b7d127cd1531498b9752c131959db0e361d7e8bc6488b60c6110dcccb2cbbd9f057e57358159d9f1ac16e4592436f8ae3b9f6592cc40d2b6251e217a6ab6f31dcde464cdced691d237c5e49af8b836cf2a7d87b1280bff54b914e828653ac197b9fb86fe3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51b1a97de0f14db15a330483a23f42accab176e1c27e1d1b633974e82c34ff6d25223033d97ee5fc97da0d451a2af1afc85d3694d00b1664f76abc9a47ebda0d4b3fe73e0f898b8bea0e3bea3b02c21a56003f344502b11340fc6d8c9e5dcbdeb9bc881f479a427a4de0bab9a1731f5b3efa7896eefca86ae702f32559514230;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf05dc94621a6ba446cde4c29b6a918d5a135ed13b23ade5b37e87fe1cb80db0367bf64f54147c4f4d45d4971cea5ffe2ee1bdac727cbc3ead8796c98f25881410cb7a1b94f5425711dcf9b9fcd47d2772e9cbad9e9fece4fa59ea889f2933ab29d7635cc8ee214456b9bef1013e7ab1ffaa67fc46e0e22001fbad1e0a0b74f43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f4eacc98aa29603ee417badd68ad13292d8b54a5d39d2ea4c2376f2f565c298095d9d62f2c24ec889cd538ca2dd2e84be2178237642009ca28a240d157e9b001fe0e63be87116ddccbb36ffd282ad55d70f19a8658c5312e3116bcd77b0d2a168aa9bbb3a6e591e7620d5aa0984c7f357fabcb8c93f15552e4be35a604d652f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d4d6822355f0ebbf42f2469d04b7bcbaa05e1dcc5356f256a9853cc8699186ed89fb410df6145d7a9a34e8f3ad0be4c9e2cfd4b0e9c6278c7e6e535da65ebb0d5d3d6cd14fc04c0966c961479e89e1e64542ca7627ef86201e7f5f194c7bad4b6429d4af7cc1b58c4eae7721f73a0a230cd56e4c11dd82a639f3d10bda0b459;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h446d7d5a1aa70f19abd9620077f0b5030dde3ee0c6f30d9e9c137bff74a5a06da6fdbe149a55db86242e4b245a1166baaeda5383dadb2537593c1be6e8142ec0d6e656c63d24a0a58db2bfeb25de088ac4c488db8d61605f01fd5d5f1eb436b80be5bd33332e9bc08cecb97756cda961f63aa5e8d69d06f2575aff067c7c857a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20fa93a27d162a4ed0de86dec57754684e2aa3f9920e753a603075021498f2a4441cbbb219deb8026d88bec18af147fabdd35cd6ab91952f5732f7a23767b971baee55a0c49a016fddce6460d4cc8f84560bd03137bcbc86422fea590405fa69fbcdc289cda73a3084fd13f058c5018ef19daaa3e1fdf4c2fe71e0bad457282e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e027e9d566740b1860abb469ae0080f55f276449f834e9579d486e07f0eabbaef2e49f4095169650fe2fd005e402169cf64573ea9f4b87e675b3c3fa4024ba2ce2dc8a1874973ffe19dcb9f8847e1684cedfb39b41ed97839ae68baf235316e26d16020e71a7ef07c7f00db89e5ead8dff096e39f900c4eb60d8e524c86bd4f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cdff7c21283b498849ceb8a9b8a8440c31b6dc35a00ff2a3f59b420abbf9abde490264dce3b4d4e8f31974683ab4644f57d64fe0f0ceb324144fd29dea28bb551c496c9e1e4e57b2e4fd29608e4633e11c2abb9c900bf91fbf56597e5e12954f84c0ae2cf31e2d651c54a54ade3c42bf8431fb453f9a61f65f885d185b800dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24bda840c09015074d14ef519113a2c1f9fce47ddbe50dab75676910b348093a1a200af5db6edd975f0f481c16c10a05208a4316fe2e75ee79d8dadbcbd2e74dc2faf1357b5392a1879ac7e1663aaa807e9ad576acc3c228efc329b11cf42fea7eca6cf41609871c4d620baca58cc2b58fd21063c13aef041942a8d6220996d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf355a2e3819384caa43a65229e37d838dc94c6cb49276cb6898e80450dd9a7531aca882f509c86447482629ae5f82997c02e3f817b9fe399a1b4a0c7d4abf4c40ffcc35d285a1cdac7249797f735f00e80722b60e7a559de83c5c964d4fd649c5d0527d95ccb64c49e06f32d79fa94316df9106e6d15b0c0b67e7534fcb95e27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca2dbd9f12955bcd75d6416f8c410413d1319ed3451970805cc0e0444aafabd65830a623745df14275ed9f29c144f6eba5c4a4eeffef84895ccf14db133faaeb7620b715373d5a16bd092a127cb07826d138b0d9a0683633844851921195b715f1f5c412db2bc5c00cf2f9a213d46f0acca7a8e748ddf3926fd4187aa3973245;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf687718840a2dc663bde95e6e5c5ba6b24840b269928be4894ac8135b2e0e38cab5f403db3dbda0b59dbf879bd60b58979b3da78830e9143aade1bfce0d1482834099960d2f4f457d88f322d6415d99258bd13b17df3716bfc4bda309eed5d0f97ba60eec7ec8fb2097b6f842255621591a8e9388959c8e30ba8cf6c5346c55d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3a29647d682aa2e7b3792e75c1a6812498d2e638470561a17c2f609b81d5ceff0463d81076dbcdb73541c85cac0df70fb72b2d35ddd09f3491eef8387b645cfb58675741318c070c7a123e7c4804ba6dbd15616ce8127483249444abdf3107e52e103d75fe5c68b0183a3fadc7c6b8041eecc9c99c2ea59a42b407b197a383d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h459bed02b12981e4571e1cc3c9609e119d07346af88d97dc3aad290be333dbd07d9124c2f6019edaf1e8dee0a2e32688207203503d1c6ad12b9f237b80a5905043a4c4beb06992d72c3fd202438775f2374551cf7e624f9793eaf3b1ba3a6ed27e39cb7ca7ad09b4cdc3778b84cec162ddb6befe8197f470b999e99fbe1f3d99;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h863689d4ec2799baa6c797828eeb310ec331e7bbcdc89ed69b007ca0447854a58cbe4ea5dd8e3488134635c4c0dde3bac736ef46f2eb04ab5ee9b54fc52fab13df3a337bff7a50620ef546cb3e9565b11eb97a90978078577c0c849387b5f6ac69c7f38e3a602c07982d5f2c7a63c62ecb6fda0350a4f26b5f9d9dc2766502;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h163bb5d15fe0d7250041fc9fb6cafdabfe158a2f801dba7489805706097fb48da4f592c306cb61b786404f3ae297688c685ce0272130a787de00432f3478d15b2e2efe3d7a9612f2430d26a2a2db5457255fbd5cf0c402aa866aa822ef08c32d1b49ae4d4e17d13c8a89d2c103d54bd1ace1fb49a6fd67fba1d04724962e29ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5936f8d82e8c1c80c7cede66b424051d4e7ec40dd609f33cc76461b8290c6d495ac5eb243887f41952ff5457f677a1713bd6ee2c076229fb2e4c402e3263afd5b64bd15c79fd59b66ec2f26e6c235c1c3f295c52ad7761f32b1dbf892605ff689d7db5c6f1865fdd87d4cd9bcee9f6f2abf415655cdef898d1e64bdba3fa1606;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a799bee9bad620bede69b4b497f5b2ced0c4cc955f3533d43fd54f13acfd8015bbd5148a23873062bb5a8d360ee425929cdb10514929f2f39968b7002c0380b6133aa5c5e64fb667415ed11ab5933e06c97dadef9da5bd6b543eb9b67ec288223803af83ff1f61e0d9bb8cd3232a26106d4797cb2244a84dc8846f3a90c067f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d9f85703e177917722e3971438f9e9fd288d0c3749b7772743d4466e522ebc352d6c8a8e9bd8cc8e26137de21fe078b3f1b4b12d3f3a45e6124ecad2604e2693fdeeb54162de9c9e19f4b642438e8e0e703e7d9d53853402211ad959149a69fcd0cb6db375b02ef481623069a5e2dc9df69e5dfba5061c8a8928309eb3863d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe2fd9fdd157b1a32b9c15cb6801391ef2b02f889990c06a382052bbf76e24ec8088a222a692f62d05ce12f2c688cd8ae167274254d77dca7324bd7973501f9e83a97c96d61242065829fb7a452241b4f5575df4ed568f5f9a9355375a06ea3c8a23d175b27b0ebc1d01aed38e2a57e0dacd662bb3aa6f2583578c5a05a5ef8d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cb7ba2b0435c2a4e29f2f9697bfbe44a7fb439b40ba9be6a1b060634deba8205280c61c7e21d8e6347557481f84b3387decc2d5acf42f649ee180bb599dc4791211f28f75d3be58835452765b6171c603914c284163d79a85df078fbfaa9029965c3af51f4bbb52393058cb41868c9553150f1568172750f1189c0138fb63ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h464b3c3117a2edc086ce58f7fef1c97e4da4ba077a32633302419019b143a12fb3b428a17a52e226fd806ff15a441ee6e79459538f5d6b12e1e900955183214cc8c5fe07e8747e3acaff71691fde714ff7486336b3675fa50de762c0d4c719d9698d0d8824dab3e71d53c02fdbabf932feec9f5ff2fe567120c3d7775e0568b6;
        #1
        $finish();
    end
endmodule
