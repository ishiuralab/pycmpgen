module testbench();
    reg [28:0] src0;
    reg [28:0] src1;
    reg [28:0] src2;
    reg [28:0] src3;
    reg [28:0] src4;
    reg [28:0] src5;
    reg [28:0] src6;
    reg [28:0] src7;
    reg [28:0] src8;
    reg [28:0] src9;
    reg [28:0] src10;
    reg [28:0] src11;
    reg [28:0] src12;
    reg [28:0] src13;
    reg [28:0] src14;
    reg [28:0] src15;
    reg [28:0] src16;
    reg [28:0] src17;
    reg [28:0] src18;
    reg [28:0] src19;
    reg [28:0] src20;
    reg [28:0] src21;
    reg [28:0] src22;
    reg [28:0] src23;
    reg [28:0] src24;
    reg [28:0] src25;
    reg [28:0] src26;
    reg [28:0] src27;
    reg [28:0] src28;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h726d1bba91453410766c126548cee42e2e4dbc067dd2960f4b2a78c5651cfdaeeda90a1cbeb987f3052258b3605f6cbd10ee2819c0037bd0ee728530820d683df06429fa0fd78a6ca05a808243a40b0e221bd6e0a0722e82aefce543d6cef389927a9be62191871956;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e294ef8aa21f3316703249b3469ae8ac88af1269e56c94e320d0f893ff67b6df3a434183a90996485df24d3d169860dcdbf63f393185a60d7f8068fa4c762425d666da99ff31fe44c5eb8f75d66ccdbd00e04759ddff75fc281d839af7205a527a694a9b87567ae5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1223f2bced4d98f7c42655812e696d15125c1a599eee935464b333102032bd69969665e8aabb5513f8726a4f54db496229e0c4c60ee82c9e99e69ddfa06941586263c4e483de27ec5e996f0f402878ae8535305f7fa8190462ac132f84f446536e8abd915a58cd9d479;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e5094b5b35702e965694dc4584b0bd080072616ebca70b7e6ac72084ac556728b28aa9b4beeb194685354ea87f76eb20b2ea967328e3342013c196b2b368464dc8a9d6f54052cd65001a2e32fb0d0e03ae9efead0e9f5bb0f7debfdb2e9f1a778a3aa1a83f8f224a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27526afd0f2be9375aff17035b46bea9f75bc310ce5e4c893fc236ff405070f28cd068a94a633618f16a02b8f35f6cbc5cdb03e39af72f7a10ed81272b19c625002bfd3ec76e2fe13c6e28fed8886e32ad024304360fe0e512ebd4a0ef7d91a0f4b1b7dc2b3513bd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfab1fec9e1f5bbbb57cbfcc159e1a86406b029b439e47becf286c9e4d342f23668e677c9e37c60ba5d6ca9f9113088e4a0f1ed3be61ceb50a6dcd9d881ebdeff1183bb515a618fbb2c23fbeb7a9b0cea78ecc44980eeffb48c2e814d0faa3aacbd5e9ef27bf2e0fda6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161c7c1cfe9fbd96145af9e4e2f1fe9f16a2c903c7ccf388b4f09f7155687834f5833fd41d98bb7538721fab5904b2b93b05af9ccb4e120920f6229277f12159458cd61f9f98820da1fcb1633954916d57e422adb0f7fb704a8088369492d78c5fddda3aa97d4f44c4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bfd8920200846cc68f7136184b23fcc5690d58fcffc7c003365fe418e09272c703dbd427896b133a906c0fa4dadbfb5aa95b72f47d637762c79dd660cef684e6d0e76854dd8d7565d6980379f3b66653f29a40d3a15fa5b3987359253054fe274233cfa419a201e14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18478281812f21b6cdcd62cab01bcad26a313abab5d502a93cdad1e9a99cdc35f785fd0bc7e1bb819e939e895ca9a1b59b026a912e4930f76bebd754539e4380718fb72a9eeecf7f30848169c7a3ecb65946703b910365857dc7a1746e83b66e81c181141336e5b4479;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4227decf12fdbee17c56b04975a390cb4d004e735014630309cac531e43431fb1214395e43ea9a7b2f6555a1533f3e18f580a469fecb4080f8ae91b353c7c8932ac42699e0857e5847c1dbd49528dda811d74482df7ec87f441be8d80b0e8d88aa34e71c0cca832106;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ecdeab439f42cf522edf17cfb2f5417b6f9ae435608be2e4a0148291a52ecf76fedec08b76cd47d71b36ff513b415851ba5ecaf18c5fe88b110a46e4856e3cbeb6a0197a91d983c73d010e207d5a1b65473e5e11cf975d55c7410298c7c8e3a942e44bf140c161618;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174aeaa1841558faeeaec845d1f9b6bbb932ec7422bc232aa01f4614b1056135a8929a32f63473592006c79e6a2738328199bf4a1ba0164ef136827c18a612ee54937a051f18cef64797b26f763da81fd80edb30523962dcb0df70e91e347dea62d13192239aba3c114;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4e39aee6822026826f53c0a6c9fc624cd519ce7b724a914b5577d89e669162228f1a284e49398ce2d7a3fa516c4c48ee346941f5c386d4b4d515ff6095cc19be9baa526d7e36c90f98218eaa3e979d9debc3d8b40d495edc0d8a38c9be5af97a3912995bbf737b4bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14169b5415f36a047137b98029f190466b35cd76ff5faca29149b07e6bb25bc8c010ec81e585741a51c3e3e5a64233f4d3844c5e38440ab4f6f0ea8377d0122fd4032339e17b3b610e812ac5110faf3fe24785586af76a8b3d764c2ce00586a74753ab444214610836d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hafbb4e9c419e91506623adf234f2679d8cc8887d13324fd5d55de2c9d416537575fc75d7885a5b0dd2a20751cc9ab0e3a285144aed0401fc7b99b91c035ef5d1e8e9712993e5a580fd0e086a871091aefded33896b53b89d7d221fffeff62836129a5b22aa40f2f4ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f28048b8b9b97e94cafd80f8f3a9a827d6ccdd624299b41db76d2a904dfccdea4183013cfbef3672d466c2bacfa21472421e98b6ecdda2745bcf6a7a97c00a73fa10ca0f050d0c06f580e5e0be74dd5d19f877783143c050e9b87dc9653efba6289bf2339526b659e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f4c286a887640e00df9f0f548071bf4fefbebbf7b12dd82cec0ca7d07bcda5aa796655db1f0484068acf7a9922f6189e00f1d186240854b6504c96ea1e3405c520beb3b067afbaa54ad9a0aec295bb27842881035771bd1fbb5f5765bd79d05c8f22497ce6e44176;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e37147f89b2cbf93165c4e25928ee3060944fa298b8f72bbc7917a66c6cc5605bee185e170e8a14d6384ad5198c0d8db2b9462d4845bd4d017c60f6d454c22eb6e5937bff8e86088e696905358a717019dd295a670a9fa986a50519ce8f64cb181e75780db79244dd5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha921a65f84d77906d8080bc51c702a8fc6094743e26ff62c693122a1863b080552be3d5586ac62817913ebdc5e584baa41c05235e72e9167c03d77f362c5c80c7f3c611423ba236a809c47e28529103ce8d01cc94503d252b328f1a59aa362acb413fbf500577b647a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcac2bdbc66e050de2ddd3d2ed8ba28d10c6443dca3ab7b3d6fc457747ed73ca02b1a88b5b353aa6d877979e18456b5ba44a31ce1d4aae0867320f488aaaf586e45af7867807716f57ad9c8ac960b06e5d2a30492c42654fd9e05382c78948c6f07239a8ec6db53d7af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b604631c1ef413e4018a3fef0b549761f3774f27525e52ddf26e008f12fe757b99d7f308322c44fd81a0566f325fc71d13cef62159168434c944ef2f677f47ef54cdd01886a99a6667efc85892c0ad65cdaf874951f28cf7481dd7b018ef985218b00d55e20a107aef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc92991844b3323d08b2cc73e7c26e397d494bfe49f02de00bb29aaed5eb4fe01cd9cf763a4ea7e38e604327218b52f5c0f32538753934f3ee01baebac283d0090316d5318ab80784165bcd15991a5e4e8e1dde6e929bab7ff4bdfa2ad2def563281a79257f41556cf4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0539be138786afa9c3271f62e3f42526110c849df2c537eb22f2523aafc57a3c73d95a06e63ca8e6c8360d09a418b0e9b827cd6ca4d0d1afc8395b9b647b3dd96fb15f2910dfed4044fc520657a45c8e8f8d458f97c2075297fb968269b096a93909775073c4bc3d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7db60754fe833afe1c0d807d9baa47efd256d055de2319145b0028f4bcf9a087c4af9f8a52af8d4d88d82fb9a87c3c50e88a3602d6cce2000a4205a2931c5456d95381893003e71307063da2f4f9ed2ef1d816abede1729add8d3409a5cea2717e04530d2f8cbe93d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36f800586977c6b2d29363d25bfbc4e4e895f34dfee5d6cbd478031ba9c236875d49e35959c959d44c60769646cae01c670d9a32104ede2568f3d49d14f7b34f6e7251adbdf65474bcdc9e0dfaaf39ed4624b3493d5d4f503f49cb789f7442b9695bdc253bfbdea262;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ce61f85016c56223b2b87addbcd6a9ebd1b67f3c5ae1da2eae1c130ddbb586c77c2abd6d9281c6a05506217bbf2213846c1a123d799bae709753e258eb17fcbf9b0cae274adf7e321d8d4443042ca01b064b6fcf8680ea475045991da757fd378763751390712cbef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bb960a0476df47ff030c688feb326f0690ffb8e3326c2e3fdc51f3d5165bbc2b09896fff55fd634b1086f57cc5bfc8ef497f8fe467ad9d7d4051d90f950ec745927049e1bc21b67cd28c167381ec6369d282e32b94fffbd7276c4bc26122c8485e9b9a394fa269f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1979106f57f50f4264184b21998132a21468b707126ee3e15d0548830a368af90d32d6b7e55b7fda1297ba9070a457a84e8ff4a513817410c6c05d8277804a25f2d69ca532c05da755781b1ea872f3f8b7c8286cedf92d9c447f767f9416c0ca209e3438a3bb1dc5db2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1142fbe00b8073590124cea8a3cf9d761e5d951c8ef5a7fcecf15be9f16f92eb82a5d6d0b177104b8740439546f32a19b29c070770760790137bcf420c5d1cb3fa4ae74610c68cb365295b8c749b01a1a295784d1924b0256ce2cb8428bbbb72186704ae458acd7485a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe593647e5433f7d4ff58699d0e940f9d108c3f368b923ca6d89bb8b3cda6228fcdaa456e0d9f65b3627a39cc465a7c9261cb5a10a5cda57cdb5d3b4e692749e38bd846c830e008640b9c0f5e4721113b1bb337c0a7d73fc587b836a28d07e646681389f353cbaec07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bfa35419a909497ac3bb2c4da222221005fcefa0f23c86c6e9f586d510a553ee973f70bfde5e556b3f3f4a2eb21db9eea506bb936a7221b85b021d96ae2daba99f95a1688960ddca21477ac77b0b2969d2784c3f6444e034a357ee89f504c65018526202655cd151d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e19b7dd27fbcb9b3c986475f2995697f7522db37ccb9837c934aed9b138ce3ceecd9ce98d2dd0225103263d21d45c8317f1a52a562437b50cb81f9a84727362fba99bd934a6eff0421e6bd3e9c15d24a631c84bf3cffb62272fc0f7e3a69171421b82b0ee178741529;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f951c0b86e3aef57c64b32a53d3d59014e13980a034fa743540b9c6ed9361faf7ce837cf8414e8366b2f78994b568b2b735807634627746e1addedde2b9ba84cd344d3b619cb6b14105df9fa8450ada2a1653673ab9845038d9544b7ee3fc1b59b908c3536619ab26;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7a9a6057c2917ca281c5d96005ed66c5912bbf94f44281f0dfabb5dcca4222c033c8b1330830dc5cbd610c73672f3f0f71663ae61548a8fbee0c838fe7a9417e4727f2a1c089452fab17d388a99a2157b6e0c5a0b74317f9d7f054258c60aa27859e055db1a2727cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87ce0f0c694673392a292498ba0a4bd6ef1c3ac6bcfbf686a0aba1f01e97291bd5578c9dd4577e28285eb7c62a751c7c080f655640e152cbe84412ce079dc56ee7fb9c8e0105a9e0d6ad804755873332c114cd0676cf506e4461d5678b4e8126774bc294a0d81e9134;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad78f5b46493ba653492e68a8566b4c93579465aa008580d7f5f7d19dad4366ff9c63b85dacda156aa220dd0c5c10446f2b6f6053cc78637d599983684c6639f8ba20c2b191c55a455fa1a471187ca4d59b854b7152ed498f1fe746e7d750efc17c9fdf2eeb7bb5d80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d96bb62f6ea1a6d16319f0811e0f7b24d36be5ca2769c99e8ebd9d1f4d964cf9b2d3e2776f0460ead68c93d71cb296f18a850d86d437a3734b419ae41aad8a36e1160f803a1a3f6481c46cd54a70456ed7caccfef244e06d3d8b166f9f785ec20194d2fd38227324da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1624753905cf1d81190b13ca2f05af26156b5b24bbeda80d6ae87b6aae7a7b8765814c3912d44c15d1514a9978d10f9347270f72b291a72c5fb26adbadfd4d05afa77d6ae2a7f33b32b2c89d91ab2f8c5af350dce11061b109b3d7c7997df1945272c95677365dab11c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151c663b95a27428f9b0b8d48013ab985ea6aff87fefae1223e0a44c8939c8f7e5839eb76558ffa1f5b5b9e171872caad5f2e15b2818a3553e96c5ee1ff0d567fa2275d4f43a49125bf05d2aaf3f549f514fa7caf643c76469156dfae8e69170024ecc413c6dfd98cd7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b9802af3059eaadc443a48e8ca621bf03b4c26a014dd7a8c76844aa43370e4a351b2b2facafa83faffdabf140a669b861d144da83a80802fcaa1bea6fb6cd7f51033fd0d33527497fd8ca305d7e435d1e757e75d6b51cbf66377dc734cb546ad6492336a2af9a9c4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3737ae3112dc94c6e5d2fb2d1275444fd74aa9ccc48a5afe6dceb5807db42ea2661b9217f439cfe83913c46e828d5c2acf76f4e60eba8011058b3fdc6bf122f844e4849890b7f709e5a410358e67294832266e01db08765c48d6a13c84e85d799e38ff902531ecd416;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130f21b64682259fbdfbc3544f7e0e9dfb17e28ec9846158e0dc44b63f6ce4a29f6b490624d1df752bc54de1fd609d8dec4bfa3a9d42bc7de01a4b156e1b4b483a52abd2320bfc5651e6792b1c35a54b6e133561df9667ecc7ca214216fd55e840a8d31c15383ed3581;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1241f3a3b7eb11b532bb85875118b5cc4fdff488401ce69548ad23b2f78a77c9d342590cb7a367276b99aa33d350ba7a04c7001756598737616e1dac11545ad02c083132d22781181fc0ef875f0a19404838e4c49e4710eec739f0a1e3f43928c0b3a465d7b2d58abea;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144cf85a12022d77997e8348424a036a45433923a0f690112de71d510ac24f02eb287cf5872d0daf1fa68250354e47a7448d5c648643d22b291a115130fb68b30bff9c38203b462dd210f124d5e315456379556a751189816c97978b78fc3dcfb87d5f008f115ec63f4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec2826c817e743350e8c6dc849de465faebb52e1a2147132fde4e7a50eb406561afabd311503e8861c56f54cbdd8d2a91f9b672a57ee595a1a5ec45acac842c43fb4c332ff603b64a518e6c36221420984b7f65e63ed80294448096c9971bd5e2aa46b4a71609df95;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170413249265596123f598b421e8370c32fa073d86f3d020c662fd60eae279722d16ac19559681db9b8a6d7ff3e7833095bef7ee686db160313e2e351c6b98c66d8900fe66ddeb903496fa2c267f2b858216bb17e4ce37564c872d3884fca0e6c71ddb37d3a1844268;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35bf8762d9734dca52cdf27c53ddfb4c8901ceb5324659905e1c69ec5354442aecc2d91490683197c12834f59fd53229dfba25763a9328cc3eb5a4717d7b4ea7e08d05b80fcccc222cc34f505108fc473fe1a30da05109ed8245f1e63afe235715c39b577ebeafb061;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b84c432400863175ee65cbfdd8e37011daf923ed4f379b6bbcb1b9ec5d7de932f51ac118e3e5876ae23a26d5213b6fd37851ccc916dc42075e64c78cea6f29f83972000f1632e7800c22178bc756145acb649c52ae0cbb030f0cffecab607ed6f41368aa2450c6df69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25a85da205fa742f818bf6cd007991b35a6f4429b1ab9c96e11302503aa9f47d04de2d2cb59227562250c620b0b53b54ce03ec46e9e75e3a8daccd58cdc30742812b7fea6eb8471a86f0c9511ef40599d561d763517380600d2b1985c0eb3c35ca0282b5b8cbae2d1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140cd80d2bb5f65e3f55d1fa95d42315f11a910422c0f7cb8bb7657fdecf208e9e21a58783fc5186a99607ad3159de0039f29eaae980bca3d46dcc3331b5e2e0420e88c6b3039b77673e7a0b27b1da58ebb0ff46d2e73e6f0e5a8e4c481c56d49da59ed45e8132b2bf5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d699740b9f643222138cacfb2349c49927e1a3f4264cb1fe7d4d71225083a54b1350b93e1cb1e6ab2e3a980146f835d5b3392411e8949d941f373abcd72b01fa82c2faddc9e5b373fc243cb4d4bba70f39c800d9f53159c0e5893895384bef6699e7f461bc0043530;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59dd6fb91439b6349fc5e7b641dc9b40bbe9d4b61c7d5cb25890f3928444e06d4d65267e7d0e168b86d68f41f3aaa3c7f187bb090554643d8c46fdb2bdb768251cf0892d6f714864651f887f97790526cdf27d8cc931ef37a59293b72c9ff903eace6ba680e8bbffc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14915e07d8c62978e8facc809f95f46fbc027cf85803bd527b93e58f376d0d2eb28f54559c102232a895868e001dff28db419b6ea68ea975f5fef42d5ae1483d0cb8ebb33173725c57d246f1007fba0e25c6611245e7841c1544d866e8dc54722b083070f11f1efe0b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e816f2da15ce4d2c1a8d4887175b3b2ec76d3e0411f9c50cbe478498ab8892cb6d793d67f02be4de43d150058526a1c442dfb2be36f445ee8f4b64e60826f3d5d569db79c623c4430d1d7fd0b21b0c0e39f9a8d606bac38355b73535e837ffe6534a734e59e2f448a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1667ce2f2d0d68f8c9127fe6557981f6129a36d5dfe2ab1cfe333c729ac9b285fe954a9a1ff0e30db4a62648636f0cf6248823fd46263752268a80a8184fcf901f11c44be60787502c6591a53079635d9261d5e0c675ff786445de1d826178eab153418f148b7a0085f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44562a82438ab7e3ab18c23248fea036affd52c6c65e3a631388b18d124bba3b11689ea29cd48f61808fb359d8a87e4c89b43b8c67c6d5ca6ce457a68592893f02ee6ce28608c0d42e6a61d17a27345501e9ee1016db435d07ae05fdde83edce526fed1e683bd550d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a2a1a72904bf83583d67a377f3d9629454c3e6061f7131f8b98f52bad1edf3368c74a21066df9709be872caed3f43dce93844d73ab6a6e13405489c2cebcdbebbddda35d119da9ca1d8f4c8b8fe3994b98e80d8eb53c358f8afe649b8edb85cf0c4ac3bd452e9016e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h997d47cd5a21007ddedfa32fdb7aafca4b724018c6060a74be8c95113a04ec21445d29da1170f710aad7f6d5989c04be6d63478d0fe167acac2dc5d1728ad84f0c8ea39c88d31a5cea399095bcf93652c8b4d8dbd5f71fd20a9ee08dec2a09f1e3f3ca93d09b7869c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b5dcd0d1e11dc593aec5eb3a71857dfcb995dfe24430e36a91493a84a67b1e6e723ade50a997c8c4c56a9e38f832e52743bfdca151168a0f03baa57d772a51d12f57eb39ec06978994786ad3fa7c9651f6b49580d7565990e262316343117406fa895599a7bd625d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heebf3c9f0e56c3c4cde3859d48bb5b23b8dbf5acdb3fb089b4df11ccfc996f2565e642a8042c37ce79fc2ad70202f827b9790628840b80f8f7db008c726f44d4e687ca559d1ee50289de16456dae8da02a1186d1dde100e0c48ef4a801dc3d1bc35b69447780826b29;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcacfb2664e9d26f958fd6fe8f0364a7e1df5b795cf730481326444d66acd9a39c2666095e73db9265d6122312173bd6d0b696f23782e7cfd9f2eac006feeac24ba2c234881fe334ee3494e0582c8e44830ceb1442b64b6d1b069a48d1728f8d99ee8a25c5bd17e8f62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3be23941c53317962c266d454c45973029f616e816db34dd842c297f7509058511da1f4713f849f0d2548fef059cfa9ec25bb171067c648fec4ca5168f5cbb9b5a7f8a57bd6b4a46a067bf2f28bf3ede52a53eaa80f6df24c11a544db246568d15426fc46665ae3bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he78ef335813ab4ac3e196421bc54e1a3fc715eba765ceb7b083bc96d348cc20e6d47ae38aa1b9d4254ba4e72009a4da9bd6e65286988e6a3421399b61f679f46d570c2c00ab6094772dc2dceb7c4d5fead0e5043cab1810a10d6e08c526dce3decc39f4f6391a1fc1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8ea38475cb8fee6745ecf4699204250ac6ca92341582ab456d5e34ed299ef305216562034f2716bcc0ca882522ae1900ebeb44729f5398f49ab484d74ae5ac5c06354990146a01fb00fd5ef7376f4d94c2db954e230d769fe5d73a6ebe9112d8ca5b9b1b40e75d4c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5c7bca94e00c409c44f73f333eaaa81080bcaa7c73481ed0ae4fd5c8ef81121b7babd4a9735dae0683cf42d70db8ae2740489791f42d3030e9e143327c89e5f6b6669880ec66bb0d5e14d562ee701ded135d9197805fb07b78f29fae22f77799b11c91f215226d49c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15721fef67193ecafb9f4d0be12366ff835c596a495979645b2916bd11972f36c1b166976d8aa02c2548b33a5ed3e81e4e55ec6951777cabeca0a9eec5d35a48312592e2c0cfe3fcb1999b88fd0e1a3c21da82d22d72c725c56dbbc7ff4d9f0c8c31a8c805d2f103d3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e51f0583319fc60e3183c3a1c5bb29754fb95bc0ad3d91b36485951128796f3f0bd4b8b101cfc4184e045b65b646a257bd827fe189b9576429f517cd7e9404f33e64745249029e4b50c4d785431bf95482ef6af999c4a21ed7beaea14aca80c14ff7452df31211d960;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f0b7a6182fc0d22e68f47b1320a8c1956d12110cfc63e459e85bc68b5676b0814ddc83bbebffbddb52c632e9260cca2cd8291cacc1fd08baeca6a1240d3a386bfaa4ff199269e0fdeacd8ffe3ab3e42a90e668ed145dbfb7718132cd582847ddae1eeed16681b30c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb76e0cb5349a68ddc49a8f2724076fa4fa81a0cd00d9a2a2d052813827cd824c311aff6292fb1f44b84183ad946ca98d12b28f956c23a5bf95094b67fb93f6e49b02c922316079384be398663169059f50e75dcdcd01247435a35d150a4233d7d5c0a469e3fa3498a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f314b7d837fa8427b0a5b653d1e62be4e1a85ec0f99c305612d8bd23e761e0b83bb9b75de13087e5dc7506cbc871330142b2e85ad73d645196f342ec5b99daecc5288583e5a174fbd5fa225901929f0aa97307d6e4dac542724e719d708d258439c9d677dc75fe057;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179b0521c5dda3c5ad7195eb0fa4c44245ab5d7357e170a62c45746f090b555617ac9fa0cf60f0ad53ab05822f15a373625e7e5bef4a60d5269e1b8040e2587c3ced46241f7420353cf39f17759bd3c6ea69f21a407f5ea5cfd0f612c2b9d6cb26b7e09eb16609cb8d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a4bade7cbc553788c706aa5dd1fa0c0c24fb9846169724aa70e296d09626f40bcc05ec23f6f29a1c91a1c71dc5a9d93ccd9e07b9e0861513271064a5010c6fe92f1161f5db2efd1fc60d26a3541843977753bdbab7c1ae88227cc3bd6bb6ab8504aab97dc919754cdc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f19f6571800b9c6d128ebc2db1440606751cec72ae5d66e84412d2e2afa8f6d59dd262b32c254414ac9c1c434c79b8056af97dddc8b4e5bcbf7d29236b1f29ed2ed15042cf59390bf6c6dfa7a9fab0df3f4152151993f71311be5f4bca0ba738d7939ec4df61fdae2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9df9da2c98977774f2d1ba0d765497546ef2a2fb507f76dd05b95d3f64f89c66d79ed3e16f810d1aaee39674469d642f231b7eb1c3269653a445141d660841a46864ace60a72f1d0292b5dcee2a3ad00d2bd95f41fc19d499c68ad4a307483d8d4ad43da61d8fc1b3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b7bf33924f1fccf56f3e9c2b9b08b1b95bc1ba8d530989b35849c2845e6b4e25a6cce41afadb2ffa91e3c7d4f0a93f49beb0d39dc9d1ddcd72f3d078a7df7c3724db88d915018d3c72e68c0b9616d9f7baf0590a34808fe8824c67f59aa03b94be439cf7654f66cae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e911060259e8cc64610960d014b857e6207bcadae3172d4749243819585e943a24c096b27de5c8ebceaf7e30bff718b059ea2ab9d7f7d05f483ecee4d871a992a94c02b62f38ab89c99d9b059e7821afa1effa53b8f2309d3c8002041faa6fd50eb531a438bcbf7a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h765b48930f14497134d5a9bf7b22c088d04cd19b329955ad7df6dc3516443ba8277784b9fb05b2d03914ab8666385c23c385c956d0dd7063b231c3e6435847a790914c0fb4ff90301bd541a760353a9a02dc7392d7bdff1a14b9e252b0a03082ab651161e4add57e62;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64acb5c105f660cacae1e6ac12feaea9bd8100ce0086407e36c4abb6ffa98998587a9361d916f66a1410f1997547206e6f30cac644fa7325bb39c6099fb404b0ece85de9115aa2c17f5ca851c1e4e9abb620e8d13a5cc00e20e7408797708805005987c9dd78173e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec46a934ec0b0e6659e3cd4e6332d639ad4b90f070e96543e9a6bd08eaf4543a79079b444bc71d9a04d79f1e1c0a9a3fe1b3a14f535492f25ff0e6b08c1434b59d6b10f3233fc377ab35b3e12dd5a39608c98ea99b96beaefee47e4e998f988a7bb33a10f968fb4322;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11830e62a3667af19da1b56f5e1fb10d27ae2962f6ad1a1bdb567fd3fa787be1311d27667f5d0000c62e56f99a4335f7a196615d4f4c15faf52add6316391ec489a1acc974e2d0d650a9e31766912f692e320fee55691c074ce760a1813c7666b49b924e023a5127a38;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42ca5317ac7f72b9a4453f8967fca5d93e78e8d3601d50c63239a429839c9fdd0fcebfd0cfafa670ecadcce109289778151f2ec8fa887e3c2874026b1fafb26de605cadbab3ca649dbfc36a45a9e323fb82216791ec499ad1bb3451168130037c0ff0265277d0f77d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a52482e890ed2b6c5b5e01bff89f5e5cea2966c7cfc57b2d12bfc136c2122d8eb9f226b482106517c164d720e0d0e7b89e89ad0a5218efdcf443728252ebb483f2f7d05b2b1cfe5ea8f8cdc0a8860d2d26b4944df333d7184fe7d7ca53652069dba7739f0b17a45ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c36683e68c7b5b0ddd55a48f8e9d43e81eb02fe6029fc1667169812544429b32ea0e64bd2d3e43bb49145b0d9784557c8e4d56cd1c9c89035e0a4758e4b2ab7cd2452be6771a9d2e9944f5ed89c4ba2fb1f5f0f441937a42d70261313610a0ca410d4f06cd024d379;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd700f8a4d6fc09905e4ed167fc920d3a18adba7e3f9795e94c554aa22a55b738651d3171163e7aba8e1f362150d786ba7459c364e36a3c0054fbd44fea4fc0af3075a6b531dd91f45065c5c4b13eb858c67985624712a6297c5ed9da6cac35ac769efefb55a9154f82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0dd51d7453fbd86a424629ad4d83c6b335f23e79b7ca594280cc85ff9e54727a4f1439888ab6a6fb279db0867ec0e08a55f7483462f6179c3205c722edc4636eee12550601075d31ac7fa435553511dfee7e71e41a037847849930e125ef1615469d636e45f7d7ccb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7ae3720478b868b4786526f23684c6f2bc12a4e9394e941926f4c66af2e0e668730412077d9ff43c4b58da0df17644ae9a325b0c5171ce29bb2cb95077bb06dced05b1e5cf9e691ae008e61c8a5da0cb0125a9b62899b2678545e98d4568d0a4b1a682f3149198442;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8935eba921b42743a33615b3a088ad915f5ad65574f0565fe46f740f8587aa3984d70161d0329c865d06ef1179608e813d526fa060027c2423c70db477234b4ec55e6e61de3f308868ad56ad7ad31c60bb7894733e612e2e1a4ab5b22bc17ec4724bb2c9141a55ec07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3438619ebb67c39b6791f686d79671dec1192566086b57a870ca8405bb64410355508b36bdfea865a08c2cb8fa888a82a1923b90016f9b53e53ca659e8d470303b0b8b606a34782bf293886156b5ec02086264178b52c91cdc050085e30755c553cb5e26e9546b6c7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2930b9fbd8720f5e35da8d21179ff0e2e9d4013af45aeaf24f473182d71dc32ce6f74fb4d45d9521afe54d89103a18774c31aa991de26990f0dc2a0ac1a8b8db203300a71e0fd49f35a27aef8301ca5e1e37e6ebe3d67bbb8c3c6822df379afff22a2b6e621c51a476;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f18cdef7624b542f0d0411b7dcc297e5f9beb84a485c52ebf33793c125e1611449f39584d6af1e09daf7d76e0958a45fd1d0910af08782596937da7361decb5aeb7acb40fb911dce263278d6794fb199bebee4c3a685dd6f65f119a6505c61b7ce81130b35c76c13b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d01f2d86a6502b4cb663e721991a8225516ceae527cc2f824bd2f913d5b1a05782c2128e77d0f66409a0170680eb3ca52bccea0ee694d559bfeed13f686176dcdc838a1eb34e2038c470ba304676a82b2829745fa274004e32db640b94c0730b1763acfdc90e94f8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18631e636e7306a6c34bc896cda589b2176d466cc929a449e0ccceecdd7fdaa5703c5b2378f5e26b69b677a9c9277264f7bff04fdc1cb451091622fdc5026e43baaf14b1bb7c8dbd101f7aa351d3a7d7b7186695f156e209217ab115956e959a3c87e523a7864903a37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142d41683053e93e08379968023b00d73631b28bfcde349f39dc1e7aaf9c57eb79c0a4e7738f483d7dfd77b1b0478b9f5744294e36c59ca9712286bc2472a3b7a03b710cdcae872bd06fa997ca273e0edf66b380add15f5977900e40f6053eaec3f30043b2e6f763e37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4fff6210168f16c972161099b71e4a4e743ae8a902f2795f27c704f7edf6746ea5e8c6b24d1d2be76153b33d13f0caf17d014592eff85a513e496ac5f97d4bc833330b35b2966657bc4f50258509a41e051ff2f45e08b91873bfd5ad5838470db8afa76f634211051c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fad45483865839c717fb83fa890ca214382789975f35fe9d57ab268bd018057f06365480f3614caacf69c27f833d59886619a07897a85f436c930bda1252ef83fab42d347e10a07abb69f8e0c46d88b777d24751db026abd3608fd47027e896c64f4dcb53aa7e3abf2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f4511c2f8e1027d5edc28afca760b701fb42d63234b1460f1d74754a7b823c3f11d995920d859831f849c28e79e18b512f05d00c78c559c4c40eea98593995c90e4e249e72990b5e77bd77430cf3abaf7ed54841d01a192b74f182507dbb27b3ae061ee0f93a074ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8284c3204f0b6bf318eb70ad4ee3123c1f60d1ffec3122ba3a3a80b8f620a5ca744011cb41b1308421e10c1390a023276777c69d95823507dee97644e8eacb73b74a1c31dca8fbee7e3bb411b3505d5ae1fcda8d5b73d117460b9debbe5db75b7c084435d940f1bb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2253484701e3f867e8eac5d8811c12eb61b6be99d5c5588c3d80454be942bf3448d4d928c7eb7b246c05e28761a2dd22010a4271933fd66bc84891455e25b82217c5221d484a067da8fcffb85f3d8d85c4f349e8fee31d6b2c20d37bfbeb2c537761562caaf2635b0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eab39b8457a9a3a916c9f7131ebf14f1c8ff5564cab1db3ba89e2468d31e5a8c540a745f5aec20dcbc3cde3782bcfcf0b39fa850b7911de5f59cd83d1e913ff9da421942f8eb012ea75e9dd5e2661f9d09b98997f6917e240615dfe5e1a6e167eea17932fdb7fd2268;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha303d9fb13dcb3000d4d146beb622e1f38826217b9b6552cc6788059eab4a1db1a105da8f202860d6fcbdf60a34fb29c6c9875e6e07d9f8edfd7671e7b45de77a921c9a645e2b395e704de10744ac7f623460a3535e2cd32bc0e6e3bb5d2a3c0f5a2bf99341593ef07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64aa8d94407fd8ab0fb7ec8aa2ce18b7820ab1546c21d262763223d751ce2dba11641f78f5e70bac08822b3ce56528b783a8556198da53d78d26dbb4e59288bff16471c29b829d1570580301b48436fab6a8e7d38525949daded692c86590d2a34f387f86b9d22b99c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117c187106dde13460df53b8581cc502377a2b77f8cfed5a089981928378c2aa0a4c0bc31842496a81ec8996d1bfb36839d41985597fdede6bf2c01feefae4892c006de13f928d1dfac3ac499ba6752e0a2669efcd1b8b4be2915a77cd4a54c66023a027825742a79d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45376113a9f102287355ea4c3f3f6efa8549bc7c3dd02918c18a60ea8328d2b9bff0302d64c3ca2f716df1e52e17efba0ecc30d2d807efa98c6e7e76399a9d551c1b722bca738d22853443f05aabc957d99ce5232ff658c157d1e9a962a16329d4c6ba7ac995c412a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b389b3fb28517eac20569da0376ab7740795b0e8f1dc1e05172f471937782f2fc5f82b09fe8be66662cdd3b3090b674cc1ee6b9080ba53441605e2bb3996d5349cf3040e3e334764908393ab17ca58691acaaa2016b6660bea99a9cf36fdea330c38bc8709a618055a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h919c86fabe9a759b91a4a1286f54bab437dcaef8a48a91629f9e6b30ff10e48e57f0cd640c21cb0eba8c9c858fb8eb05d098f0d50ae28dd0e61892f10253ae22ccca1828f8632635160ba1299e39061ceda6fe3f1f2a65a1b84babdbd9fb1309cd2d7764b7a35b9636;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138a5b6f32daba840f5c00966f6e4e8c5e566b1c6df566f8d9580728a6c1673d0c84480373fce5b764d06cc61febc1087425f02a14b61184eaebb4bf218629a05217ca8255d042bc6b98488b1171f2161532cc2922e8460563021e163ae76a380fe2394a33a8168ef3f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a9cbb1121901a7a3ac2442055bf116cc8ae0943bb7989c2b7dc07c2fa0c874341e5a784aa4e6d35f03e304a40d70caabd3f7e0151338ca1632eca6ea62c3c3dbb2b066103eac4b15193e01560d366af41e03772c88145588f5d77099d17b9e3aa88f5e3c94e138309;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d93a834d15c59eb8f389bb02930f76b96359ee960164eddcf40a84decb848739b58ccac8ceeaf8358f58a4de7b48c9d7ab8f79136bc5c3b8867e5b8890026c9f107f3e938f2678827ce1425da6b9a358a6938ffe7698a260a417f001ac747db53b2b28d15b5e9db5c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b42d498146914b343663441f5333c9aadc2bd322ada79798c17e523a11feb55be62a16be15fb73faaf1b2d1ff07e7c0df35a333a24a935005335421b03cdb8b7dccaa7185e095ad889e3251b859bd41e6e8c8a91235800117802f7499ada71267ecc02f2faa92698e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2bf9b46288c9b10750f11cca229248c1408b6c9cf529b6bc37fb622361ff904d10b0fbc1c442872c9a74ca96b844d4e2472914201c7e2a76bcd93c70da4af48e5224780165d1f605417811d9d8e2ebf3d0cddac8faee2f9bf9cbd88607560b9ef191c5773cda729488;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b79018b21c34d863d6a14e2a5a01ab0fceb16a9a04515b6f4f60501434e0904ab03314e7abfa9403d051d0132b68551ad1f25ee89cc3d9a9879a5db58646b0facae43ac63268fcca57b816b172830e7a0994f922bd16c4654389a01742d088e76502796bfc60b34e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1193c4bb8aa5f3776de2bc84b056b11002b091604af97d1ea2363957e49bc29ae70d77e319ab19feb0d7701ea42846700a1cc5011a849927b680cf2ca69779f8e390b69ff34bddc6290837bfee28a194161c1818d367ee1efb5dadc8a69c82adc4f4334d336f0b084ab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8a0f0de9e027d43fe12f49c2eb15adaf49358c7c2b257cae5016d138b97cbbae9917507fddf45b30fe0cc3606776674136fd976b96a3fac6b9c93e2a12b97d6a6fc14f82ceb4ba35fd2e006266226225a12e3541b7fdf95aaa7f83fcdb258de5ada77dc3ad40c0012;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae8e99227b3f79aac6d5d83af6cac466ee91db97bfaa615d438ce1648331dd41783f77de447d2f97f9b57a4a3a904da89b27d485ef99f704af44d7cd0454d22fe7b98bdb0b91f279a0f2b650e800f7c8989e8559fdd1f1fe029cb28f491a478cab73c2ebb3644a1757;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1896f35ec02fec50a9d732cbacd0a1d975bf17cebc5e9041e2d1ae849bf356f9c0cca71c109843ef2372a08600a5244ae4e0f4a44b4a067c3191154d955e989465fe91e234d63e55a194f9faa186ab5e2a57d75bfd02eb00a1bb31029efc825ef61180aeba761f3be2d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134b8963d99280bdcebda4f21bcf3f41bc2ea7d6db086d3d2f40b9eec2cd0d42908247ec62fde65e9221a82a0661a06930d59d667b696433244b8f69306ceedf1d0d63acc5e0c9017038ab339681304dba067b21352b44a98e51ec058eadd8a041d6aa9fe6ad7566cfe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ec5ad052a6b43ef910a9b0af8621979dd1c14269d389d3a764457d2f67e28ef110dd7ecd1cfb16ba7f2cd469ebdd5df0829042a3b9a78a6619787ad08ed7c65d23b2c1e5e2621a53bfb6339aa18afcc008910e88dcc8c9ec2b9c0eb9338ab5fb0f4084da7f2bfdec3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13fd13fdbc5c7f96f3900090a23be2b0467318158c4bc0f1c0b0377dd015be63fc9b98e0eecdd81456b71dc4c3878ca5e502d6f7e57ccc8db5bce2b1ca1ebafda754ba8e66c415344cb44add9890ca78eaeac024bdd8e54900d17df630d098330c3d99c59e06a07cc97;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8207fc6f5042d7af72a84c835dc7526932f131bb87587be90a9fa6e716c559ae3d07d8d39a66a24512b01b421f0a98c45e4cf67b44d5d7b96e77339f31877dc77db59dcad94a01bcf48542701061c86a5acfd21942b977db6ec3c6028dbc75c24c4bedab64034f731;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he81212b084aea11d50715e3e394a8072e359ca3c519fb8e04fd155bcf41007c345d31ea1f101b0f285b77c6360dfaae26a85af289365a2f18b2c6433410fb8971084b3f8bc0f1fb684fcdae1ceedb42b7bcce53c1d3b8835a4604aea017d775f786c4492eba6357914;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1669e9b923fb6eaf9c9f9cc2ac22f06260d70ef1baca9abd5fd6585beb2c46747075e53b7178a39213c4a643effe8aaf050df657e044544f18808bbfa8db29b0f9315b2ee15ee6c246cb67310e9eb6fa7f77f2a6e58eb1fed46996c542d2568961f66d69bb4a5760f0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7992d622cedec9dc5ff9379f5d1444d7046c04ed3798bacfc4d05d409928d5c8ef913fdb44a32891f1dd6312bfb538a2297db644db331ef58d1fd7b817023376d40c259165a98352f55becb2619fa03b02b1ba24d670711a145c2a339362badf3a0026dadcf0e60368;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1590a3fda5eb2fe0ffc0571660fd1da6d2d9a2c8efcd318dbae831a5daa2729e7d34079f7472584657871fa894104df1eaa0312d04010b14b3a15044b24f7adee40cf91fca56031f58e16baf7616f249c4eb95948ce79f03dd2c45e48a416b7a5d8376450b9b66426e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h967354227ea48480d955d07c87bea0d7edd1820711144ed870b136531e9cfb60be6d4e36865b5d58a5dbfcc6afadaa9e302840bb407d4d75b458fe37e3daf5f30e8dedae361da2c1a18a752986a886f716b46cae16717406d54f118f2d255609e09acc98232914f1de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfbb323e9536657811a7fed244adc1df0688208b65063d0200dc7a9b762b0e80c2edfdaab09fc818e0ce2d85248ac2175dfc95aca4353ae106d4128c69e8d9ea79dfe0f40bc0d2f4642226d9ace18f34f6bd7180a0bd2922cc9170f3108dd6a4d02080010a1a423a22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d569688ac83ca7adbbaa427894a6c10b2243a6018873f865b689d56b45d253e5e315ae3537c23810014b02c44fc5bfa3ed7a7d64ea7657ec29480ab244efc258b7ce6ccd0b78aa4c4468f193bd80809dc091c189bf19741afc6f483371943aec7752124359c5a2d3d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h304d8f470ca33c9a1d28f2b19b43e1874093c73b418464ef235a1ec48824d5ce51878eeff470cba5dc02d2112564e19a2ec879bc938073b886a10d8ce8796db3dec8449942a1cf3512f7cd1ffc7a9cc05da6ef93380a29a326d8e884b7262576950823ac58f058ea0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30b22861944696ab86da4b76c923874db2a74d69f3aed3599e878ba5a3e011ef57f402afc391340a7aac13a7d078dfd204b827a0fc1ba7c8d79dbeb55ef4bbc050fa496c9f8e3ee12fb113891b337193d2ac4b6238bf0da5d48f54bd804a903716135b7390154aecd1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164f9df4f7cc64ab337bb936329b5d7ef39cfbd8fd82fa0b4968625ae42dbb47b2d697557d721be62eda9ef2b406d9e44dd27008718070d26ef50f92586d572bb060cb637f63d316b61e7ddf069d67316208da5ff601568c13d41035e017515b2f32f25a101cb3ccd2a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e048684b36010977c9b2ff8aaf63bb9ba16bee09bef3e1bae180dfcc7d88d8e32c422cc5cdf3b9fc3b6b13a22ae92f400c599755552f6cb7e348875e6d3815a2de9d26fbc17e62385ab64af30702f7c907552333d8de14a59b245806344ff8777487829437c291709f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30b212a9f35f785ec39c0486ace50aa8e024466ac9b8109a51d2f58d103df1b91dbdba4cdce0c2d981814d02def4ec2dc5afce1634c4aa41ae257ef958448ce141afdd4e26a0ae1f7e0031a46fbd7d83db98f880559abbde0030e79a2285c81953e115307cd6e45d10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a22dd5f5646d0f7ebe9c005b5f1239f2c6e068f6e0e92686f35e336be35e07de9da628d18e0d100207c250e3dd0a784a3fa2bf351b387b6334ba62065e192de2bf16eecd073b76d5bf716fe9ec917d30df8046d3dbf317151f84ea0a8828806de5f690b4150ae5958d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f0b77f4244b5b730d7700f3a0ce764d46af847ea2e7cddb1ee105eede70cb9941767a218f0a332613fc3c8f3231f4598cd288f60fa568dafccfbcc5c37186944b72eecd33d25daeb28b7821d15c5c0292dbd25cadcfa1803fb84fbc45c0359973fd7ed08b8be9fdae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f24b642cb1037f690a145920577f2cbf7c9a213d2f6d3993cbc43ab31cb55af7fa8553939383e70a68b64911b4ee9eab6829731786a3cb390966e6e6c1c26d942f08575b2cae0520a1b021c92038042d74315edd910af0f9cd7f96d7625410e4b812dabe4ac5d28230;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94f0627db6d25ae69aa625ea731770ef0fd5919af3a117658fcc8f753bf626b7e7fb9fe784218de6663c5f9fd4d08a33264de4d04988e3411779a8d0d377904dfb91d2cc93309e0e855755ddf8a9e20ef5e40ac79df5a2d7bdb9238904df2080f976ead81dda6e9007;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee261dc487a059c079cb02aadc4eb2c83b2e2c37f95e6fc0e8acc41b7f05f1c42b75bc9b74ed3242ae67da19a47b7b313d82f410b0c1039acf753bfd2f20d92af1d414ea1cb29e56a7a6864123a5ab334fd1277ac58adb2dfd653c18315bf67bebbc881e74743b63c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa8fdcc66079af000666ee3ffa7013f1dec8af50db6cc48370eb11f110c7026e5f2a2ad484f88fe33af97d63e06e7b2f8a5d339ebbe728f73f44fbc0c3a6a28be380c20621e29e5c36f470107eab5dfbc92f44a6eebaa2e0d38a7d04ec8d59bb38c5cf4fed1243a7cc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102b6e5ecef39298560f647005f1b244f3b5fb255b9c8fcd5e85dd27f7ffafa5d60cdea30a969c779c08f6027da9029e101eb6f238b2285b1654e111a8992b38edcd2dcb44c2b1b5044c55220e2e380f022eb1897f1a749790447b9e1e7c8dbb2ef0b3c7090a0a9e590;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a185dac4c56043dc98adf1bd4e1ff879ec43b57f2b7ed019a3d99a0625dad4b4833a609418b69fe573383ee9937c0b9476f9734e05732b7d83f620d78bb644628498126e217e741b46ec2f2e4b417df89cf3942e6f728da033ce35f961b7839fd9cd8085159d5f66ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3e942f565981442057fa96f459046ddc37f56cff6b0244952b77c32b637d781d7477da07bb141c53c03a1db750a0ba2f23c2e0abd7b91b3c594fd4af6c74b215699d9a5b20ec11aa1c5852bdcda0b670bc0123d9681be09a22ba510662e1dd24c27e4b58561c34f56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7aff30aa4460ce7e3223412cf6fbe8839823142ef91aaf8fc4b1d2c98194dd79b482e6f7efaa79fdae754b22f8b2817c3f741e96aeaebd206a48a9fda2527eaafdca49926866bfe63a3f3df580d04c7390c68d30abf639999dde04c357dfaee95ab5d7735f530b64b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18aea65fdd3cbdc4e89aee3ea9e60ddf6769126689c495363ebb7744c7cb49bc9ba02d22d818f4402053a1eb3c90d21a15d8b9cc0517aef7b00a9b0a99206e7082117670b3ff6a890e189f99e2fd5a44fcde877b312594fb05e8571f83cb1412dc2cec2db4591aa0089;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6646f71b6ea6fbdffbbf79aed70847f7d531aeecfd438ca3f9fa3d876b2dd40aafa47a5b7a36b95fb2879cc03f8299f7d2ece56d755abc7fb855dc317ef644ac81364ec046604268672ba293d785605af95db167199ca89b5960aa76eeb6b604fffdda11379fc3c99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cdc4eaa154a680704b13245eb75df9488a16c3ce27d63f05d09ec8fb2d6c4bb22381bb6d191e0d2d8d67c8e7f45775cca1d53bbe1d338e018d0695b26bb902f3974fa57bfe423068da22b53c3bf61b93ffb56e5e548e552f008c0da389c67850fa4634671791e8648f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1278038f6f60628e279fc88f60d68113afec2197397f20e40b1ab2d33f15d068ffd9e93d8003debf306844b63f3347ce73f13c46edc4542938d84b60813bc70ae80dd16765ab39c444cb7cce394782301f57b647558ea48ba727bbaf712b78e46819e250f0691e5e266;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8fee95c61f55f7cb2146d56adf48398f8675aa323815b00d805d4fe2cbc4b561ff2a91d105e22bbbfe8c9370cab0705056ad5956da6a305073e9e8dedfb6528b1c7dcc72fa86c5985b7b43414dfc7dbd0a212b8edef1b08834293a44567eee27abaa8a32ff765e61b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha008e8e81b577296c3d1f71684d0d961ad7034b2995d009058b585145bc3145ad6fcdc487b62b3d321e01666d9eac13b87f51482821ad836c58e986af6acf870aa13041f0a41857fc9ed9f51492e2b5ebb315e5d1b961ae335c005e6c7c73be72b22c4d7b331d563e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd45e78bd9d4cc238b15710468c7c9d4937756e380e68f5026932e3f6ef8382c4449044f84cb6a507374fe22b7aa9beb3f1a1844750d80772774c410da99de3139f1cceff89e9aff8a47d3569461f5d41049f503974a7f102b0b7d2e554f6d79a47dc202c3849c49a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155de6f2693d179eda6d7b351beb7c7eeabeb2660b005206dd4b3ede3599b413f645012765b46cb866e7c99798201575e7044f9fd8796b37129f7e5720743ef00e05cd4856ee4526ecfff2c2c09b02621dc76d9b2b73a8cb764b433897347257daec702098f1e29cfc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa494007bacf29e46ba960c7d4d1224560a3d1ff104b4ca064d8eac5c4807c113736a03641a7f1ee99a02ac3e721ca117120f5167a4cc082c4aad078821daa9b6d846492bafaa289ba6273eae821d0b56582726e80a170550b4661d104ab143824af252818e0204f02;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73677a4803b0b55f8ccac36d3cd12ef8228ac19493d25b75f325457d1a6346d05797395a563c87b9e5b60c5b8dbc945bc61d368de0719dc9bc3cc1eb6e67b0cf600e95cc529c71d920068e62de0a2a77048b788545e24c387a53fb4c65929f01b74163c133fc500a20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122edd6eee2c26076730737b8b0f1371a447bf2031a9339be87ccb06b342e48727e3a35f97b048430d5564e19c7b7df517fc0ec4d4757f2b0b1bf71a4d0c5eff35f33212e57780d04a28e41e6501d9316ac4acdfe23ff487284113b6dc837433d85c48b28284681765;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9b032b12f75b474596e3e5d537fac5a7888204e7fd3dfe92b581013e85669856857ae95dafcff0cc644837ab87c1ef1cfb146ad5bdefd89acc5e92b9b95ac8c2c4440ada89c827627bd2bccb616c937bf2997d328c2caaaf858db995f715e92c565b910875d38eea8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h709196097e196e87903fd10076fa938eeeb8964569fc8398f1109857580549e4576c395f7b0f4b1355361b260986319c70b560dc885f2c17c84ec252b6678d9c54beeba17b41e422bb8482deba50010636e9f44a5a56b21e6878bcbcd4d7c8dc292ece0b1f6f6b21dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171b4d1f6a62816ed011fda2c7ef017966c4b3c6aa6c871b98eb2e936a21f7ab4c36b50a6dfaaca0c31058bd10919d872b4d2d5717bf3309608f20561c467f261f1593b5deea9602c0978f999dced99e55cf7ec6fa9375de1c521c453e9f4474b470a2a10fc4389f7e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194ceb8f974b96394d8a9bfa580f990348786bba7749c8a1a3722f8e6d1c959f548d4892876d772a159abd69afd7cbfae59c52e82f91297cbd48d4b86b9634c4e823abcede72b582a23fdbd41a968658ecac888bc45a5aa2c425a7ad2454abc653bf2d9ac7e539e13d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce141d7a746069995ef2c5ae409cb6e7f93a3d8f473e4a048e5009b63d7d537a3c9a18cd4ff25cf5b8a20c48edb0c9bb337a620691a5e04617fa8ec0fdbff12e22fd29931a26fd8f0a29986eb4b4c4f680bc1d863e5f7ddb33b4a6fd6d9929cdbd48e21ba31ddf2943;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6413cb86f238e9843b9839d247c72110af313ab17d73594604838ef54a93f40cfa213f794ed2b598981c2c557502b858e83befc561042a3a0a88aec2e5967c63169502c521bbe99a53e1b66cc78232acfb60cad33fb440d7c6e251e4192bf92c021313e0882934256;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1222dee213bddc6251efa796e920e0e6a50f326c2247ca87baa25fcb1230c651fc64e86883f1f7d5fe9d72dbb2511ce1e8a926004d38a19fe889ecb2101210477a99daaae7fcb5a34d54cea167385a7362c8aa0a2b159cb410dee001267c192d0d9ad30ea727b829808;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9526daf980666b1ab7f550af3621b95ad534e0b2c24eb86ff7c539d1dd1e0ba4ccb97d9dd1be5951f398e502fa269e184566e2f4ed09a8167a7a7b8c373bc11f76fb5f857410d16a4ec6df19d54ee73ac1b05b814f8e64209d3b93bd51615468466c8a6b9a516e8253;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a3d577e2638fdd0ccd45a5b87713bf98b7bb8a8ad68c9dc03cc740129cdd747f271cd50165f575827a8f162e11595694476b68129ef084a189647a9479b35ff31175fcb57ab6562a5df7ab4922d6734865bfedfe12c0f7bfcf52b3680b91c3904ec7aaf3599acc19d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f6a01835b60a6bd09793bb57c315768f3db358f7a711c67476ee1a63756b740184aaea27f4acde96f911fcc7eee3ac78909ff01ff1cb41f80078c0ce8fdf287f60a83b61631e9cde4f1aabcc1acb51f8c3a8ef09ea184ac9fdb07a39f3a76d76dc05f68952179e539;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1351f6bb40f0ba05b2aa4ac5070c23a58475dc5f8f7a4e1fdec306cfe53840b202fdc05619f8aeef870498fec1ec527083ec638c8cc6eaebe3541eeda4e546bf686c66a80eea36427cad0f87d6fc2adbeb79a34e1c3eee3ddc93299ea2f1df8f6293cb9eb8d32d6a914;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd78fad8b262853c746a26e09967d477891df795e0d28e0143a5bb9c82f437c49fa038cbe1504297cfc9165ce3d47abbf41c4a4dd604b28b840d0f4b6e901d35425f64c0958b3bf34e4d43e4935131b1568992341084cd7e3ad143de922c532a48d3799d9bb7a8aa61;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ef2dccd6ac1cc70214f7ae2970ccdc474a78fa111010ce1460d38595fc6dfd08371851dca5fe950a6224ce74337090c8fe2352e515ad6f993026fd3c4e781965603e2ff687b1ccbd4bd6d3f39066eaeca35ce18d4182d4bb93c08c5523c5ac087f515ac6f2a384a2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd0a9fad253de66e51fee174cc425b9b4811922b7c728c63c60e4105edf730e8dd512e84b41f628aafec3b4cd1917ab61234bed9d965f152aae875160b760b84902287ac9daa3ab8c6f72b948823a0ed81d80d125767961039fe10829ee2254706e4e5f81a3a6c8b06;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a31b7ce24c7708589259bf5dea5275ae0c010cec1bf5574a84f39329f4e9cdf148da088df0feebb094f5cdc74357df044760c5b585022044231132b3a9a3c5c19f288d9b8b12ae1607f77fbd4d657221330f81d0a3a1564a7e41a3286b2d3f094492ce6f3a9afcb28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd2a190c8401b982c1391623d92e95d90ac97ee0e5a6868274e9a23681f1f882e7cad8d877d856bd0dcbd58dd6d94b08a072741f0a6ac984afa4a098ab31f96332afb2dc0ccc7d9c691cab442bccc0d893ec428e2067b71bb3f72a02044f05b2e37a041ca1ae026b26;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7c51ba4489381ce877c42aa4946ea14a0ce36e75b75eb81e7a7c28e528f893dd08d04b5fa3e2c4f6ce10fe15b7a46ad670fc708f67b1fa1652b8b462224dbfff06e111081668c6a7039116170f5aa48cc4065a07935070450942528867fd69ccaa24f10052d1c7f7d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb0cfeafc0f9d8e2a703ea31559688c31636613f3521998e1b0f93db68660d57a63c92c23716ac2a6673c187f035d6a83e46756efcfa67026f585eac27cc35336bf45c1b4f23b08f85650cfe9053dc2691f51369e4899a7d0d8b332fb9822be21ada316c0e3eeee835;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84caa7de5518e12b713a0b56443713321e1f0edeb654ee5183e1197fca25116a4f3e17b925f70af7b41aa2d3fb44dde28886507c5e649fb64e7a4224423101eb3560d6645264c15441f35fcff3c45b9a6f9bce3993c7e24513da39feea51603ac6f45a18bbbcaab154;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151441af08e9e8adabd28f8eef32e82dd62b5e309b35e769e64f402de7b908f60f75e3d380ca550862b088a73e13a99ce3209616eb3d5b6ba2226a5beb03d3eb2a397bd75f1009c81c9e69670f1b51480098dc3b86d424df8b376c5a0d4d68c91f17021007651fcd75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5002f99be1b3ee4adf79fd4084224512da947d3bbdce565c670677e9a7495458b55ffeba1a9a3b42fddb342e283d4342d09ff5a226ca8970fc548214668afe061544b464802a4423c5d485541314f19d86599400e74f237702760c73ba2d7fa6ea01c2a8dcf379ef8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1944ddd9389d5c39dd5b82c2f019dc3a4e8237b3f4b2d946eaae8f603d550c375343fedcb7394a50b191ccf6160fe5aab3dc0b595b0c0d2995c0aa6649a2bdcd1020092c3c9b6e56539f51e31d43c6f780b49193599e9c73f8cc86f5c2724f46c96fac4b0a7e1b0dd60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f7d557b7240a9c13697626b2da45b1ffeba04da23eb7968dc6e36e4a7085af27828a69042282523660e91a34ec2e8c024d9b07cf02bb8a7d9379790fda7948509f71b1498a336e35bb2892f2a655530996435d8a4c900b9569d9705782a718b6050bf15b81e25e9ec;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80ee6135808b5b39b450c63501858ee9d5f00be394db266c80e6344f5e5718d322aa5a2e62ab650d710f39f517f95f68d2056d92c2d334c2657e7a84ef614f34e0d5f0cf5532c13db0e6ea0b3cdec244986daa5f43641629358d1de17b866f98bd4b85eb985cfe9f0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf076d212f417ede34ef1a3c60c2755fdce6b2726e391106f259f0660c93dc038b4a5a5f0fab6eb8b9d4004ac042b0214fc3848dd43338c3d769e686359249f9b5fe738210f4130ff3efd2a8dc59c496a35abcf1362f6d4726027b024b552e3b03d54a25a043994ea1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17178c3edb9a8ef659fb4bd1dae04c6dec94f689c6d2119c0df4b8bf7cdfa9b6843009fad6a8e1deb0beabddc736ae5ac716cc402a6938c8759eae86022c9e85ecf0ca5986e33757c75972bca100f7bfa1e906b219784eaf0820851f1be1dfa3f36da7e31b432303df3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbc5537a758de1c5c911ae3d6e6dd6e9a3d1cefdaa57cfdf027e44184ff183774b09a86688ea19fc4080fd5394a7b8aeae5405edf733683d64f2f5059a05ebcb412b0ea77c14d8cc6fd3f42171b3f813ef0f7b3e8673b7b297b837c0c9eb15e5219fce8b933ab34f4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1389fc414035dcfed634ec5921e264500187199c4c2483b4b8c409b8937ee3f281d18e0c17a143118cbd0816809565624dde4cf12a5d29ced482eca7f86dd68d02694ce6017b95326fab277557324d6828e55c809b24a28359a34e5a33e1c438daaf0a652ca52c139f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18cb7332ed26fdb68139fee531a539b06f684a926578c0b00ef3d7fc44fd116b2267d32addd25681667ca108e473d6c972d1f9c891b729d29746e068807338d6f587fcac108bad3b2d2f634f800146b2c380879dfe4bc3455e7e6bdbca62b4a56d87f0d2cd2eff4514d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0f86a63b5cfa9031606d04089498dd92beb115913307f6f61b7315949bf9e58a99a010fcbae15e759583df1e5adb02e8a8770420fbec45e23de6561646733a56384eefc3f7d1625f7c6ade9a4551f7e99480076955f3aa271aaf9b8952c2aeb5d27ff0c226ba99793;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8315942d0da90ff2f43b97da97862dea1a251084b55b2962222eb4ded072a2f856812c3bbb420c12ce1c0072b1797dd1c27d3b60f7c61b401edc1ebfe6d13c6d48cd2ecdfeb7ef55b4be06ddf7eab418f5199d79ef403ff18f0760d13fda6b01192db93350037ccc6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1efb70cb5d22341569d269e5486331c16e9f52c260cb0637c1ac06743de38042f87638b219739746e10e67e20111b01289bfca151bf3fc7c5dd7f9a961ef63549f8a95d02edd4a6e9d72a669f303f8449b1a0b5b527597131c2fba1d45348e0dafc29542a03bf25143;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2154fe4f22d0f26d479f0ad40adda11983b8969f25de43a30a05db62b5193049ec20e557215372c684bac5310337cadd1bea7d0cfa83a1eb8ba43395c301337ed17b5b41f86c937a689e53773082e954ba60f0ed048b5f980d6acf1ba5faeb99a877b51316646e1c72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181a4ef6e043607ed4e0e124012605bae8662787d3d653959b248693d743a2edf687aba6ef31238557c3ae31ee64b70b0af201e01d93bf86b85821890453ec87b7f3ca778a0a689081887c31937c8f5704b56c31efe71844cb550aaac01694e72b1c1630598463ab052;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c8aa7c4d7cd8749b4f26daf7ce643e605abd6803bb89ae76777aedb3b3bf20d417f7812c2580a1a3e17ff6ee3f9dc415b312f6d4e38603c419ef0a9d86980a3471b8fbd2c4559bd6e613fae6bb98d28bf8a8076b8c83ebead583ea129829bd6dd96628c62ffd104ccc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5052c69a5438b0f2707707577879f4b7a70dd0222db9696ee37ebee18632a3bcb4083c554d2969bceea3926f9662bfe6102943d6d9b95e6748d3dbd72aefb5e5909a02eb6b563885ac56ba6e26cf93f781db3187468fcdac99fb0410c3c3f0ae8549407cf9b0ab6d74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1983daaaf58e80a54e5dd259be75680193a55fceca86ca86e67edd49abf9571c9830f2bd227e2d447f1e7759b246c959ca9dbe7ed1866568ea2d235aa6bd11413c9825849aac016bd5297f18de774a7d52bcc3bb0ef2a1f41264438a818f809755904559a0af93477;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40c141870e5dd6b83986dcf4faf6f01b2d466aff794eeff334e4a4ec4ddcd2a557b91cbb88f062be776959a62dd4a5629c428c79cf507d8e20e450de0bf70811a9a14c39c5084ad9cbcf7d11a592489555c72d23f3a40a956cd312032b105dbf3396120f08c41be968;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha322afe4767b2428659088700a741052c6d1f0eb37af096c8f9c34faa1ff8c6c1029fa7536a7f0d0cfd088ddf32f3902167c977b95d422477809255d1d9aba305157b4dbbc91d3427c887c57d04999e1cd12eaf4b88ed5855521510b9c86b2af8140bf61fae7645457;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13337d92ddb17471ae57937b25685890c89c4bbb98c43f5109fdcf6019062b7618d20ab29d647e43e3e2d9e6c4359798341ae91441f4b9e28579fedce6ed0ed7de45d45b326f41f8dd96a14c7aab3461b0e86994404feb695a4b56cffda64bc30a4afba2d45ee7e8220;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6378de9d072e1c0187dee70e61c31d334ee3799b9de6f160284fe66946daf010709eb90d79ed1b2770ff198488add5ecaa624f61cf38be62bed80e292a7ccc60560336afebeb1ffab8e7386216fc26833095aca09f7913b2b40de0e698aad6b88879ab7cbe5a2e681f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe534e196c34c1c2f3de813a0a9fe5528c2cacbe5cd0c31238f45d13dad05da53fb93ad78165b489ea12ca6efdf63e91db6e8997178f9f5f664fa9f7188b12092d5156b8699f5f37ac251a21512486bc6b7336851d936e310d0fdf485934f9e9749f23e54538dd7e7c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50ca31cb6f113267d9214866152a618eadd49da4f253a65d4be2991429e66d36236ea6026a61246f13344c6e5c2e1cac5dec71d9a9389be35924f9109d3f013b58d9b1f5d44a27b6dfb81783e204528ddadb44f72983032b54e144ebbd1def9348a991ada116ad4564;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15689e36bcaa8bc1f68b8750c2d75101a1cde6f4a2cf6ffd61841734b0ef48e486932cd0d7c7c7bdfc11c910f5f4bde5d071ef134d9d90b5faef50062e86b2874f9f92753c6ccdf6ad2b5539aa98cf6505befcdf4fad00f310e441f825fb12b054d5151d12b0ad2583b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193b6ae7b761cf681298f65e0109b2071d66cb3aa7e35f99269bb58368ef8dfe4dfc20dc45c2468e11714e3d8a77750b6497b92c47849618ee32acd8fa31a760cbef3db917800ff76f9aa9552998ef1c674661ce5f01d2fde919efffbf20ea08a2f4ed4447e9483d7e0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a931219524c5b79776ee93d1eb31e4146e63dbc5d132f86f1319534cc99a47e42e08e692d09530a9dd9ebeb8567add31414ee95cbc31697aa2814cf628751cee37ee8d0d984e0a88257dc43e040778c3b42677f3fe77d1a4c2842ff0b2c7c34f06ce4591482af7d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ad56eeb082d63aafa79501e6abf24f25da4a49b3adff9b986b365f539939a8b678dc9bc1cd39bd35e7389057461d3aa93849d12e531a0db0ace676a2c0acb3ed10ab8cb4162a20228523565b72212a69a31035b5505858b7bd5d5757b0b2fd217ed2819dfa3fc841;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he60bcfab4a176dc65547f3d3307eaa78c741a0de252317f28819e839b45d046de89ce1f479cdb25b117867ea70c276847f5d39e10ee9b21d5ee51ab2a4e2343d1966f073e4de4025651bfeab82c4d271f0991e6070d8e9b8571fe3e37b06aad799e863241c3203914d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h392fbd7a161b29660eecb9aee00127b2c43a7d478d6cf2b901ddda06b2d572efe036a3d7467a75cdb8d94dd6f53c3e780ed7c8259aa469d629d3b1d50be2ad6629e5924786b5d5f4e5566422796330ebbe4e8053babc9a6c38c7c5a2b007f632c3037900b5501d190d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc3bc1062d06a119536760fe7393855f4c673de87047f5e28d56d295c0877468b35323f9a1b9126a3141e086e3e56a37f41716e25098d021f3a1939abded77e47fa052770f545503ed17ca3d846998d06f15a0806570205168a7ae1406bef2bc3d6897fbdd777aad0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cda2590f2035049781bd573bb217177a6f2a92ac8bebf23905987c9ec972e7b2d5bc56a8db75283fd939eea1d439b4029edd7c996d435f9edce067033a14967fc025dc98b2c40fc836d7a9cbf570c958330c7b121d3a17d5c5d3db7cc1584f0dd043d61ffbc5b303b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1449371cd1fb5d80231c335fffa76e7e75f5c1943779461e348907a96e4b6a59ca77a455bc49dedc2385154e09fb8cba8e06aeb1a02931aa2dd8289fa8af30b1f2334dfaeac3e9ee97021f19c58f9bc708073ddd4d456b8db79cb1ce7b22da995aba80f54d80e1bc134;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h693b8d0fea12df339cf813a2194644b4b71bfbe5e463c77e5a2e8c2a0d7a2abf1e9fce3492ba84dc041df0aae1dd02a6a9cdc8103b33adf8a8113d14ea9a7ebded8a9d9beb4f1108d02a6fd44cc4926452cfcfbf7ad6123508adecf73bb0e608cf873377ee6559c238;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a86d672199bfcfc5bbc829dd3ffd312a6d024506b69968651542892e30a49402d38432abe7b157b9ad767a92e0f27d5e9605cdf64439f91d262654dba4f82f200c1b28dd84208562647fca7a34d929b6a60aa569c6f7162d128d0b94770e431202810337fb35983f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85d8b3f593e4fe6fb0ce569d2f3371b5046c8ba39585e13d7249bb3e664fa055827e9c5ceca644703c1ec376b40f95464098bc7c810e019823e525611a3fe0667b9092466853830e2f4069a3f7b5f05cac79a56435abb92048e0dcf4ca472a331be300abf1575ebd31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c1d2c2f98dd16c8f38a726d42d0a9671758ca6e39bbb3551a00071725ddd7c22e8b871b18c55ab23131f19db4c7a37bdc062fdeb66dce091607474442367c07d3f97ae2c11a2f488d1b2fca281ac4b8195798ef76d0a2bf266a488964d832cb73eb4982277613a2f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdce50e3639d4411c9f68a103a6b17d213c77324c6ef4e77b2db8e53e6bef9eca09be936b82cb21e24f207289a65b7808e6d29166b365fc3b7f2c7169ca32d9864b3bca4d96a240fc0af69dcbf19f8752592a6180cf95ce89352afa751246b47fec5dec7eeb81fd4f9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7235b3ac57239afd3af222f4a6d28d5981eeab65da25d707029add3c7c91b5d9fc8b1b906830fe1be6eab77e3b5c97c754e24e7458d9fb896169926db6f04ef2e5ae7bac26e68d106254b0ee4d86767f3e41d93656fd8cb4648c37fa0546f5453691b27796373b210;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h985f56045b0f20d5a24913852a2ce1ed10bc120c373c88d092e71e9c0867939368aaa0f377e62c77f1dfbe33cf4c0f8b4ae1ef198865da9135f298b1c66e7551dab449453887ea494fa3ee35b6004500fa19e3ba09c0c137569cb1ee6f54c07d72acd0e81d8e48282a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb537c3c3afea3fc5ae0e0bbab3b9df77c43ebb28e65af001dec2f2e4f726b5422cbb2c47327179c0d47424dcf96ae0cdf25406fdb06183a1cb43eb3becc5b1855208a47e479950ffa9862e42a72eaa83a0aa4420d84b428210e0ae43aa216e302ec736a4671ffb050d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h307ddb8524b2646c1b153d414c8567a8ace06c8979605d24d57a77c97b2979cfc3625f644bb773b5bd2a0e6aad725dd078576dd5d5d3f93e888775bf85befed0655c642a119e366060af835ec8f9a9ac8d413d8f30a8cfa4a9ee09998892b52828036f7f8155c66738;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79e7e196923dc361fe3a3ef6f3bbda780b348892ccb693ed787570e3d26cb2e55a46f2cee7ba16691046cc3f7eddd8a8c8fbe23f12d5a4d391342b6d2870dcfc11e7ef61490dc7ef8c41e833bef44f7dd7b4be036ba2be9a2b31b0bb3ef971167c1db2ef81ab3b3135;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42289f93fb2f60b47337574e07d419a9be691389af08f1ac69b0c443336da368fc6ca0f404d37b1bfd0b896bea4beb94112b01e7530c5dec182c1d09c5d7884bfa4c753b57b291e289fc86ec5d02bd90dde8d32e0a720fd656dd8f1435bfa0c2b2b9c8d760303f055c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1908adec0a38299649bac48c3a6ab8f79b40366ca30713ae4add086b10d5cd51155ba310615618e17e44c17a77f52f98f2d1913f39fc6072d67ab3b728c8f15790cf35f7add8e21ef806c9339a0187ed40b0ee359d53e74abce110352164d8c36711a6045defaf742ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144055035db4dcbc8d250e31b6730e5f35071fcecfea3b125206075a729f6b5253c39b88408878beb51d3b5d34784808f2385b8b436b449f1ab2e79a74418c0b267bd57ab322369deeeb9784e08a94b80c37873dea35f9ea4b0eb0d3163769959eaffe73a4ecb47e9a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36c42a13b98d03c291cc3a8c67b92cc0e2b3ad5b42308d4c1c4505d858d1188b5de28230830de46798ccd18b247497384513f0c5551126dc029fb6cba08d5bc19eade1e49cccd18951db7d7961c04ac258a0589da19d96eccea8aaa7d49b9d000cd646a2d8c6930992;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5b4d10a239d8be568931937b0b36c0a3d28874971c9f1b4e1c691b6be0b937ae8785ce562279f0947ea944eab1e0f532a029edff9e4233ada1fafc17d7b860ada859a58151a24d27a5bfaf49148ab49f2257ae6ce0cc15c56a6d8cce7bd1ab7316f56c8e324c7333b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5138b80875b728dd4260c6f688c53ea22a7449bfeb6e0ad2d5f52ace5563922867875726fac0049ff7997b9b212bb4e30fb054c281b052752ab5f8e6309cb69652c19c71ed6f3d7f878e284f36528b04026ecfd8d43dd57a8a94266c8db5b937466c029d6ea84f7a9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c52e42d059b1e4a62467fbe391db4711b5edca3fd2c425b638746439ef01e56b5b3a696c3d5c6a06b5fcf3a7e27005713a5f8d1bb99b80dd7e79ef29ec04ebe20208e5a4268ef39269e112a34bf23813576d5394d0127c917311f6146e4a95ff2d275f896ab31b72d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6cc96bd97af05c00abe1b08a7e7d3862676d69d6f7a6b20d3dc59da38994c579f27d4356fc1d96889bf1a7ab55db226dd9ee18793112595dd7c1b63b7446a00ca333bc6b5708fd924403baf4a8b2c07616fba604d9c7ee77e576621e1cd1d22ab04619ce92d6752b21;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3fc7276156686d72809554134c86014abb0a14648a1bc45df2f332c5648bd65014f1e04778cf01871ea1f00fa626dfe2e4a1086cab4026e565f372fe5ea0e58517abbecad201c30492cbd613b51e500a230642a86e239d517fa998793330a0066d1a775e97311304f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10972f4834a051f91f29644953706879236fdfb236888fae7a56407109a561aa555646191df304ef6d9879c01f83e9800302cbaca24e98de44099fc6fd226a2e7bd0b8fedd7bcec8f9d81627a58e086ebcb3b291be86b7eb9191d738a86701a224dcd1f1333e0cf231f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107959824cbfa5201cd99ba07745bd547be557b9217676b780e018c5b67f3efc87c3b629738ab18bd95a169402e0434dc3dcad30a26d13d21809662f4e3cef7a3b5e524e286b1708755688f366ad5ed54ed1c84c9ff87b51437f25fe307e342ef6cba22a12a9a5413c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h761a2e062f85e8dda84d73b3d520ebcc40dd202e2b8eeb1357ab3c8066de0826a6a4eaff3dafb10f78d9dd7a732f3d63548e2b4348dc6d7a2f9d0f246ffe8f19477080c945e236b347a346dbe5f2d1f34f3af689da4a168e421b81efb2a0361f2b69e1b31c45e483c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12822cac9f321033653c3ec80396fa37b56ffa2ddf6fc41f65e5287003e47e884972ea3c77b29afe644a64e39d769e8ffaa6972519e448291c4e07d5f2f52d205dfad25df7fab1eaa97234678916ebe9edac3e3c62abb1c81e35006bd0bc2dc28a6410847c3e388b2ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84c61e658e5815cf9ecb9a3877b3ee4cb0f0895a5d2a997d15f61875ab5319bfa440c62596a6c980f959a2efa40e713e973bd0f1f4654081e726aaa25e66b0b25f2efd7ba6ba6d5191e855bf837491097c65241198649e6a2fc3fa5e31f62354751ac92362a99db35e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf165f51076121416e47eeaffdd4f08d1fe8ad335b1c4e182b893ee5a41d46f644b7afe44ae913b48844792cb588025dfb957cfd1cdbbaa52dc295f7f73b6c65585476811a5df4c384ccb7a91f70116051bebd614de242b790320107bb8df5954a8bbaef8ed377c60d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7637c17f820aec80a0418cc477e9eecdd854f8cb27824383fcfaa06950d218122c62e034fe02fc2825203c0c35ad52effc14eb4ed9a76c34c2fc5901cd313a1359c71dbf1d1bdeac6e534ed992dcd31cb73f1c24f5c6ed2eb3e1ce8c6261a8762577516498f2542d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b542c947915aab5ac37acd082e9bedf8edf757dd6eabe21086d15d74d81dcbe7b94d69086c18f9f9ba8135c7011ea78b7d18f2b00d717f731d43ad806248149910f77236aa822df59d4a5966c7909595e0fd2b7456666d141fafe859068057cb7eeba5ce511f46117;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ba26df9793f754b7df8955b74dc137f12dfde1a0616ccf8bbd3fc8c5170051beeaa4f4061f63d858b9341469c847de71aaf8ed6f0561b34104cac02ba5b55bd6bd071a8f8876ade85a7783bcee2008e51033a35d5793c6d50cb39f2abfd0f59e3081f6e3506cab591;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda8bf792dc7bcd14c0ecc4fbb633e1147a0cf2df51dd14ec4ed8a342d7644550bdd674dd8c7cc3d7c3eb0ac5bc7d82a197c01e2235a92aa4c3a8aad9d2aeb8b1639c276323a7ba654c377a1827165af642f1e72a4f8bd8f3495d10ccdee898cd5829c3047cc3dd58a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4ba2bfc152cc645a9a9b2b3c0a824fcbc68a0c8c9e872fd34c6f8988499b7ddd76c9c15ee4063b54ffdeaef4bdb55957149233e95d1863039a9dda4cd3d8f2a2a48acd3c072ce30b8ae22a09d2dd5cc062d0c327dabab89ae35fa98729c6e2b092ebaa376b88faa97;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e378c6dc2cce20ccd5bf8f2df8f5e96ea75a8e2f6cfbe0ac44aad93a8341496f34d50f5c6d8735ad1cd859e0099bf22c9b795ad77bfdbd9e75e952afa69cfbad832586812d63224378dda2a66e32b38765ecfda9065e9d467e50e73ff1fbbf2931610e8da17537c25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e3f4fd56b6124a98bd1fe92f004dff94b5eec2e47d702b945596bf093355824bb6d9519faf28752bc4f14f5431666deeaa4f0349bd7a4b0ce32bf64e64ec009f57b7cb9db54a8ffaaafa18544bd7a9093fede57310524aaf3cc0f748f8daa7a2d4362bf2bc4a070af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4275050882b0001fbcc58f524d32e8ef0d72048be24add44336104b68667508aeec762cb5f231db5a0f4d9b1c18d5aa80bc201f059cff55d001a08e10a29a5eddfb8c3f33337f4a5ad3aa5cb59818d0259b197fe8157eb4354fa3d7ce0400b35f5dcaafef01e8c6dbb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e9b05b22dc4223d9f1ab03dbc72c17601d59e84eb288d2940a71e4ce1dbcfbd34a35019f7527b7795992a6718a60d6d450510712dd03ad63f91c0084bfcbf4d17f6f4beaf6878bf78397e70817c832f5e5353200087c21adfa84348c2b5abd1a7bd586a301af23254;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140718f9a72085d2258b373d7ea244298654def922d5db421bea9604afeb7b4379c1aa7886fb5bc8d02bb38ea209251085b03ee559ff77bae9d81f953bf66ce6f367a92f8dda855406474f56af8ce0a89c6d0fef391b5f950283daa8cdc46a895113447c09302813385;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bde361eb2d1bf50d2ed17f5191fe1d136eaacc51bda57edd5500abf28a17f96baa758ad506c67837bda0b323eebdf82fd726fa7bde168349abbce4771553f6c8a7283077ffd2681b7403d5631bca00b37869e20523b2339cfe74331d2d04a0881903084e848534136a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h589e7868044ec06e29b9f1fbd70dd35e1920ac66283a50dba94de1a495077ae0b9faf79fabcdab868923d9e535cf3adfe8fd43b70b214ac86083b9b432862f5467a0cdc12d82dd2986bcb130131224fe3425c78e42ec7f1fdfbe17a9ffb4396b7b294d02a8e019b05b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fa8170ce5cd25299c9b87d9664874a26211df229f145a73232e0550d37449c266c63ed936b048dfef8a239f8083594f38517c66ebe9bd844e54724a3745e3e1a7f00da3e3554f42faeb21ba7f635be599e0b579e7404b38e46d83516d9ed64003f74adfedda2abae1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6689c61cf20030ee471d71b7af60d408b8c53f5d22e3acd668965e18a078f6c4e9d4839aab4efd51bf156db7edd617bf4c86d0b4eaa961dfe65d6ad5be4c245a19d0a09f16f00234c0d5cfbc49e6cba248baef5b6c90a4d1f73165d3124cac4fb4b78713d5aee2e350;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f9dcedcdc3d70e17a39e0bd018308199f905a835367ac6554c0ec17df582bcd2e00fe0db727197ab0ee6cff7f890b9b37162ce440821dc8361c44b040ccd5b67ac6920ccd35d39e711845f5f577ce962a912bc63f594fa05b1477f863b415ed3de144605e5bca26ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5e71b73fe027b143091fdeb6ef96c9fad98f1cefe53181a7b46b4846979ed39a7990a9f55a60ed09b0cea7dab4bcc4ed2f7f164de718ac9f0962491d7d27ebfdd8260c2fc4d3620f3bd532f3de51ce7ad56e0ea55d906c02af5512969459768635d5e746a47c8a09e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169cedd4319440a8a5d5efd110925d104565af5ff12b73cac341d0f466b16b85fd712828a022db0a83582dc83737520383e26eca43896ed94262bdc2b9db909b3e26a284e2fd3efa63039df402b0f8eb9b87bfaf30b856772ad09fd2d0d236bcccc983695f132ac83b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4ce2157f65c8c0f4957c67616e6b48abde8aac2ce1bbd1d6ecfebc9db5f26c989893ff631aba843697b563c43589afd3792f31fa14fbf986c77f523ccc270cff607fa1e2b2448d6231577ddfbea97da44af3443d6e9e37d45b27b8b87e3c3dd3b248161970366fc9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5036e5321928e88bacbe47190c857af24f1cc422b2d286bf78323af868c8b4b12f9f2e0be9b7ea5d29cc390c38507b0f89f388e6ff505b5cbc4788172ed305357a0565a56aac4c26c85991b42b2a88914b17f6c4c2f9bd16513c5b353b6efd7bf6a77736762261d6a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1668235e511e4f32738bddc55c3e214763c550a684a5a8800827820c0aa71b364a10ad4f1ce55b8a27a4f20a8a4e4f61972e5de95f0234cdaeefeaf817afa9d5d3375c4f29f63b0ae66084300ac41d46dd758d8c578b1a424100cfc057e45a8163b547b89575fa8e924;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1409f1fd406226e81d24ca617f7fd3b10f6841833c40b602c3de4517f9376bad7c8da3b4ca71ac72ca58d0d6037028d58ace3ad7b8816953cc7d6282cd28e09676c1707b5df73fa6f45d63583cffb14854f4b9af81db54c9ed70277371470e423588279597722395af6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1505d5a113afe4d19d4b1e4f19ad8e0dfc28cf5b45446716a4ce6adcbfa6fec5115dae943010b54370113f52b97fb2732fbe9d7dbf9df9c675497c7e2f8bc57068cbd5e35833e9175007c1947e28e43637a507e0ce2460b1ac7c1a4a7b04be424b782f0f1f688569;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h97394b1c3e619e85f6c77cad21c26659f8049ba12fa17f3a3c15f65f3590254ed63612847c208ec7716ecabe40c2197ed87fc043326de1dcc446cebe21710a6208894dfa44c3d4b073b42738c50770698e96ce9b7cfcbe13e624e2a042b092f4e1cd1459c1cd02ec67;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed5b5944084f83e13c8938d6c360a8078ad9725a5e2ebddbc6772d5d6db2f53d485b03461f54348843c4e91fc0c84603762d8ed471ca7a21c96bdfa8640ec976fffdaa93637a0fef5ce576f49ebd4958fbeab4bf5078d32d6dafa332236a7a214453c609be2c4c5091;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51f7c16ae3b52b8372e950ffa840aaa92503fb3495d698d33b5bb1e024585e969a2362d35b9c295e9eab640704643aa69f61f6350b8b5aa820a2b9676f24a32f2a7b61af7d6a1413cbe8fbd60eb9d811272223a96d97a60e679ceb30c970b885709a98facb6a4cf86d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ab02c6743bf79278b0b401fa614f732009ab1d3bff424977ae00eed529749e02296b115d947562e8323bd2568819df52c49ebf49954cf9740165977c773351676d89fe58eeeb50330abd50d7d93af445f9c1687e613e5e9e9af0d75c5f9be487a64c90e017a11b842;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf332755466b494d785a834ed58591a3008a6a5ae8a9a0d00f626cbabfe2fa975c65206d797ed3b4e0abf6cfdf7272a41f5d2a1fbc0edb1a39b42eb6fb0fd08327f01800d5cab868e98c6ceb7b162ae78b371ef769cd7b1f1269fb0a9a220795d1b0690d2f30e5f6e00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad6d9e60f7ac4103e206ee3edff78b538ec922d0674bcdd02670264b4524aede06b5d06d2282cbcf6a6ed1e0a570e10af9e68fd2cacf5f82348934a7993bcb66adde6c0869675b3ae606e37355c94c254d5054b7ac197f766f743651ed76969fb5c827c4682f5d38f6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1a67ad8175fcffd94a1552db084d31f523823626ad70a96554b0808f40e64cfc1fff7d1d7c7cf559260248d3b293dbf4d2eb6b912131f61c49a5d816b4834715d19f2512e8652ac4cb25009cb0ce7d29557b5c6f55489f3c85b5f309b2e11b2746f97e2aa564eec89;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0c9bdae43724f93923d2a672073b82cadb6846190587a8515b571afec15ab59dffbf34909d854c6f72a7652f0803230f3564b7effcd8b18bb91ad3658db05b5b12f0ee88462ea8cf45c12747cea764cdca0709dfc03fc86997b582895d73349e5a9cc0029d3cbccdc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e735cf25e2b8f5c329edb9a4ccd84fd9a78692e03707264c68811be8154e0755af71f73a6322b018b09ac0d09dc453781115fb752d4501caf72016d95c387a81ecd10b7b4a2debc4448920c2bce97515376c2bc494b44620e406cee75ab4fc0b73986868a863c612b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c3b2894493b8f44054aac7869a6b7fefe79f41c2caaf3cd204ef81c3c6832daf88a0c4d65165b12106985b50d914eb8112711ea56fa5dca88d9ad3bd106b9d69e5412935a53a144016caa843509d95b4276dfd712278f2a45054715ab482dadac37871e312c5068dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5381e2d8e746f0c859260e3a267612a638ca4675cc4e70c1010855f9be9c13fcbed5b9b5a9ef6100b33f20486ef658f95e2720fd42a0058cfcf11407d1fe5405e4373e661bc467b8cb54fbe3d8567550ef1bf17c0598ba4111323497e9c5cdfcea4e44e54bd8639d30;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb34c5584f0be95b162c20f066037d541ef7a054c1e15bcfeba42f3560d803ad19e0f47bc9ee9d10e11430f2f3dd09e18151e73b7fd75610b17a68ed1956b58e79ae503f02ba09de31aed3acee615dc715c60125beebaacc8d7d6c4d50f570062a2d853fd1d9e0e2a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bf4c1a05ccfb188e218e5253b2dd3253b40734f7a825471a7f1269a67f9e3b5b1f5a71a2da3f536765b3813f7272eee1d4e67ed7f7f9fc0abd457047c3ba29781d6fb53da94f93c2342c609bd0562e41534a75fd9cecfe74b38608877a0b349e2122a8fbcd750f1e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c8b0f38af3a4ffe98ea2cb1d32775635b2a71b8d7c6a41f0bab014d9c4c1413c50dd747d138af098c94d8b5ed260764e98272ef4d372788ed33e60a6a5daaae0513fa7f186c2f547c7010f38255909d861b325ca5ba32399986663786e866194fd639d49a231102e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1083e0b1313dcec4fcb36ea6ef3be22b85b64dcaee724f7679ff9f46c39d82f4f9e8d12aecebb2a0feb00e6f04f9e87ec4fe3b691385a55dc5ce2b21fd1c9a6cfa7b1fc5f728a2e4d175b210c8643af9355a8c5399ee0c8634a76453812ce7f2a1b83c29ed7903a9c22;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6222488221aebcb5fa93a3e9676f6e15225df6c637d1752782bc17d569e8e68d0cd4884ae06d4f8aadc1df92eb01bc504fe1ba1ce97e0fefd57dc7cce71525b7b8747eff637d8f0bf846336c9c7246d990bfc51827633348b115d09fcb1ba0a05e479f630d3050d90e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109002903d4adca4d3083f47532286738c00cec64f9cc29fc47661688fe30766cc94a2d5b1764f6b9af65970ad511a96032991e4ba45a153a71e257987b5c2586955e2c5db6f891f142d1dd1fda0a7827a4a74ac2007d9362a8bd24e1ca3e82de38359dea000b9dd4ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25f28e18d6a52bd50bf1229d1ce0db726c05f98d78a5ab2c514e0f2e9580cad29ca67a798cf1f567526332a6c96b609845291c948c0eb1e344490848a71900be773ad5cd0362227568002c57d69b7a75b38e8cc96491661826259ddc2ee7d351e652c6b392a07ce3b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a080036525f3a6209aee026221ce87f3f2e60f67505991dfe030cf5704212c30d86c093050fcf4d768b71290484b6b4ee88d0a1cede94d8c1b10b47e74e94064b1dc9edf3463cd38bba254c34252675b8770c25d26babb3a943a02be9751556e4ce139ee8561b1b65a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h455b93d3f1301c2361ab019bf131fa3f0813fa2ce2f9f03f5d7e278f80bd4ebf6dd4d9b091113b8de0295e05b07e9d3d2c6144af2bd4c4eebe4e8801ee4408b8c96572645f08bd73f235ca2ba672e66883ebc0dfd422ba86f42b29e0f10ccd3bfeab0fd2ba65cc2bb6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12250066a4297d78c5cf8f082e2db978dea0766b7005e2d10c4498c8a58a07200b46522914effbbe903f5a5900e3afddeab1c5ae8e510e22ef4b5f0176a4369051dad9fd45f0a384dfd776b2aaa56c5185ece206eab3b379f0d4c5db8a8c61786196eca05072b10c628;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19282353d55754bf406c5e849f2adc34a753b0d398715f4c4626e4d4188cc5384fa5c0b422010ff54b3e7b4b44fc8739290dc749390c547095b7efcd2098b2e11c04dcf6b75ef0535dcd0aaa940a1b959e894f138562f507ddd1e1ed0241f4914e8639bc20bd34118fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b2368320a21a866475f4609f84b02652aa43dd55413d7601caeb159ab7a02f70835cdb93324e12dd024c3c728f7d800e00e685106610eef3b7a87e6258c23958de8003135632056f9cde1ac6261b56908185e31d1351eeb85a5a3a64f61273c674c2ba246311f091c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha844e0496e6487d5a9d8f808aed38af7339e7a3c2c416245a0c6f39b8871c634a56306738416f684850026300bb35905f3c57e69694d2d234ef7697e7d065aa516e2ac90de6b60b30274a0528e024070c5209e506194a2085f94338490389e0add24310c28fdb9c3c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191285ae3af8e9155eee0e1f5002bcc9c71251c64a071509a5dfffbd2eb032729f874213ed360cec5685b6f64041245ea4db3771ab07ac6d6eb29f8f4d5546852d1829d6596b1b43d16d4a4ad35e35894bfc75fabca5cb8d7775b98166ee13b007ff4b185d4393c7d6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffab41cf500bd3025a94d57acf60b2a0f95165b9d21442de524e9b6441ca685c8a9f883647ae283bbddc0033b0ce1fecdf9888f33c310487770c9aab56c33c76ffc8fefe7f44ec059c6ac9ae6a544ce5f5d68a769b9b371fa53b8b5525567d0b0c83321461e42946ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4957fdcacbb2e3ddda74e374e03a7c7bc6eb64b8629ade477b26ae9f9605f4d1e9a02de0146581dad8bb9f7849d9923d345a7e787400d8438719e8806ac549e10d77e3e4400d19591d0fb59c26ed8c13028eb13b1a8957a587d6cf0ca5ac90c0c42b41fd41208e420;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100dbcf203cfabbeac407fd0617aa60aff89220991b68e12b0443cb5b852ebdaedd5087580f8f9aea11843c9121e1bb0a2124fb88dfe7784d3253754c7a0c6bb98c4842d4685612610e1a7625ce7f4fc966e9b317141a422b0b644ba0bb44ecc34ebaf6f5e6445642f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8e3076248df15b517c2c7c4ccac9cc7977eae122b0d823a2d0f32d48ae11a77ce39dc1253a45030240130fc4087d071a4a67cb6ac5fc78dff9b8c81df526ae735179e59f759234231c3b898ece52075ff1a4e1489810a87a22f9dca0de567201842933b39786e58c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c334246e40734a7bd953c6e6cbaac0ed7e4576f38df8288a87aec708b83905a56061cb4a9f84e29521b9f72490a6feceb8bf324886c43dd1a242b69ce905f906f30bf30376ec90d29dfd613d347cfd8a6e7f9f7a42012ed34fcfd88b8122708806ac192c7717cca1d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc6633770d1eb0d312726af94cc5591ce40503526238990fa6ed313b8b280b2af93156c37576e9fc1ad9c68c47659a5ccc0f2914352ea8083752883bccdecc2feb82184eea013bfb81732fb3d2360c3660ead2e7a1dec2fc32590f594925c2e3af14f96802b73b33fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c407eec8ab4d2d643d7ca0d07cfbf58a273854334ad015c7aaee9902e38fafbe29ffdba6d965fd6ab64a5f8708582311855b07f28006fee9ad6bf34c38ca2c3292c1fc08ddb4b2224053743759ac7fb9480d8fb1d4f16155cc56a1f99a90fafd4d27ef931e2373621;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff2fb5453e71b975ad0bdc6f78ff47946b5d06a62ac1ea178156efbd572413c9cd1bb0eea4ed7641cd3ecd61d35f5581b8c6b3645d26806bcd09ea5cfd5090dfd2fa7a94c6dba45266f955f0d8c7fd5e790779e4efc6e2cea5db892af5870246dc3d0eb40165c42bbe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be61282d6344623f27365316d947a6dd54f94b74514ef9f056b88767402d9cad47ab3472a8e9ce50e552959ab39105d9dbec664ae8b648a340f796d37a976fdea84b2fcd52b216dc47c608c1c420834991a144a1a7eee05882b64b288d6d079323d342a2a3c3880b4e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3312bccbd84caf3030493197e30a42fed35e491e024ebe58ff6ace9d144e407d9000dbfd555a2ea17a8e120f55a3ad971970bac917b3e810db52c95e7feb381e6fe0245b0a2a2b080ce0d6a3f99fb42e8c647e065fb9ad1d72bf1877960b1a565bc7fbf1765ed8fc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d209e09dd3d648463d2d66f98e6d6b69ab2379aba9a9199e3490f184441bc3d6ccaa315abd1faf7ea7860954f215ce5094b1e0411a0fcd42208e8b07c1e4b2cbbc5cfe7b18c1a540bce2213fb1c1bbc5c8dd25961cc1bd8da6f50f40c01ab2c88adc0aa148cac1e7b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156f1195c13eeae6f015e52bb078244a27236790212238c61ee939491df14c4f49397572ad353d9e2f9eba588ac3b6ce74f8ae7366f2fc8ec1b8e0b7564dde305a2abb5efb07d6d5556419dcca9b8ccfbb5da92e3ee8c2a55e02a7fc41b14f5098616230f28ee4ccd0e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha18124c22c2f46f7a985170529f37342cd7b2cb3403d9cd029aa1a2119907fcc538a101cad0473813c1f0f0d148151292b1ec75f644ee6041577287bbc4b9b2ff7f4add8a765f4d9789fbca85a2681b2baf021c17982cbbaa5ea8db3c2a2cf2b6cc8dc42610ec518fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134068079cc83ea40a3f6d4ebc852f71cc6ee46287d3ab950d51ea427c4781d095f482e650c9d59eafca482f7a68a9152b8765047d2b0b3e52e16a55e1c6a562d6a1945b497b1f7da6065c9c96d64391938b89e1175552589c79ef857b832e3dab855266a3bbe4a208f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha45434656f8d024047e2a2b221a068b5a7faaa21a222a2fcbbf621a37631e27a5615e200081f6beace7caf8be84d65487a3a9d71db8991e394b5532e8b7f9b50c7a57cc01aab8f850055351dc72a036371965423f3ce998993aa9463af9527a85069b5cd0425953ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he619c2ff1e511aa8fd08f9ac5c2c186091dbf773df938c0c7594f6692f7750320bcb4c486364452fac19a30e3b12d98838b7510257f06b536493149d4da61b19aa4bde8e98283ee0008c2615774dafc7405c7f1ea784faf9ca20616c933720af00444077b8037d52d5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5479e666d9ace10ed2d8ac34a3392fae751fc33037a3b1f64f98be0dea5a6af051dcede73f241d17ebe8d604bcaec0bf5744ab78595429735698b9aa3547fdacc3963234fa76835b88ee3f425cd43bb67e7ec107773122f5a6f08ebf5cfd77f6d9f6dc127be5a312a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b634ffe29f55a69ddcee304a602fd860319c57f7fcc397c6b040801bbfe843164cf867108ef8bc8580f7136421280d19d52b819b2a24a12c908489a19fd4d3080816e6ea2fc00bfacb3488ce9a345893c4bc9eb07af3c9083c553f0c5ee24436c87b72f205359c8d59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa6f15bd6fdda35138024d60edf1aa5d4d2a9b6a1f61ae233b0699cb61acf160325711597133a860ad73effbda0036c5ea84f59c4bba5f7eabbb0d55c136a3c0b32e8544f600283f905292fcc88c4b6bb2db2fb6ce45edfa57e43df0cf98246c07acbb0b29be1a0f9f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4662248c43582e41ad4083410e7b8e97c874e01d85ef69f70968433cf060f44fb672ba039b326e3c77a4fa38bdf5646d392985a820a8630f52492a0cb428036dca20ec24d78997f6d904109bab0509cdc46587c5bd46082c63e8a0f1bba49bfff8432c852c6220d4b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d5b13f975d055f4e7412f10fba29efc6d5f5322350d4c77607c57bdf683d5ed3561ce3a0224d0ba8bb52ce298987062559571fe0550fd83788fb4c26708edae52e2f07a00c2f1ea9272a1bd589eff4b74f900e90866d568ebe2ebe93bceebb1b0316e5ce1bc88f6c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd0efdce4dc3c5f80391239ae0b91aee730c51766c5a0f74b7ca8cdc79323ac5b591bbe148e500bc625b8159d5ef7c84c2852ca40f921107aac471fa8319f691d7abfdd75292e303d8f915992b91776a50617f885462bb29900635b7453db6c8ec8642b5ee3d0c646f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde5b13fa8c1c260428bfa72f5d2d71f9aad06a25f1f16b281d49b13884c00d1dedd9f1691e3eeb15f23af554604cd07c5416a7e861397d7a68868c7f7f0509da36e22c52596adbed58d1881a60a0edc15ed0b6f402a6fc0f0f2aad141e0fa6071efe318e894bf30677;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2afbaff2ea64501e6f6318b5e001decc2cce8448c77009ed0e27a5b562af8208b687e58bd60c7fac4cca948eeb367e27629bbb296960885181f836afa04eafbf928e4752785991bcb5661b3fd2c331892a4e7d95253052f512ab12951db604421996468a2a2ab6a75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1841c72c863dbd1a3ace8b66e2652961e4153902dcba9748dc7cbe3df821ca7bb80b30005e9bf60d4a6f101f434a1299b1d2322a479bf3d85bd16489afb364a87a322b3c3c21975f4c31dce4122386786afa75639ba921a46cba3be35548f95a42b9e92546aa602e652;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f5e3bfeed0f16eb35098351b8c163683aea22511d39ff2c7eb1aa8400f964c22b44fd11f13922234d16c8082f5109d3c2ee44c9c36f1b1ccef2f7bf72cb0d918aae9a09d860045568c139ae9edf570cd8e2e9e191681a507c9a85323216f87ff92787e09e4dfc3dfb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15652ea9cc75afd3c13b3367a02cb96da9085ce6c79cbfeca55b23427c1d9f54357c62e3c01a939bc38ece06afa432b66f93611b42dd204a034e355e014d9f90b09dbfc73495a651bad285fda45fbb1a8819023d138c285b1f44e89db0af452397281896d1f4ccc666e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he32ad1fadd7a285ff3b3aae0000993eb3d9d445905b4f308670aa437231c73b1cff4cef725abc8ff47c50673f4ac7316a9a9c3ba63833ea0d296384cea3c6253689fc5cd06968e311eccb10e0d8c1c55c2e3bd4ec8c17c9035b4b91c92bf747effe7dbb88d04042403;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h908fc9bdbddb531cfd95bf1b43e576f57a9f5e8cd62609ab7b37f164fbb794023bda162de581d8efaff05fb175a4d5b4806d20ea14d76c9d070d80adbb9519c9b866a86c10fdd638cdea9f20798b32c6b55a60c0f453c4fc33445317592d5e34a4f7d5f44fe110a1e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bae8e5854f14cf7b7b71e2a76cde3928a0798d9cc01cb9c15774242e334ba68bda0b08a21f092be0521807cf40bda84bae0db351638a3849bce0f9c4d1df5be174191f7147b6c1e1f1fc0f5f039d5b91244f84be2eceaa65fe69f0938cb0a97186df8388a7ebdc3c71;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha87ac37e9a97d049c13d3101174a14b20336f68de5dcb4e495d1770f3e9485f2c237fe85b50f65ce099d58705184e228d80e3746193dd28399a31cf87bef685927d09b09fcc5c554ff3a2840bec46a0c32ab284be564e2fdd79571042d0520ad548236d1d021b9e7be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a85d68b1c498265aaebd2610a2f7cb612153f1b04e8d92b0ae615092812f8e8694480802cb9fd876ac1c483abf9df22052fab0e45d9738fe36704f8ce5b700fab07a4c8ccea5c0052add6e186bf9c7ec9fb9c3bc5d0bf90e601d4da4f76d05a55b2f1fd298d224c6f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h899ee24b7481ab4c5da668116081bbc98f9319006f3378ecc42b271f6954f36d48f12954b2ae4189b70225fe3f066f6deabaa67436a3bf1931bae93f300511a34cfc12d8fa47d69d79160700090cdef7762424dfc1ac0b9d37bba2433206933b09e1b0ba7549948feb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1370b62fdb421660ae430eb1b62b1fb12be713e91169251b614b5d51e9a3b055ca8beeb14232effaa1f9bfe67270d2fd07e6ba0d94b22429231686a0a6cfae4047859b1a3af644407ea0f18f330917b86caca25bc7ea4a54140a33474bf4bf41cd47fc7aa767a91779b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c8d513f83cd46a5a5b772c392409d572bedb940b8486a8a6d336337a8fbf8c3da99162819cafef0c0607bc8ae7803002b3cc048f2dea7ed1d5aa411c68aeeedca4de2dab6aa4f92414f20bbddc21e025ba54b91963aa94a2f39827d22766805f24bff5afdd9ce2916;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h766260f43658592b7dbda5540ab376c971083d71eaa06628cc6f45e5fb555eecb485e6996fc009692e0c68ce30cd0faf5f78df71646d76267dade0465b87843759bf190b725950c8a317b6a1a446c22944df12eb6b52df1165e0b2b61a6839125038b772220e87d2d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf045e6dd811cb812b5d94944d6a273c192f4368449a5c48a0de38faa9932c1a327a2ab50d3e3074cdafc992d90fb6cccccf36d898dcc8e118f4a491c105a7c24f5ebd74624d45377620fa4109639a6293da8fc964035ce508928786e21d25e506295ebfdfe70c9301;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fa933da5b7d9d28549c40f9763fce76568fc4b096e991f8e81227aaa8101330b9eb389b8f81c3edae5f6004f64e80e26df7e9ebd09a13bfdca67839ba202f7d8caf764560afc8175f5ebb75a170be6b3aea9f1c6a1c247a4e66e4599eb99ebb105aad7a4772f6e3d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19975d272c20ff26c0ba359e374f83d92abb345d1bbcd4cfdb979e42b76d08841f4ef3fe00e5c59e90a55493e49a81670496b770e45fcac1ddee5960e371d55bc880add960bb164351fca27a930508995d26718a0d648907162dc8120204f8207e44bf95d8a95b1ad79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd31818c4ef8ab0cd1327c31efac04dbb5d0231b9380b733c8827c8b78e08d054ae65fc0d912684069496cacca99f0f19f2eca18b8d69105473153a3c8010f176fa021bea818a719e4aa37a810aced4e945f04767500c172e2a7f7a98d314baaa0b22f32f0bc7a35fa0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae4b00238a209affa46b714a672853c55f3dcbc0cdf4c22f9544b0f6b6912a4f69d73745e6e3a23b914ee29deb30e9e5aad68b5076a67cf72fb90c9b1abb4c235dc8387242a8dd632cceaf14219be85d82e6d24837d586bc1cb67c16f2d8dfa85b007940f914419c48;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a8685e9c3711c23fcd60d55a3421b425004d7a995a2a6d64b682dfbfaa08841ed222e23b4fac86783ca753aa6685678740ad8a6dc5488959b6c54db001f07953ae5921790891aa266f81b20bd661207318c5677426b398d1e35de4e2be40f2eb5ab7bff6bbf4b375;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9832fcb649a944c3e282a5340e3a6f94ffba85b0e679766b7d14ca596e46ebb9c7cd3db672433291fa1607ee67f64c93d61a1011bdb02bf05ab3f95e2e7c5aae54c78f8f5563988de1bc89e081be6351b8cf9c423218915f4a44198ac54eb6621992f6f90d891576f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1268a070da81dd6a9479e9feb3e4d84de5a6211ea32387b8c1c1639eb753cf7dec082ff1b1222978b691ab3b0daf0b4855d3589b1f103a7f8e6ff9a4ec85feaae5934dad11965daa16b54350ca2b4a24d6ca73625f61b1e73b9a7fe4464151a92b7e9eed632fc2b654f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50a677ee46887e4d8d2d4af5abae24b1e319f7510ece72ee296daa432b35767b12bf315ee10f6b2a33a663075b2bb2c736dc659f7ef0a680ccb96ee573f9fe4257a73af4d5e7db8f2ea27a4a46a61d87452d2af77e21bb7f03b5111843ab3c10584051091aeea25941;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11bb36bc080a0be08c0a0ec6ee9b143a07dfa5f17929361154c35b5bd4b71a61ce6b66e6fe65b62e8c32e623e9404c7ccf88bb20a6c7b0b80219ce7c6dfab05abc75b397c1c40b8375b6629a9671747bc1c9a7c51f2f1b1200da8d854c3d083cf36740f1a65de0d2804;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1914a72f77f1aef11b1e27d5779d7e0ea37ba9ef045830a9f489e50bf726fb44485ae4c62161316e8bf9c3dbb73ea5e6fff40a8aec89ec4a48f03ca77c44016d48e52babb49b32047e1259a1fda8399e33e12288f813cda0b0d064f77e5a7599bcfd2076bfc2845e94d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8b0f3cae8e7e8ca47134bb957b3007ad6c7552ab98efa7923b4fe7cb16bc8c1626991cc9b19341ed6f5fb50124809029a9be5c080716b30101c0209840402f009d2f91a20667fddfd11ab483b01b9d9132e4ef229831d974bc709187825448e0357c562531b49c065;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fa202f481c27953c48e2398a120075e6ca7d1af9e7765b20f23e24c24252729636ebd7ca10554b7dbb2091805b0e2d894828c934a26774d664209fbe8401e699ffdeffacc79224d21c93108e867e1c9af959941df04b099a6c96df27fcd5c3a28255ade710f543311;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he99a2c5a8a56b3b2e9a080309d5a9ba7eb213a4678a8afd2353bceef6578bd375f52ec5aeafc812d5cbd204c16adcf1078163f196606871ffd87051197946e280d479b21b74958be7cfead85ce416d8987f619c9de2089fb393815915414b1d97579e094286692fe04;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h715ab6837cabb7fd3f47d32922dd9c5c3dadaed12aeb8fca13a12267d4423a5a6dbf22b2012f7b95dc44bea30205ab73a5c38484de9baaa9225b7eee06b2ec60834e7d809160b91e0d4f7720e57e3de5c695b7b99eef3aed79a7418b2bfc99a8235c491fc8fd881e09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb6f7a02ee520ce3700b8aa4e48ef78efa6b09bcf9a490f05fc5924f8f586d4a190155345d367b8f77f7eae1f1e996bc3911e15592770758df8e3cba25bc8a07c384b1ddcdbf36db66841edbe8a35d994ef8f0e81e0835e2d84411920f1492b2ef7ded41ec06abeba5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb7e76c1b7e2b563b71a6cac1a2b5016540b4ebb4b88d19828bce5d70ca52c6a363d9cd29713b22c1bbc069defe250f61d5034b906d8f1c5652d80428814da8dbedcefbfe813515e9bbc8ae4cae69512a575436ef87203d61ee7f700f641bd96adb225fc8d0d75e6ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha680892ed35e2b124b76511a778685639811164962b5b39a61a0b971ad772c467f3485681c0282f149dff0cd727314fcbb608ceae61d2261c2b4e3942f768113b9be97194973f1c106eb17c69321420ea4ace769d230a06d9f062ca056ed91a1b5c760cdbf652ed71a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc44053d3b04bcfa679038eb2db5fc0df518256ffa2b95b9813fde633b0a8fe65175ca5f58b41266848b4e8f529cc6855ec3b6c71d1f208e92da7b9b9bd7d9b85617535bcb4d3433d590da9a5a0712c17c4180bc59c687460f3d8b0d697a8d2e68eca9e9a242c58a814;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a67b84b842e353dcceac8860278534267c825e91c131b5b1d59572fbbac3171165f93685efa7763c04655b95bb6bf7a8fcda5630fbb645bc0ed5987c5e9a420d872a6cd775b88f64969b1a1d3af8bf3242174c2cf07cf5bc2c038435dd5adb62bdb4a65c4398ea5b07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc919a0574f9e1f13dc6c9b96598d03dda1eb28b82656e49b1235fcab130917565cb3c3ddd489fffc319b510ff0b5b1dc1b7b6b1a557981f655ce6763c5ec974d6f3e81cd1cc2e5c2409350b988ef88e7ddde3565a27f9fba0e3b46a373911f7cf24ac0677606839bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112ac46d265f6b16c2da8a92b33767ba5c3530dc7830d407e28ecd6c403aec250beef4adfeb95a49ff265a2acfaf2cf5aad7760f72089a8476433ccc8776dc7146c91dab8efe2d0ac8be22ffa7cc1851dd7c8e48743a6ea5cd7f23bb65c524a74f471fa7ebd2ff4056c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h440d0c36fb25347ecc855680568f8495c4e7c1e4d99a8ef2c9c56ba3ac1580539366f43c584082f9a818d16dae1747ca3259ec4981f5725743746829d97444828f23c45fd33fcadfd96fea274cc6c90adfa7ffda97345e761685ff21f0552f64f825e6e104f3d1feb9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3a3ae6fbadd088c9704b31d4b2f5b7e9ddc396844c836dafb7ebb88fbb59666314be48eeb05b71a62087423a314d90335d49d5907ca59b873b16890ef25b574fa363a2c4917d507d4284b8535af90569136c99968818c0f02bf9288269192e019606105a3b24ab1cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b702d69d471eba6654ee71ec8fdae1889b225b860e88444ceb6f66988690cda0e426d7c42f8057209cf4c61068e2915a286e3376c2fd174cad75557aefde58c44d59f7e3ae60fdd23f3b70a202325931d9d7a1a80c9c153eacc7159eadf3b10e05a0d4cc4a02e5595;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42186b9b7a94f308ec311d4ccc5c4e33ade8e85758cba8cb495ff7889b87c0113bc34990331d99a22041cebb0788a1c5a8e16b6dbc509e25238e0cd2b751461fd54f716bf4111a3feeeba5f493bfa7d1ccd3c46d7b14308a9944fa7a2a13a63e56d1b31f91cded4eb1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aaa1cca51e83b6ba01a4971e36616d06819520f09f97f844bfef146c2b6f540e903b823641e8060dd20231c7e497eaf886e9a66bd129b171a5391f2592457d1b8154edfd0914d59c47660bd303afcd15c8dcf46b49861841df4fdad7b566ec074a170fdd8206b1a8bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1c5a526e11ca1603b8c15fee4086c7dd7b18dbbbc2cdd848987f223c5daac194f6841bceca0d8552996029ed5c1746ad472173fd2f9d7e54f3a976a115f262bcf499b71093d4cb5de89c116320ebc0ceaa709d24f6002f8ae98624684b9d313fa3ce136e97e39d34;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a47e2753e04be4af864a08666700fa6bc242e3fd1fd7ad8d655a508995d4c0c001914eaaa14f3c2d06a61162ad16f8ec536d2da4a4ed05129526f7d39bf593fc1765c176a4811b58259a04bea746b801e39d77d4adc46c31f6d14e342d81c1751b63d0984f202dee2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b72ad8515f0bfd70661ecbbd09ad3bfbd28988342f449f8b9d09c9804278b488651e3f575b2b789990f6dac7cce22af8d84a1820c1b6e7b9812536fbaf4e40cc9a551d4ca21379aeb7c7ef68c1908973447272b352f0d68a5b574d20e99ad9037b4622ab02a499318;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192db6466a3c739ce18104b657434778933b5d05a1d146f0e74745c2c3e8b156e0daa15207af291ee5aeb47302c4d7834bd7cadfcc3217292ed5a836f38ae30e3ef3b773aea754a574cf092bec74793ba054fa03556e162513bc26ea88653323e40ccf16194cce1d651;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c9a35d824a991a24b4dd074ca744528b5f9777c3c310701bb546b61dd7ee7de1c84076ef472105c95232fe39cc0245593ada2e736376d2f7c2e2914f83fd49b3401c4f4b1a5f9e6105c9001e68e6bb3568ecf96853ae0935f9b9fdab9594ebac89a9090be19e6d3be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193e34c593a7745d8ff82c0069e601e20f97b928ddf3425b086b9105f17645f2697a87ae6ee5f011f49dd0fa37d236fd3540f56ffe5462cd5105dc619e581402a2cc5d91eab38728dbc717ba19c6f2627b4960f66bbe03467900bf011cfb1ef78df134ccb7c60ad5f56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4734cd3807fdcea22f70e998ebd1289b3802e12817b3a174f6041f6206ff570a557ed6600c435df7ffac10894ed9906c4df9efe827048eab9d51230e6812d79baec3169ad6e99875a519af9cfe3f77d63e437b7e75ce120612df0e557d8e3d1c59758b8e5d8a2836ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c1c79b917919415a6bf21b13e38428312c2e30db4b75182944df94e975cb9ab4cd045c53188051491fcba45df935eb3931761a0895d255c4a87addd81711831a0b18f62f41381617dd39c0c2ba68d16e0098ad44dc1d9ee334ed2bddf2da52e47b8d85028412a4fbc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he497873fe41341d8adea99cc6f817e935243893bc8babdd0057f4423bb45a0d7e2547846e1d0e7219c3117a8777c8dd6bd98c38432a66ea23e295c2440183be77ebbe7b271fb911cc851cfcbb5defb604c42e6c226196a2401fa0b8a7e79cf0771c61bfb34e298b95f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51d1708d8ffc63831f642c0e2edc7958188fb22bd2f03902871bb4d27e34fc802fa39f82418b7a1e192702b55b4a0851ccdf94c4b01ee756379746c39d2e2d8e473e468b7289a7363daa3f1aab5eebe1f4af1d6835e78314eb2473c523a0f6b01f7f0cfbe46c73b422;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1397991656eeb84f90ed30a9e686dd7f4b9d650a9dbffcecdc26349860b19d638943d663b9ec4c034812a6886740a36483c8bd443cbe5cb4756cf07c0a8282605515cfae942fbbd69cb59e6524c6e0478d64b290df1fa4fc75c348cb9f916b12eaf624b544e7eb762c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd11898760fbcb897d622439d05f8d764f577ab05cf4fadc21a536c9a411848d3ae415f720020315519e2f29cbf177b5f8d18822c1524ddffaeae20c75550c6f03d69444bf1c36a9360e6a52cbd0881ebfb9297e57f4b75bc6aaa3587be76b667ec195eb17f689e841e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a16893760004a748a4dac6d250d52b344b2a3fd784cbf5868a2cc74c5cbe8e3d3a87e9974ffb65c36ed0038d8f699a84395cf840320a5713a5ffc94782fbde1257934caeb9b0c2109372df047177800ed1294541dbe6ee6ec707cb05d865d74e7c75b42ae00c71e2c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6a99ead79eeaca8fe6b76bb2b69057ee3acbbee4e37c6700556cb20fd416bb4d8150cdb70b3f085027765033040cbe10cde8da6a650f35125ecec8067e4df4f2f5ef9ced935ac8530af9493d953c75869466dde81c55eead498499bd96294eaafef00a94a7417017c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cb15aba59d9ce65cb672d27a9dbcba573f0faa6e386108996823212f09253ae1aa7745e15b23d8217a70c1fe6f9df086cd54cb3050018d3d6b8e6fe06b58abb67fb7875dd0f6dd50f232e021f4b00153fd21376ebf13500521ec8f2bf163f4262aee4c309b7d82ba4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9d5653866093c1aa5f4e621941ff00e0cd6605e40e3ed27535473254e15b51e7d995bbff0c574abe9c92f16cc5f5401d1e40cd84783580170c2e1f0906cefae7db4084671ee9617c4499687bd24be2007fabc5378b9955164d59ce8454eb84873b2702153c28a1079;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3028aa6094fc528f74f2cad4a421744dc0c411d97706e21e202abf509202c0b1f30b3c27785c29a102fbf9c81b43784bd8635adb30979847470e29fddd59bb7e07909a1aa53fc6708a9de6174ba0f82e25309d70a69a527f69a109f90896e548953dac20d3237d2d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173a77fb656690359ca1f77faeb409d5a0a596bc096d8eea2a185bf772496e8459b3a50e7fb217345df78c0fb108f3517d2e21a12bab5ce652d3421072d32697124e6eefaddaa8868152ed58d182b7fbc85b1fb6feb890d082aa3e31d7f5a7925c502b567f039c615d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6eb0a16ad4c89ece4c60a964aafdae26fdf5b45102cad13fe6b3286cd3e10395e7d154b4381f91574d31a75cace9fdf1bf4881a6d8052476197929f0b1d25a1f1d07c29292ccacb7f8db961249841585f6283fec8496a0c8962f84911d7528b9e4c99499eba420c29a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1735dc27a679c1c4cb6f4e80600351a663f6130fd84c859f81215f835cc02817ccb3c5bd6c7dd489e910978034caa84a76ef6f0a17803b09a662edfa90b12c2f5c1dcf609c57df46228ff6300ca736fbd48b934d94fa307891d897bcab1b6e8480974e81d7c0b2232a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14794130570ef4d169ece1abdef11f545184581ad1916599b42d5e1a79854fa3127625e47207a218768fb058e293e4d76cfb888fdff8e1d06f39cf464e559ef6093a248b9ea248dce2b81e917fb24b19c0f7a7063251ed2b2d79f996907860e6796d76709273af30133;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d1a24fcba272426e93b1cd992a91ae690c34ec1df7f29fe1d0ec91354c096ad12409770ed2b483c61cb7dd910f67261cc67fbd095eb2c9d1769d8c43df04f13dd603d256760d95980417c94c695da71b40bedd92246909f803f7e95a8b364a0c3b1c8754482c24fd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd35fa709c2c3524ae930f856c22e43c238dd1ddb48d35189b49ee8a89ead886fc2cfd710504d5ca0b8cdddd74b278279b378ebdf870442b1441c4356bc33ed0659945c342909b5ed963ae724bfda995ed9762bce214819b43af28cd5cfce48c729f68fd02dccf5511a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef62c689b250dfe8e6f962ec5ab3eb76b940258d067ee38b04a9c62a49ba89c1c42d94dd57d2db9e9d9376f1b91961b6e11eb01565d3d13935a1aa83284fac34f0a820107abe1976da38e718ce5dfc3546dcf218090057fc3cd0c303897897eb7bc4dc52e70e1a3312;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f37bc518eb07a6296d383f4f9d0f7903990d5f4afc3afe1c81f0a02693bef88dcfd0d4852c4e0bd4438d92e2243107c3a45b61fe3ad8fe774270fdfa44dfb1ffe570c7d5b854692b299429496703b843f002da3b69239c730c5068a7e3c77c8a3a32de3f8db64ab826;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1327a46d66e1b6a9a33bf1eb01452034b6b18cbfbd00f73b86108159fa917b9c93ff3b814c13ab3bd7ff95f14a3b815febfe90137ffbad6549b46c3b386d59e8175ef5fc906a5fc2c97c119da697e55b8decb6491b01cfceecaa9562a1269ea1916fabbcc65a17480c5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d584712d762fec23afbaf2938f7b29aaa5232935bd1599bae0a8b537a54a17890f0c1e2430008473ae0cec92c09f0bc7a5f320301746a67b2c43d4ec80c98baad7a62f75c8639d9b845d6e2e68e8d37cb5442c4af42b621298056b6cf19fc8daab730b605269eb8c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13cd22ad6cba94a6452a5237ca7d3531a568d300069df4d3c2fdf8b255a7ceffa807bfcdbddbec9bf4a890b5d89445cee0f2201b801e03fe4d46a7bba0230acd824b48c33ddcb3b95fde8c711a490ccee064ac17181258908d2cc8ed0f3930931998d447205e9a9732d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3cc5cf9f4908c899c009f7d4e6a2d7f21dc8a9a26aa959e805396a39a463c547305feef196f9665f8fc75e3dce5eb3ccc6cd1ae5f8039fc37515642cbc33155c3928f52f3a3c3d431b0087541e3678116c38b425a97d6462af65ef5bf9875cab4aac931daabca0226;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58f8402c0bfa70a1960a42e64d568a481f0917c42976e8766fa98851561899ba87737dc5f8e4c977596f98cdfddc11d3ca3edcd83ebb2de1f2871e8b9cfd4d5139dc86147b5e2002bcdca81e9bb4c3ad1b7ae01002fc8f2979b94ee4d82710c1b8f20573e5fea1b186;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3ab4586d54ad26656186fb2ec8bd9dfda928cfa9f94e558c4a6897c1ab8dcf59540636ec757542e8857acc14e4772e981709d050e75eeb01796f0630852b3543e411bdcb35cdaf6fb4eb99029a1e616eee255f5b28b7789595e41a1bd7f50a5af40b5adb2c78bcee6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1949a60b2fe0a7cc283ca005b9ef8cd9c59d89bfb56f1a24b647a018734456b5aa576070440beb327f33073354047ebe022baad9fafac6fb5ff495ed0a8a2f8be3dbf2d99c03af25940a9fb67a6b4457c9501bea1116e0ab44f60ea9acbd21a89ed455041e82f3cfdb1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b3b6be31c2cdc35be7a0e796365b76744a8a94b007e8376ec2040cef62e83d3bf06e9f128eb352a24dc0443447eed7bd4d0914d69da6bdc0bfd72a79ba0513a7095a2cfb1f1b02850a160cc0efa0277905eefe01208030366971a40596dff678e2a644849ebbffb2b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e066eaf9ece02cafd8b3029bac96c76c5762cfd5de58ea1682e80143ba12107fc5eab4cdf1857a74a6b75b1465f0499d40ef3eab9e2896d0e3af3b1ce38a09946f7eb7cb01c77c4c3cfbf0fe7f58cf26ebb782044b425854091b2d501f5e3a044b2a364c8622f4458;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197b2c14443ba3a6bf2e7385caefc3d8a0e661bcf93c818364595499ffb48e7aa47c5a6d5172365873664d8bc3d716c025390a9d564c4a37d5d98ea4322dadeec2340fedb801fddad22cf404e4fce00108960cd76e645513edb0e6c1e06780a9da6bbd9ba02c17826a4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdcc80d9507c15ba1c65b1d9e52347542af19af93cbd7dba8ea1b86b26d07e2f70666eb8a8f3820024f4a694466454508ea6f2cd39f6405687b466d81973d6820a2af5323a71d1e16904aa14c8e4f01a0e246e2fd85402cb29f605ff7e15e74608f5694d9868e0813d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190e1d3516a28678c14458eecc89886b98d22b3113df9005cdaf73894c655087416d32aa75a70b8d096e275bb2bddc569ee1a0c2138d6dd0176033ef56e899636d9826aa030df90fecafff10f4541fe12e27bf2c3677e9edb8ec7b462640c22572ef3bcfc1c8391d6b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55e267ae2bfdc2d9d6e19445598443aaa5a7a8beb0ac8bc9793840f5bdf3ba4690be7a11e37bfd66bf6432dc03ac0d29e1a915525e35f8b4f05ec55c1f49103e835a2d8f6cb992665f943e9ef412c19ac1b2ccd5825e0ff6bcb75f6fb84de267710ace003565236b5b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ba83dc291b15587a81346c01b7fe4cd3a027624232f8b6f4425d26e266465b5b644be5af3a74ab2979c3ce8e1e58deab1713af98f7596cfb1a211af3bb1a2b285b6f0ddeb35c3c912b102b94525c340c6e0e51174635483b38483a3ad37b1cd19698a849c66ee7b6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcaad11c4badaf0b3d6e18330d67d3817ce18c35ce88925da2c435c247c76fe2573d525a64def5605bbd57582dc863f15edb854aa6b6f34b4c713bd585c72666c607926dd3d8166f598832ad9660a5fdd55d69c1a09ad8bf944a34f02756cef60b081c33e65976413b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4f6b8a3bf483105fbb665fc6d7a2af60441cb971822854509e878e421f0fdd6c21498c4bfd69a3bfccc1e6a9a6b0fd13c6a85e054ff433ee0c657bc85c372a50ff4ced42ef07ba0986858bda7cf39cde9d4a2deefae41fdbe50baf360f1e136e72ea031535dccf606;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e3e5d715daa377bf07ef7b4226c5a7f397868ee94271f1cd3d7dad82f177f177e0cbe00069a99a5eea2e4d2003be4de1ddd684fa526dddd93a272d74a8c70b4fc841d187e25b96554f382f84a0b36a8eabb18084b5790a633132f65f0b684e7b75f7d008085da7391;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58fe6dc2cec08f17f784794f254cf890c752f997e0d2f849b9e21eee8320c2bbf51582063502bfd790e7a8cb257911ee267bf4a4db82e4e5aeadb14330853c07604de51c59bdc9d0ea3d4aa83b4aa8a9c9aee3a000c66b83c1f8020fefe001c5d6d3f5494ec481d7e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h462b51db0ba98dba4f90a23d3ed053b0c94a19ea35fe65b41208f967cd51f68fc360ec64b48bcd645a2ec46ad00dbdac39a44f95703f451c84b406f7986a03e1ddf2bbbfd915633eaef126725d0ac6f66bf98f61279aded0e03512d990643beb86478d4171bb6d65e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abdd213de079e3d5ee2229037513c53fa27921aca9bdd8888ad6d03caf4d0f4edc197cc878d541e15ad56fa7348be70956795eb2519944c2d6fb864e9188c4ac9031fb9d95ac9ce2bbfb6b4637d7614021bb1958f5175848f05e25c8428997c572920b10f9b884155e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1963808ce7addb784898d26ef798c7a9318ad89d2c2119a12cbdd58edfa4bf91ca4ed8540b7fffe4bfb16cbda0c64acb702df136170e6721102ce447c2ee13cd86886067e4c7436a890b1b027b8cf21ebc177b579fd1edf166f7fd3a7df9bc2af7029e5816723aea2bf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ae7ba6c533b281a0e8c3ff1a1db070400e1aeb7db5a6416a7c920e03911a69e24604010140504600504a5ab0e4a2fdc97175e23f44cf14e626fb140c51d904f6ae842c22786467a9e6786fa3be3aac7e034e62f4453a406923567da3d1e07e39b37c5e25d21bc5e12;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b84f3182101921eb8a2ecaeeb7446ca240a363ce6cf4439a9ffb170edbf6c128e5ad76b15004f551ae42ce320bcbba550d3380080ef2611c50f00c7de39a195ad667c7cb23f6efef7500a6dc0f8846978c43c687f2f44812beb06c4e8bc9222bbc98bc3c6e2fc0157;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f82256e9a0e6451d0027810f21ff751a0776cc82f671fd5184da77bf9a4c9820e7dee66afc37d27b2c8363a908e949d756fbf1187e79ede970febbcc94587d9af24d4fa28b5f9010e2c87eca7f75310115b7cab736b4d9f97bcfd2917876a07442a52c570d0748864;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5a588c3ead28a9f20505527908f75d120247866e2ab9386e8ace23aa5821affb42a1da549c85f40deaee1ed7e7cb15846ce3fd48b97ca217d5a007140be56129628155c18d6ef3ccd0702ffee91ff7b7aee76d5bc3e08176b5314edcf69948c51980c44b9ccce6595;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166f80017816a00aa077a56674ee1a17331200f03ae3d531b8740fb70ef4627bb30f7acb58a3b8438476b46502e8baf0dfe354583fa8e1a4551799b237e9876a1a0b04b82e38c962652504c3d0498faa63341e1627fefcae953466333a2bb4f21f92a42361836a02a52;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf23505dccfd1e306b9ea3038819ec8ed42d659da9b323c6ee2d98ac546c6999954b77cf0c34bc09650f4d33e872ea731bec6b8bc9bc03dcc36582f567aa43429aed31ee1699ecdde7f1f1bb5a1cc4e6386ca4aa2a8da1fdd2fb6b188031453283a31b62c9062afbd60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d48c818355a5ace5681e41b07eb4944f781d45aeb5105883e45961ccc36affb0d832d8e52738e293517040cc415e0fbdd8dc5157635efbd026bd7109c7e4f5a6868df32a47f911f30caeb5cc8d3187ef49c21ec98ffc78be223c3fc638cbfa3e966a443cca7c2d214a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda022c3ded2b7dd023a5ae6dd57c7464c2572e5c255d90313a6aa81dbc9de02f509c543bce4c441e5e7882fd129124fdc653b419fc32ca3e20fade590bb8cc331c4f05f9cde033dd3747829b2ef13fadbfa06fd2d1b526f2ab94e96ba3edec89f2d8439ddeb0809b49;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f95f1ba8dccaa9a7d62f6f34cb4d99e1f4070da4d202c3fa1894c69cdbb22894391696f4b4051a22335109e75c6cab0f4b652ec943806a2f6251b0d36a074bd250e1164d5159eac12b92f8053dd4f0cbeaedb45d8558390fc03d01e0b2649923eef36b8682240ac013;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172709a494cca2320dc980382943c318847a0b9a428cbb90fd400e73684c863aa2cc32cb6cb3d24ac958d7951495c0665124e807ff0276ffa2089feff7b13ad45821830217f3eda69730f272309d2c22b849bd7da20fca13d346cdaa56c798102815bd8cb398b574edf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a42fdef6cd44de84b7a20361908013ceb858f4d435de9092c025991daa3cc5ed33828479cbfefac56a8533def8fdc258ff26ed501404cb6ebc87f0ac362d8d5e65e18edfc57c5024167406748aa090d9f9fb189d62373e1da8a0623bc1e0fb8dbf9377a33207b0e13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145c7cb3ab16c6917ab98fd0411ec84d9125b383687f2669b8695de586c9de95a766fefdd68241552fd9386a1bcafca3f1a55007bd77e115568886938abd30b157c0cfbc02be1bf31955e35869e32f7fbb1e943f10e208f3510fccb8f68045e34e68bf1952062a5ec3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc03d118b5d6be0f5b88485a02c76d33c54680a1092092e469278930a0d07e7b5a5cb755015719cbfabcba6d048ce81f3d28afafa69a47b248bff4c6208b8d81ee354be072a81fa4c94d7c039fbbdfedca81f9c5168388a3374f00e5e80767a63f7bafe1e89463aa51a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167cbc28d4827de364cc7698d4d3a4ad2862fab7cf0927e85f9d656111c2e82ebc8312ff21eb4def5c549fc2b02b1c779a4e3a1ec393765aa511030d21d7d9f86fd1417a820dea293b3f9dd3d6b3e22aa82e4f31bfd33e73ccfd4e0880bb9c9bbb7b07a23d6a2ed4251;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h98de05925c56a6acacd49ece4f49e57163d55199176132fc8e370dcc0780c8b840875fe69e054b8884fa13f4f532d745ec55d0f9a8f33fc1c7d0cc415203c254f91041d11734b9a5abb932f08cc84c50807a1e047b02379b5f04329456f389adaf43083a834971fc54;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56b0a6190bcf71e8b0cd45a23f952229678165dc8305c90dff5472864dca8b4d2926b8631ff6b228da5781b5b9c1688a38a32af737d67a8d41732e8ef54a005cf8517b2bd78d9b75b262a770694555e86240f293f7f05166f95be5253df9eb2546e353d8142dedc675;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccc3616e1bc7f50f0042e0e23698f3b6e69bef60210caa9b07b9b61a5cbcffe66e20a5547d5a27496ecb9d1e4aed84a472289985fa0a1bcbc447c53fff5d07a2b2855518f644fb1e63ea38519201c6ee65a1f8eb2d383528012e85fcb6b996581f7ca58a812e5a4615;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102c2c8fd32a1fafd077089f24de08b4d08539f6b279ed1d408d8d4e4548a8f4729bdef5fd598ac8d0f627b6fcf903f79f0e9e8e6781ac4f3d1763bb275f23c0a5f61735cbe5c5e347bb70c4d71a086fa6866a608ae857e91b28a61a9676d532b6ee484b6da8e571d72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36f22fb50a1836691f0c1c733566f1b7b0ee4242ba560e719cd93b91ff5431233e2cbde1c0f66b3428b4fc953492894eaf64d97592da742d77e991bd021faac119d6410f60a27e88868d0441ebaa2d0bf8d06dc878b4002102fd4dd2f6cd21d3e8344515d7fcda448b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e1adc6ded18278cf91e97e86763c16ac5338b1bbc27df1dea560ffe06ab2a05ad00b5fe753346deadc8fe5e8c9dcec25d57c5ab3e0c4124ec5fa243d0714ba3cc9348c184bc71e0b386828f35d6a75204ab1d32eb3255dbe9eb3d9091e8a46d180a629bcfbb45b1dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbff9598bd8faa75ee0aedf5bab9624de6e2967dddfd396f31e26b6d410fd6a593edee5f0b26337d1a3dd657918626f261cfb95f251ea7c0cb1090d67c10053db909302701319ff28a275bcabaf4a236de0bd13d2f625a4b3109bcea019b475ce34761727ff8e682c7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108d325fe20cdb5b622a9bc637f6c37bb253177b1363c226bc35d323ab90319f457076d01e6b4e32bf56a55037f73e16a6d8b2b19fc1e87d8446883ae62fd8d207d29bccc2c9ab817c09de226be3d429456d6178b368dbc0f98d8e2275be8a2643da9b79b0aa79f2084;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62b24b68a0d05ac6d681ef4fd665cfa9393c1bfaab137716be426bb347849521a4470a9d7ba9278ce30d6ac679c3e8cb348eaf8e3cdbc681f794860eb9acdf3f14655c4337ea89da1508d40631b14c384330bfd5b89356156413c531e0c42398c1f317fe6486a12f63;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95d69ca40c7bd5f4862b839eaa8dd1c73d7b190333d2fba0f0e92272c9bc502806b6f4ff8652df38500d64099842192d49abb17e37805c869cadf798fb20a6ddc6e1c3396d499642b71e640456a1f25f088e7c7794a108e4cd5d1a8b0cd1f372b0b40d3c0c91008801;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162e18cbffa7a0fa600a623e68303c90d7f4acc24e92ea0976f5cb0384e4508aa29851093140de48b7f70e7d2b6036a59897f07aa45dbd866722c27d32619b19eabbb05b83af6d0dc04c9163f248b4f5b5eb6aa8c9f3a38327e47ab73a29159e1a1738ecd5e98c7660e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27c77cbf78ff2a9cb7f23a1f8f9b49285c18b9a4900da0ae33849370559514bc12b7941b9b15e705d768d4b6796c63f115eb6ff33aed0e8800af463d4d2eb0b79714136ea4ddb7c29c8a7fc70f63f4b27e5fcae0d17e7d53532e0026fa66fb98ac4dd5b7e50828d428;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7f6cdaecdb0f3c85ffee670d9acbb7d0605635a51c7e1b2708f710ae5308a33f9dbdb9a85a8dbe22c9d5cc0053d5b2b0a335c86d80a526141b8161692264ad1fde185510cc95ccb5b2bfe7f4b2e128c7c34b56a32ba95ebbf11545dd7108d59955061d2f3e7af35ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75d5ca38c862f2d43b048557008d996fc564ab13e35daffaad200920b021f017035609d8d77a414689c7bbe9338d5c2ec1fcb8e69e935728c905cb41dbc47a281f9cbcef1783b0fd5f4f62b49729c8152d0cad7b3034c87d8f5d98d73db09d3b7a61f817066562145a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6fab08bd93a805fe838ce8c4d118650c705670b7882b14204300e6acf107b59b4b2ea8697065e747ec5ea0887181572901b38b3eaa53c4100b7b4b49f7cf2417b5e5bf1a988a81b99310b00681f400cd77d9f92b98cacd34a9f3c8af605e6b31665dcc2fa50c98d006;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da50850c388d3dadf0f234d95b1c2db39d57a91910445d31e80bca01048f95658586c79b7c97cdce9d64b4e8999970f196ec12dbfcd41d4f806e68f94ca6e082ad51fd521033d35ae44ccb7e08b4a241e6d862177fb005a9cbeeb169439d59614a70f2b43cd4f1fca0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h524dd67b328dee52b6ad6140087754b9744bf22155be32a21e1cf975722a6332d8f37530f2ceaa0fb067b54f3ac3f9f8087af4a52b5df565c35321f4c1c798f552d8e6bc976f260d93cd4f16dea3879e877110c6a437cce7c3c32a4095fd9740edabe9e9401e2e343;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de5703ad97400311a440816f005a227484a5d3ae86932412f9961355692225e8a90b0f3ca013f717a522057d6ec0df9397823cfd73c6e62187144b8eb803d9a2bad0cdd62e9db1cf0cb1bc65df4695997f95c20e08263f804d04cc5c304f97d04f655ab3edb13563fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ddce95778d1613785e599288d187a903638c780f61595276b31354fb7447c30537b57d3a26d80a1a66181907632266a1ef5202a5479d03c4e076abab487ebfd636c41f8ea0f64f4ccb96dfcbf02d84ac8e880a5a9e449f71002e90cdca07ce47500632f404812465;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b011295c031256c4efb163d591451b7f8ebe823db2bbb5c95b59b9599d10f51b636909ffa46253e1caee3cf7c84746ad9c7262423ca5efb6deeab2d65dd606a0bfe73302695ceaf8e45ab75eb01fd2ba7e1f879a2ae616b91e3cf3767856d4b5ba5534844f57dfb80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd9eb3b2e7139c80f91fcdb06e3fb52c41ea6fda160d6ee1ec4177f50e807e1911c413ca77778eabc0b400256e4bef4fbe6fa0da85f1e3f199081f053c8da42a9c7ff2e1d361b95969ea39c3cfe04409d1f7f46c8055a4830a4cfc1713d43c3c75fd26e73f6a0da08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3624e1ba9bd5c7e78f07731b696aba1e4f2646b54f33752b27de6393b0ab60110fe1357f595c299ac9e876fb4727699b65cddd87fd45970e920b195c32913ca08ef6fe40a19f9da4031c1bf7f41646a98ab8f3f529fb56dc37d231439779f3a8e48918b395a2122ca4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd97c2e88839bc356007604641899875563771ada929387a157f66249ac6e8f3297fa13c8b209d7c4c54dd4d5d400160a1e22f5bca309bb1365a43907236b888cf7f9a93d26cc9d06a17e130f490edbf37526318fd996b522961c6549ae476317bcd0f4eb1553c96a0b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3aced16fcf519b15a0374a8fa9dd07de0e4680618aadbf5378c5c001cc046423259f0dbb5b3c6a2837c30c236b9b592642dfde3777c16607d1f37601557584157d7d030c5c0e6dc68fb55cd78294937194571228a2fad09c685ddfc30ba40c5ab0c996db319f25be08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e03560f591be43afc091c8f7e0c34fc8da23b9f487137b107ad4d91316c81a2a69b191496ca524f587ef75d93f13c1efc0fb76ccd65014840627bca5135aa9daad6808ca4e370f60827772893deb93372d45c53e482bee691d91ee8025f6d4175229873aa760ac671;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h71fca63826781c59b6a92425093ce5ad91fc381424f7ece7cdf2e740c1dafd84477e13b93c95498f41bded261caf3ea5f3a283424c60e04f6d4b88a22fe5b9b46df0798ad12deb5e302f5b6a86200583f6022053d0d0d3c0c85e6068dd3aa39b223e332142d41ed7ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd82620280bfb0b632092e021c0c1b9e36b7814d1b26b50f23b34f2afe89ec7f2869c8be15dc7b8f8ab89abd884e1b008185426ae368dc9a87e7b8666cdf50f6ad6a5ef8247adebd514900f91ccaacbddd71f8970d6816ced6aa3c3ed1b0b2e495c0e33dec8abeb5ab6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9163e27b62596768e112b6ce9824fe4ead77852b01f84ed59a3510ca84188fe29767136c12a110bcb565b7c536383bd2737a8c5c0cf577071aff55aa2b022fef4ec227cfc42c2c218c9c5a35fe3f45c1427d38fc74cc4de7312a086c5219c8a29d236068a0c203eff9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fe530d50fc7431205507681648ad80ede55b6150db8f8038a0e2300c3c5ce8090b296be06e880f9e9c1df75fd48953d26c428ba5000bb77dda985e7eff4441e4665de04df3c4873500c9907648fdbaace971108b1e937b925fc852b53d154f5b6feeba90a8bb8a7d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4dc2322e57328e24aca4fb94c0e85d86b0c6b395e73535db4a8a012918326c73e7f67e124e80772b4091691d4e2ff0403509af879ccd8b5b5b6df29fa2279064d67ee169e41243fb3d52a323392d230b6e30809825f06b171e88cc2bf8a73192e5ba3366047179cd8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6378c8c8005d1931bf3197ac66fc4b069c6475ff737fbde93b6765576b1ec17358261706862fa4580033f0917decd67e581ae087b3628546e0e1387ba23016b277e37b910849096567b2bdb25e897f2480f6930b4bce43937b28e02d2752bd8e50afc481a52aae238;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116a3e68c4367ff8279aff37231c7db03a7dd962edeb793fb9507c98f50774aa7fbb4ab3c5bdb71b76814acaca3e4c74c6176c4cbc03ec61b5828ff8b2ed76c0b2608bbfc70df68a8d56d5501899007e758aa67bbeec2aa9593b577d3e17dfca35680ac557664bb4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h347b19adf1a472cb4e19d8567dfd78a4fe7e5e8f84a709e601e53f524e687850c069778a3088b32aac5cb4f604e67c987c703777c3bc57a388d79e40c698adc69f7bc7d835c2707a1391b8a6719974c92b38955e7a5ac1571e050dba181041f91ebceeae00a575feed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175ec09b70b6696ae2adca67c86066f7ad13b7576463fc5ac1417183a6d8b520c4ca4aeefbafea509f574dc89d90e7fffb57538c15ee0bf2e887a598aabfcfd4df7e2ec4781aead156ed25c3e1fe8454cc3a72e1cf9a156634adb33386bf52ec37872a5770241cf1bf7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf862d72b2c8895c17b9349bb7979f806743be33a157765c47d0c7f58faac31f7eed9477a470b1dab2a7ac2161ee1f112af1b45405b1529feca79ab596c81357a07098ff6d6fba4365083fb50891899368a4b8557d35820dc3513b16dfdd9bfd5f1fd8558c256c6c9e4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1727926109d596f4889af339f2d38cb909e332257c0bb19f49e8220ccaa0c94a7e68087d2fe3c10519fbf07a8d2df5d724b4ac0c275746b034c994e3758981786d8f11191004fc28710889c7cb08847c7173de927a6dc7162eafd62495dff7bf8626b2035bcd7fae412;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8549242594f8a9647a45ad4d0c27c386c0106eda6bc1dce51c0c3248a4ed25f18650dee564b778b125ceda7b0a439fe0d45ea272f58f187b87061fafe267580f868677592aac4686fd10ec5a7d5bba04f0dd13943776a25bca470b55f245448ca059c7c697857b15c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f46fcf386a71760040448da26bf8516de2b35a94132dfa4ffbb305a84b36968cd852f085b346f8e91d0e9f15f8cfa9872a55c448a6c7020fb6b2b0e8c8a6086ef98d4c3ae53aba250eb045bec0e6116677bef15fdf869a68b71431421fe228adb789dc849e883475e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d9b38a43c5c2d185c58e55da9cca7959c02d56c610888b91411217df204687a5914ec75e2ca13901df02a564f6e28008afe8b87ae796b5ffe6b054fe0529b5350433c4b97388027c2afe6b570794e0ca8dd2e3c6624cc8685e4802a10de38e85478875d3ca9474f15;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e236f67abaed4d8ad564f3ddf712bf24eb6cace0cb1681f50f3aa619804d843646714af1a8317461e54475481c5617ff0caa0cca18a4f7f5bc3224a1abee054d53de118f3aff515e786090711521ffcfe42b455140689a76c0ce42029e82c2803de0fff62eda113854;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eeac6259ba878130979239529f9d2e2f302e38e8d1ac68ea657a235c498b710ca196dd2d56e858cae41cb29b3128137399f91681da53eb828d8efe5882d14dd586fcba409c2ecba5fbd9e5fafda5c994081c0e9c7fe34e6190010420f00f8d35b7e4fbf6e3c8fc20b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0958f3f26ce851bda75859396ea0cd6e8c8d82467a4d874102c514cc5a9d1649389ea91fa65449a820024d5817e101cd98f45149273f3ef456579be581dfaac478e33d215eaf3f47445663329fe96c510cbabbd9d9e46131ed93f832b50d52600f5bbfe6f136d9f6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1229d6c8c86ab0ca9c34ec66ac49903acb7930016bd1a70818bf522d73d2dab7f446b657117a68ffc7ff5c08f1e05e4750942e6dff57c4a227ff8ba9992da66a316c2b3b064b5dc145f74ef6600caef7dc8adfc60cd71f9a37723273ed57e966cafeb97e3b7c3a9b78b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c1a57dfcf118e335575955335e427bb04f9b850f26b416c9a21737208a83c06056a7b4c8c076dbc99ed42bac3224767c7a229e2d21193e4dd686f894077e3bb3952be19817cebbc1d7c74a732022e1a876d4b4e259d6b6815df706522805c53d1fb7857141bb3da9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1574d590fa20461379405c73e6ff6afdfd2edabfdee5752c79bcf3d0b89cc0436e9d1f4eefb25ee0c9b523322b85dbb7b8b3844fc49d3c2cd32ee60f0ceed622fe5cd60eeea88734c52b177a0365a3f9cdad3e59657c6d9e509b4505f300db88587e39e6655454a3d5d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb933bc0777287ccdc55b2089b8a730eca2d1e74a80dcff0300c6f10e029485a311547b2236a7427bdfc7b6c105409b664c7a05ab2d8877e90f370f4411d1ae27a98c838c2d2a1134d50fc93f81c1c95b6c1b9c6568279ebda67e63806143825535242b81818904628c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdce991a51168b5ee594b09dde9dbfc6d8512dd2bac5f7540abba561bcd31f1ab5d26b5d69dafc09e3a6788f935c8c0a2c55cb1fce99d3e7d2ce8343f75aee518a5c54393386eec6a41e5090f82134cae461d6fac0a0f5ee2c24981842f0f8c63349f2071116b13634;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c260de9a3767a099e5f33d08ad182c047e818a3d2ccd67133c96a9ca02f3d19ba8cb60723ced69a739857040c8e6eb762d303126cc14ca0be3332275a2683385902c9c8e894393a49f5751489380966e48527aaa620bc95ae2ba46887dcf869b78d754c5e32d77eef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h440cba8324a05bbf740d3738bbd7973cb6beaf35d7125099403cff415d3ca355b461de3f2e4647b32975069b935d97e8baf843c78e986fbe00af4e62041ecb1e234d7c3108ee71019f352d4a651726dc0158ba7eb2dffef708fa17d730ff8b704dfcf6a95a83ca1778;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bc28965dd1afd87901749a15dc775fbbb0e4c80b3a4b119c8baaa5c545ca15ce48b58552d0fc752d6b7ed92b40bee66977dc39c161cf4086dc7e93062b4eac14d06fd3cb2bb1b38edee8cd5fe8a97df4803cf4dab26835b54ca5f841afe57563d35960563baeee5bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3a7bbb8923c58a69241c7cb43325109b01ebf4b4e144ab9ee28322d4e96317ec5d11ee07b20f855787b191f21a66cfd4eab4f160159c935e61033f83be0610c57b21011760a09370cebc62ddb08015cc0f1a4df69ead027fbc2419008cc4ae5536f24b1a74b996fc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167f538f1ca3113aface5b6da832f557d59f0f6a54d78817b267e434b2add07b3988ef23afd92e89b765818be2c16a03270bac5b8716a41461a30708c0a6337954ee9a829ab63a0a95796346c7d25343365e52a6f0dfaf49c4c022ac2d22b8673f464150b9de0bba9ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee1e02fe366116d939fb2cc622e1b9a4a01951dd14328701934e1bc3caf4ee9b1add157fa00e39a6fee4897fe6ca71044e3f88ea50b9c2d61903ad50bc112b852e71048629e48b398e30d49218cf05e5527719171e7f7f08125c2169f3f7d7fe3146f56691dc987848;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe7b1454ca8a9e7b7bbd59886697f4c15531d359fbce7ca4fc043a35e2d37dbd95f50e6fe346042bfa9aab69bbe8d081d65cf5e959090963d13e9e411586a5cbef41b0e2608e204b7de23b582a190f249ec81588faddacf79939f8fa6a66af47406cd94987fa04a989;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha029c6c72c7f766dcf39768b21e0a87597910e38f0623f4143e922cc28ff4daa61d9e06afbc821977edf48535ef0328a441e399de1258a5d6bbd84b8ed7907e6e2bd1e575255cb2543179088483c92beb21b87b924871b308c1896efeee90660d60438ea333a175177;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bed48b144b93fa618c9bd460c6597d1b7e5021f08032af538741a1b7c0454a29fa9f8c166397e154adba07f23cfc046e9c6af067dd258a4a03439e84709f7fae4fba12c1b3b7552d7876cd670f7bf1cde44dd349325d61b88c88a638782d5a8a4d237edd8df7555e42;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13445c0948bf07a2c44e55a5c36e95d4f8bbfcb1cc509bc709dad328974eb1b831cf383b384900ef1313653c07a561253a389e02b2644f0c7182da16a475f8a258a81a985b5e5371d3ac200a2cc2892d4c9193c6219aa04b9797c5d3a5d71113fe9dc40e50310099b20;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1202549c7d113b90b905fb02810b3e848e3472897bcaf43df4da812cf1bd4426b054747d6a9c3213d31be591a63217e919cc8ccd95d8939b4b69a9de146fad24809c387c305c87300376c2e4e837ce22b300c241be578b8a5982f8a7bd1453871c49ae8806ec2c5ead0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c183c1f353d3e176bff67af0cecbe074f7d690ecf64e63703fa98bced11551d9b1597f83f13e63dd3fdfe47ab077ef857f20f49350f6a54920b7dc60161b5ba3efab3a8c0342b46661fe9fa3d581eb21a734dc1701274b54b37516bcd3add9450d7df4b84556aea07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'head5df8b5800a657578280a0b656577304b3ed4655bc68c27aaf4600e8f457290861a060355b9916688d5176118fb9a4359d21b3a64efab095aa281381561c5d9c72c6b0e2be10fabe50c0b1a7c44756c425f39cbc789b9de67767dd8721b3a4f0ce8e35cbbdc3e9f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b655fc737c1135b0e7a143facc7e6ca1b8e3a09466045b703a104606b1c0f082937c275fe46070678adafb64305a7b7d5f069ef3392dc3c707873acdc7ebea5cd104cce5cda284039781eeeed434b7480957c1a3adf58ee8ff894d84b23ff64484b32e5639c2b5398;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e68ec0734b4715fd89c79e0fc0448513d66b5ff920812e4781bba59618561c2ce626cef50520e1ba9c9a036faee720413189bcdf210562f50d5c2c7a5829f80b81e7a1fe7d2a356828092395848e2617666cfa2746f7aa468509ad7099d0d6a86fc0f5aeeae579be27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hece0bdc496a3dcc7a963877607631a0cf0913135125863b656e2ad07ab72e9247a82d0d61536ad64721383a91a390bc4f17cc3fd4c7784a1b3284919f0946c3507eb40cda17df36f34c8efe2c569fb95641d08b59d4b9d49ca85a89a3ff81ab3a87b9d9ef5a9168265;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66c78f05e50b55ffdb9a0399c521c78372ee52ffedc36119c5288f2242f7766eb82fa3470f012420d1c8d5cf76cc52cd67615264f7e4b148aae8bb7d145bb426ed71b2dbdf88e49830ff8df66e16ec55f1daf9224c02b86b9208d353d248b9878b38ba962358363a28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a9217bf9cbc394080d4dbaf68df71ecdc3121eb0872fb948a766c6177090f4166438a7b5e9afa09b27695278d3f9fad5fe2fe12b988fc8705422523386946e572029396db039a395df2cbe97b864483655cc14cc0de8b255dbd833be87e0503bb8977b5098dfb8a51;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h248ee4edb6ba4e388dd290270b60c7c8c4f86afdb563116d9ce45c33e849f100fb4f02fb938fd236a1a458c6ef0012ae0ec855707c89af9c315e2ecb49bfaf93e3969148dbe3cdbc30d9aea62e6a67ee9498c37a0ce6270679d0f05bc9b0878875a0988ec27b904e5f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbd47644e9e9183f69a95b4dc75d96276a9b8f56dc3c29868196728efb812d5cadd7ccf981920cc6a5972e0d681d59a5e21853ad7eb3ff1ba8cc7f7b2f88c46d32e896131ddd4bc5a377fe083f3cb2083b191f82177ab1312da3c887730b5348a9d9934d6a1ff7dc37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13490921dc009ac6cce0d61f38722c8f15fa29d18f852584224b4cd8276aaab6ddc2b079e39fb23209f806f6eaec600e5fa20b5c6c37086a8e8a649f715c782dc72a7969947fbfe558f6e556085bc1fb2813d6fb4465e59d5247e6250c929c33934911f867c143f9ad8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10096d31130cdaef11f4647b7c7340f97df3f955cd52f486a38736e8853fff0794ae2617b94a148778447df8e3cf501b3abdef55d97327cb54a183e3360635e7df4f39bb8ca5077a508d9b8ba550d9040ba44266e3dd8513d60a27dcd43eb772eb3914262aeda2cd15f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103248f2fa89fce9012452cc6d671111cf2e06e770d9ff06758ca65821e6cae4d9dd70c07a1ad070abda381820bfbd0ba1ac803a047b3143e319f7420c8f5bbe179076b8d72af87b8ba00209319c6f1056c9d60c170f5613e36371877746cd5d4b91012b34700f7e602;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac22e4e105185ab6c95898339ef3305e331d067201f8e3f756c3e5556eec9f475b83f8da1683eed39778003bb931fa3200a6555059d3e3a98d3b0b7c3f85988c064ac9ccbcde6220d3bde909872841a6b3b9ecf053d5a2991176b88a22b3474eb641e2215c8fcc9a0f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e924b891b28473c936b3ec2c973e5ce272d61e5d260204b0e630d78f3c1ffa3560dac93312d98d7292574d4c3a86929c132eba7cf62187775961819ce4c3ffe2859d8e56a27c908f2dbeaef152fddd93453ef0bcbc0dff2dd84ca903ea39f07a9e4c7699510a0eff7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9bcaa9eeb3aaff37285688b9a889f4e767cb217bf6fad8a63a7a540a815a6c399e6ed85a13f9cd4ce3b02cecab6ed0fa08b438c9a55c2e859060cf55d2eac93b152ed1d563b33d8be7a2a7e92935f110188b2bc5b92f0456f983ccdd24f7a09ea9ef54263057f2105b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h110a66552d57d75742ebf88c741126f210275ffd9e25aaebd07f9f63d9e48081a5d50cad495df5ad390709c3c9693d2d6807be1f5a3896aa43054d2c4369334a12141276521513c51ec396f2819935440e1bd3dfce8e4a72484b9b3aacd63f966ed0dd08e51eec347f8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b5c7f84fc0bf3ab08c24c8882f147dda538d75a899f9be3b40f58291a6446e850e3abc794db35cbf28ebe0e0233bd86c049ee997c86c0806cf21e04d52584877520dfbb008428e50b871e45e14e04de92ce551634d0f0cf03862da31b96c03886795f43914fd1e570;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7e1d94bc67a323bf6b4259a7844f9bc5fb21ec4f2bb18f57b4a49af2d12ba140774b7496b45dd6dd0dec42e163eb998606430922ee9962d086a169af6ae9c99f6da68e9b0ac809043964470779eac1a29c821e05ac2a56c627a0f45a918fb0c9495f39a5fbbfb2aa2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6a039689ee2348a04acd1ddc260609b50f234cc6b7a44b43397abcddb7105038804686fad9a655bf2b02a730f798822a141780f9c7472eedcf579d560ca6f61548c7c4eab024c30bfb5377fcda6ec904ed1f0301584b83e74352bf51cc14a584a91e36e28e2f07b14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b04624e46aabebe0ce6a3f54fc5f7581b7e1cb250bce3a11d5180d9b242963020496e5417507365df465f7a3ea162d985f0217054098607844ff739432bf5852522f4b83831125c8e3f06d0d4b908e1e2a13f7439effa4e57b42dd849365f28f073c048209c8b4367;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1158872263adab3f307c7aad47961fc811137f2677aa7b1cfd1e9cf3feb02fe1c06165dd88e12883c0e33aabd955b8f69c64432b4280c17816dd8cf9e86a15833ecb4cb9ec6a8c85bdfbd5187ef7f5c4e723ccf39007803d1583dd550829efd60a4c240f654d3c3dde3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16331bcea68e321d4d64c7e6d8c97fdd432c7e15274d48ed6f633a59b8dbb67e57ee4dd2172ecb5a2f8e2f0b1320791195fa84b61d8b9df7bfc12bf0557137f59ed1940f07b91d7c781b75fff2469f10fea77299cdfc6dfb036791eba0fb2909c8b968d7d8952035555;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118b1e21fa817b42b82c1120207257652b7acd48e2c712c0ed74432c24a0cd200bb1b9a23e0813076d54d452b14278d1589a065ef36ec84334577b32c6c5734bf0119e0d88aceda84c0e259d9f40a2b8cb342e051ed3e6b28ff1762ab0cfe418bde6e755fc8eec9bc1f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae6290cf7df15997071ee5ed8a6e8a757d17ddaf19c266b27998efddb1a93800423a9e18997a5d4e09e88fff9c83a16526bb267a82f9118a2a04fcce1cd2f52680c3860f2970616eaa08ba192170e21e3421983660007d0367b59ab8919efaf26231ae469f8142882e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec2f3be9f1f5b9895ca158c82be933588792d2c12889699c049fa442ecea526aa373254c4cff6269524fdadbca8b14de2d620e8bdaabaf246aa0e7876a94cc074d3bce7672869bc070f8ea87d5090ad71b08c91100fa71f75f81246ca93406df70d4b9910b7fed962a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h851b0c57685250c922d8ffd65c811681a271b40b1db9ee4e1d4406615d25f09970024949cbce767e59ec6cd9e9c5fd8fbb665a38476b7a17d1aa73f892df5d2054ded980698df219b7d9bc54d5fa995abeacf697330115ddef85e61283ca08ccd89e14abc855abdfeb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e6a76a9b394ae425e84c41e1a403dacc0376772a9400f905fb8b65de4ea8e1dafe8dd713dbf13ac6e18499f3c91cfe6886ea00fb98bf4a12ef71492979199a48e6f3c449e41d90b4c1c6e859c4b9be1f4432885c33dd361ba4b20938b9e90cfaadd24f7d65e2fbca2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dfa1675cb995d749ed3480a14988f9ec17de3fac6025ae7da0b95d57dee88b0f7a635f719128d16a9ad9a57bc1899f9152cab3b4c2d55f1de1f19ce7b0e5b476265e0e175e9912bb1f18df75fba3158c13392adac7c05191d43a7858ca7ca316fdc2a335003611fed0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3078111a9f4b09dd4abb84fcf54aa8b68cd416b2e8f7f16e0072d582888cfa25e81dd8c6e14e9c36fece57d9bcc9b833e291ef7fb78d228368441d17e974caca9ab5becf81c578b6e7c394194ed62d82a1d68e53824ef58233ff2d4513fda0e00267302e9d2170946c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d4854d73772a2249584c8419e31fdede56af92aa4d2197be57b17b9f5b86eabf46abd223cf4bda4da5c6e59289b674a83e280143d420e26d702e1a61c6ca187829251df6c3aba68c871aa3e2b8b414928931c09f4b103eda8ce3847b3ec5a6196da55b482bef706cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130a9f43d6179563c413b8f31ab3eb7e175f6d9a64d76829b904fd195e50a7fd6cf99f35e7c9d352a302414808b262cb48dfc063c139708473041a0385df2d34136dadb8261cf996d875c9f5749d05444019c8308ac0944f28f14e09aa61ba1f8fb46151db3a4d19747;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a94404aea638e8108453215c1642540f22a997b61fabf691efa6452d58a93337c8bf05b311f857e3fd540aa946b5dbe7a1fce321d375e5a0b77b5029f4bf1e273055a6b6e4734ce322a62e522b9964a945929313b05c9220f7edd65c19c196d48732afefdfa579ff7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14aa7ff407ee6ff35475a7bdbd3c28a51e9bca830fb16b9f9925cb2baceef150dc3794c4389a1b6b40b51b9d13b54c64dd72f05d7ada95f2ab331117e1320bd3c36983dc652e38221d4fca8fda89082f303c3257fe53617f54571220d9910616173d409f4eb8473e6ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca8db256a2393c4ccc5393a8e8b87b5d51f5c7aa62673113fc845986d68e30437c4e8bf9b66e1b14e3b708262ab2c97306cc68c350e5fa11b8b49f50e03ccaae253de64a44a3b02571ccad6a5e56d1556bdaefacab6f37e7c190f356f8752ee238a893e24503a03ec0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc51aed80343d7e70a2c9d980424a7a1e010620eeb875b305a89b731096685d169a3fe88fe0b7ba57b61914f6b786688148d6d5e213af74c5f22519e4e0df0b1ab8d52ba1b7e5e7c80ddfb395fcced8d154f6c53d164cad6b67aa3caed23faf13e2d8d4398fc8cc91df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177739344e10e00b652db0857d26381fe951319cc6a9c45d867203084f0ebcefa45b7b03136fb3a5a43739ab5cc7c03ad0d63ef7f3c4da395399776020fa11005f4c63f5bebfaf5f7f534f2679e551b116c44683dc2605480cbb3ee3d80268d822c7cc9343e641d93f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169c7c7333f5917db0d165108030dbb3be665e05da68eede5c0f2db28c74d75cd5170977bd0da691ec9c176b310ba156ab898dcec5e77973f62815cd853d3000adea0961d965cac585e48bdd811824de5a8a45347fbec11f9c2935a87015a2c92502609429738e8fe9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h224ef8c13c43d3ae0fcbe375dce91aa1842eddcabf74c457ca29bd68143a8a8f9456de86e53ef4d354f45a55dcd321770aa3693bff67ca4bc51d63392c999b4d47097adf74e75e81481125f30a5e91b5c49327d1b0c408f26c571bb0cc547d184a6d250adcd410fe76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14209ebaba1b41b9fb94ea8c219bd81c08620674328b6d7b3ea94ddaaf431560bd08b65ecc56047e59925a537ac9d13a6bec97446828e963f52d2b4c887a48df209b64811ae51417ae8dd7209979deb0347b19ff9d69194bd596d42c0f4727c7ae17cbed2504d53b0e8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5d2adac81533703987d0230aedc078dc9e77676ae4300e3867ed6862f1c438361793fc8f10628c3013f26c8fa89f5aeb6a4f81cf0e923486fa1538a87bf592e9777b39a9d7fd111e775fb64aa5f695726849f8307d188d0df3a2e53b7d56d499b0811cfa8200d2341;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2cfb2f38532d94489d7bb6fcd3630faeb8bcd1d29457e297d32ff6e66a24c076086136cf1dc6283dee05bc0daa539cd63daf3c69b67ceba3ea29f537b77bd8eca230638ad3e186ccb40030c9bd1340fc8f4ba283fa8a2b892d5ed01d20b3ca57396d83bb89d157d183;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd912bf4158338af553ddc03670aa0c304323ea4dcd2e3500c27a9ca4406bfd0c2c904e20abb9034d09f5f38e37c54a9ce83e59a9a825993a4d3674833e9b70f739c33a4478b081eaeb811dad7a3a811231a2667415802231f2a85dea2a21c7335a3c5f908e4d4d345a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7492d55703f27e0d402a2cb0c59b709f12b2113f062fc04a92b6f280822180bd7396120c8e3635868c10791f0f658c0afb127aee2e63f5e54f4dbf48b9971f9c3d81127c210962626b918acebc9fff8038db086ee816853a67313f9c65b269036e4b83b5ebeb33131;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbab2f390b3a25e8c330b8d85a0e4f1e38860f4772dddef2efdd02158f5e7d8209cd4bac19d459cb501470ae49788a4357a56636fdf7e7e2434e25b97b73288f330414c8615db212d983a4f38db543ae1e6a1dd3001659d1569b5cf81b671805505feda6fcd9ab090cb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1913fb08ceecae288d5a148d213338802182a037292745f1139eb238406b5780fe67b2a7cef05c98210f26d1f10244506193859f0075710f7f80c7cf22250e2449284591dea1af5e7a060e48e18a7f81b5514bcf5dc4776576e3c786fd688ce454373650fac6cb14d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bc7149d2c5f8bb253e128e5b013163704bf9ea0eef03fcfbfc48e662c32c17de88fd0aed5250631245e09842b8a1369275a08b2fa4f8b930ffa5dcea0e0e7f3e99a52f504dab83ca7fd2a81ae6ad5d4a19b65795e8daf0f041c75549ea0b77fe3bf01e7d1bf63cfc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2363c09141ee55a20dafb88163d88e5da5917680bc7a33429113381c208f3c9264224f0bb34297982839f94ae8e1e1ff5bf361dd4e0d067be9b3a84b0ce212cce42db3860358cf6517c555c770ade69d1f46c920f8f0a76628fef351dd7d2b046b7fda1cea8cab57ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9dca5616448a2ed04e4275f43b3f6aa4607a54f0c9cffe02e3c720d54605d3275a442a8fcf992213c837ec4a4404ed484fc8abee34156a986e46e9a3419933ee1d62245771302139dabc405ff4e8a6a22a5cf0b570d03ef3a30b74b1e63bb761615068375be927f0a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ba593642cc0508922e39812516990551cb59b00b732e65d0619306ba551769baf370ca7bb9c7465a00847cb79fef83900435435de160ec9e6ee31384dc8b47a5152dd23368e29602eb736455d39219fa00e14e0f7cb4f9dc6e093e4ba56e0586e45253eb9ad9fa731;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ea26d16eec27024e3818c626acb94511bff685a531626fc92ca05d1e206101b335cf21896969ad7c4b2348cf621b1cc753e775c63023cf73e05b2676492c3349aaeaeb445db33de6dafab2414c54017dd9c325597b64c97f9ef709c80a19c4ac10e235af76d3dc5a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82ceee91ca41682342dcf26678c570d5af05ec8022bba64a0f8de07106cd70bc813e183a853a4a9e34ba186b54c9e860fb48ebc7b24838d1e001630529612daea11cfdd737d76713e0348e87d3d2bedaaa89c3178a2e9748366693520dabd97ead0f2e918cd89173e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h495885d9f3f54efd51a950385637f5b077cad6d0549f062e75e09109427866514ccee22644e2402b1f2975eee98c032919f2bc49ca4738f95e618a882b25cffb4c2c1e0e59ab186bcea38fe55c98012d8670e283e803b00fec61606889e417e9b0f28887b8fed68233;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84dd0386115e802a6a1685adc51500bc4690f77b5a360489dce3df619e9f74e3b3d747ffa68d647920406772b1a0787e9a9851a3d6cd6bb59b494415398fa6df4c556cc39e576d9adaaab72c143c557211dd728dd678187e6271efec35c8614ee64b25e163c4b02ea8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1355a57c23acaf53557dd2b37e82b3b4b1eef0cec480b4b99eb7f8424debc81677b20428ad2972c66a8e7202f0d78d01a76fe01c136f962b20aa8b5b39c9c294cb9d92e605fc06fb6655a2a4e7df5df146190b4190f0d8950dc3fc517240dfb8033d500ebb34b4c5dde;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1e5611f8b0554b54a7315e5f9fe88855bdf1ebebfadae1e2942298a727e10e240d523a7889d45b3f0af51a70a97ca161623f7bc05670d948d70b9e07456ba17053ecab39c841d9fc194360d7313efb4bb94335dcd0c096203812dfe0ae148e83d262662d1a78d9cf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h708c28647fa1cc4ecc4712cb46c8988bfed687f4f9faf733ec20bb973c5d3de348240f62fbae58a4c7ca122ce2ea9d0345ad87b71ca84b63172fec7c7901da739a357fbcded90821e822142359e87d84ad51b0bd80c6317176193e1b6bb05565df233a7dd7691dd5a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183fb4ad42d35b3468b326ee05411740a0826a7cd64887f977f366f39149ef783a012768c1bb0c6d8afab6a39830f8892e8fe00f61684941768d90b1bdae9793ae0c5e0b52d134b4de9920ee7944b53936c378bc5bf6f977a853070f573c64d002bfd1a50ab02fb6715;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77f439486b0180d20f69c4a4e081c19003220cb40d1c0213b7128419bedd0e684d090b869a6723d1d404d8a58ea495e17a73d66405739cce406fc034e3bea0798310c4d66b7e5a268498d8c317ea1654e5f4a946d0fdf9b46b44dd12c6e0cdc3dbb5776ab32e79ba2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bad6d35ef925a8189e329ac257d1c8a9b7d917d82892f370ec7682a90627cb4a998ff7eedbb1492c414201f3e1849711d03b65282c0e2124ea15e1e360bb573fc28fc5c2d76f8bca106850c3252627b0d04551dacc64f10261967ea1bdfb4f2c198b21ad872ae07bc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1553aa9fa9adbce047b3dbf518b3af5c96915efcd6acb8d6d52ff3fb4104284c22a47e413ffa9b9ad5ddbcb044d4a9250f27b6586b364e08056d7ccf4dcdaf044610b6b04ff6b4a182e114f5ef93c67c73509770d05d45a6c60028e56f4035601eb58fdb7e9c7817a8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a35e5caedca0d4f9df8bd164534ced91bcc7f178e05fdb3650a4ac945bf1a302c2eaef73b9c649559a314932a476d66979d79db9c7c6c846814ef6ad45ca811e4ec826bae3f84938ec0ab10edb8dde7f5cc45db42eef633f594d315f9d033b1fcf88e08a73540c025;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153878ea5064a99651b8da35430fe22f7310961a1fc79d36e10c5bb5f8cfde25dc800fa8d9d748b0ce4b58a862bf0c9923457c664b2dfedfb30eca0feda4f9c43541f91ab2e43be1456e3a07a11583e4a6a90f3fde49e5034fd0c9e4d89f311582cb9f9bdae44bbcf09;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a36ad93c739f28063e17587a4b1cb4b8962825f8408f176bd5b8d1a2c734c571391c221f5a90df7fb92ac6e3e6dfa889761484efb3e91ad6b3845eda84b7c14209b626a7ef26bddf64d2cf84f6a0b07d31cffc028fbe13952fd68a7239e9a302e942905df7f194da64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51675fbc2c221886f4234852575f2252c03aa48bfe16f4d312fa2d45b46a1bfe1017bf1aa60bc009f7c1da615363f051972d9e4546cec7f04e5759f73e5fc5f73f38941b32aaf32e84f341f4c5db9b1c4e490485c1ba7c48de53380f59702357153f8b23f47183339d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1228b2d73c4f479524a6dd7e57cbe72d0c403d9921ba35c72f37d944e4ac4101fd81667c4da332add0de7193f81463ed90291801163be3bb982b38008ef7206ed791b22a6966b2b5d5678380febf8156a6c0260e0b2bb9e8ffe0f5139502797d8aef5d047bacad1ddf9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bf0dc4dea24d107bb0947931ba84dd6e97b7ee38a1c65c2a57cd0d5b5e8c53ea5363f78c8d5fc2957c5cee1e1875fec8ca6b4eb9f3df81143e9493b11c5a1346e4b97e92cfd32ce2be2c615ef4c216943471d462d274a00143ab6d3a2c65f50cdbff66b88d92fd389;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1149188ac38c98662323078585d2f7c14c5da6ce156997668030bb7773d3219f13dd6db60c5e64e797941c822435582d948c01897c16bf667cb5b4783225c8aad8b817b05e1f60230e21072cc824cb5b4a32748de5b47c10a90c6bf85e76988672752720b3c88d0f64e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha60df5a52747e2a24bbf28fc0d792d101ac5a04d78eca68772c4453d19bbef0cf179862c6c093419b0e136378fdcf89ce70a2491bba595d285a3e9dc3e0c71e1d210e242d063f71b3a6bfc39a9692ed7bbdf23f21442095eccbfed0652a1ceef9d8d7162feea66ad3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51f8954c24821e3e5d54b2dd79d63f1a7c4979de2702a18d26804aa4f51f5f2769f056fccee2763d4942d4b5485f2ee79beaa8cf3ee4562bf2721d9565f2b0687beef73a2ea9f1a83e56e2381df988b001a7cc70bcecadf959f4bfc96b631c1f651e3fa896c1e4bf79;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d70cc94d155698fce2bbfae441ca4ab509ecbf5f747360be9d9ace06a6940df19edd78bf7252415a124ebb14689776f51c1f3f374d025ad407d7acbe4175d04a2d65d20a6d35cfa7918b6622badcdbd58146efa7803f3d037c9586cd38f5565dc4f72bceeee796346a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffad5009776698276a9783806966baaee7d3ef93b6558eef3a76948a44bafad689e0f763bda09ba8516ad92e8e8ad6b8a6a2cc0df9cdb5bfb15f51249a5d306da50975ae7979d88847e8f631476137b63356262e224299a03678f189b167f90a827be2a53c59d03211;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b5da6b3981c88c6446cfb70471463687e99d0729a0c76f6ef72b3b8e71bb090e51a4242d069520aa94eda3036f34d39f290d5d7a273ab6e52894fa99aee6adba210db3ff4812ea9a0f8244e3f85386cc873f18c5ecd0c437f5922a62a196d4601675b918e018d169;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15aef19ed3aed701c8d64ed588400b093d3adb8c4a01e4771c69da0b7e847c508bdb869798beb5e4db466f20bb3c0e723d6e3c8da7ef71bc642e74e2b630aea743d96bb5e52ee45dd01abc55ba1906b1a1423a5d43f4f91f9b7e79fb98c573bf96cfd42a3accb6fe9d8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h402c54d9caaa3801b111108c0c7001a6d9f03081990a9222a0dae163f8b0588e44b41600ebe73effcabe34b19b05db4514049cd60b9ebc49b41e82ae0cab4f383130332df4e7592b2d9504f295c98367a0f0d3714e86a8a427e506ff9fcdfeedb10d99f174b73fe80d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14335c54591f684a07844ba2f68c0ff26b281b7a86c7c0f718cf49eb4bbf263d9545d3ffdebe6c97a7f805d159e1484b84e337528141b85c7f0367fd2d20bafefb8c2e1f5ad1a6934c8d82bc6aac0a0d82a8b577ef33d54cec532f77e3c7e97fd3df564202af101d4dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c4b940329849e4b80d8c4fc42b0fb8fc8d5e4d7c534d67e7f18e4cb17da5df9e51f20e9a4899c7d2fb6bb3e10697c7274026c5ecdc75c6fe32ba616bd8d03a6398583d37a2159b302da7396071ebe8e83bcd544578ffc20f048f5048ebd62e37d2037633acf072ec5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3ef382ad0aaa85ab4a863c6aff3614cb655c25b7837e8e4f1a741d91da8b7ae53456d05dbc4c8dded1bc95018d5ebee95f91bde1a6f613772da423a677f169c57af1c7904179a5dc467d5da9de4a52842ba4f5dc9f817c50c4de81b1f0fa9358f2ad7c201f665db64;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7f0583e598d89478189288b9750a163765804af9c36b06049d1d742b0d1282ab3de58850ba54bddcc0f7a836182df2608dc0e887988b0c33390d79e91e5014204a8ae635090b7e0fc3148387e418cb18a29549ed45f87b094efa06ef8b9a83a50e183ab778558d743;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbef9d1b8a892d247995b1a1a2d48241ee9be64346aa9a7daeaec0f004f7eb6b83b30e2f43f379260390894563e6730050d88e8b7eb9467984cedd09609e674c122e9bdafbcdd229d7c979462664279234bc708d14ba72b6ef98fdeac0df60d73e7558ce71638ce9ef9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha158822f61210a4864d35165d59ead9cb8fb78355d44d15ef1393914fe80fdf74e61464b8a80fe2775ee32f200cda0e0217c366f59d51261d861071405e2ce8df075170a370732e3e4c088864aadd5c0416a5179b7c26ee00c523f2edf22b3eae0896a02d89b27fd76;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f3b211491b302ce9fa83805d9392d2fd5a444070ce58ca2c60634315e99265b09666250ddc7333cc23d0bbbc05bf6908533d92552495984605cbb6f33f75ef7cc45db52d38a9e6285481e5b3b3117038609e05ab8dcc0d6cc4a6711e358edc17523f79c2fa9b3e723;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d881010f9e52f142073f443ab2e44749830941cc49e9042c7746832400c7bbc1b76f91f439f0fe6a9fe8d20d363c261a9078da15d1d4ac7e33314309b940a8b95db5683dfbc8123d3fb1421834bc773e0a750b81f0212eaab63f8a8247c495b79fdff2f90606450e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa7c597069ad2dfb9955535bd780203362546984bbd1ed14f3d039f3a9d289e663eaa599cb24f4cda2fbe6127509235dd62591dfef574ca479234877a0df3fcd542f32faf3982a92dd3fe0b6c2636ea6baf3a30863edfefe53483e2d31b330e67c6a8bd664754f2e8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ae4d2780b879ac30330c7e2279f967c297c46fd65c50d47ca4ab7a5e91bdeb261de84441a60d521347bb951bf9810c104b74db5b34317535c5e14353f926e66938977fb22522e5e1d5fca929e677b068e60ba2da4d0e44e76431f42719cf591f094f6ae328ce525dc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c6162a6768cc41eaa7dce8f221255f263510163525d3a894d9e015d639e712dd1d1bf136bbfed7245f62d8c319861b9a02af6f8ab80ec5b2306410c21802359993affa3652082d7700e639b8a9910146566eb5cf220fc1b07a65053fb6aa55e3f657b96869f46f098;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e43c5f966ad165caf65a45ee6078b46f5a1abc4797b31998f9a8845d41a20abe9f5d1a68e8bbd836e5bebc7b8ca28a615ca0a1e05c2f19edd9aabbccb910b2692514502f0cf0bf35973eb02947278e543c0732faf3133514f92d90111c28b6aceca813210a832d2ef2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba2017dc5b61aa54034931d13c13fdcd7d1950260284f8ce912849e86d08fe844bcc223627fd0225d26b7fddf56df60e2b5f4b5e048fe027d8be4b6242b4764132e2af266fec33b64e1335d5762f48aa4ad0167decbed2eceb024a929a1985ca4dcab95d7a69fb91b2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116b219438cc23512e3ecb0cdc46afbbe5f7ac1b3d1355745fcc7c708b8427c5dc80bd2c829200d93ca2b41895c6f0023f1c627b75af7c8c4f9f50d06c7fb432997fd755176f9e366eae6bf46e8bf8e60fb559d516e8075353b7cc4a843c4276d1c762a62696205a15a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61ed72b95e1a81f0a49e4d90b531b812f8f9a94a8cea49f38859ba975cfd59af5a091f841c911f141147daca236d837fbbd0fe6c49c07e4a8e0cb7933dcea9989a0bd8dfd9354a292a915ac4030d9bef8007af98cd00b0f5549f7dcc0f4ac66019e46694f3459166c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f2b06b2adde16f6629b82835b488b1fe82f368c587634a5860aee2a33c407e6bf1f267d267108775af9b4782fe910789c37fb3d051fefd994ab829561c0bdaacf4a07680d7a7543820c97589d1bdc47d3f35f732cc35ef735e6de310e1faa42f9a37fa7d1c2594c73;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2e02685aa758b8819f77d65cc8b1704e82c349d0ef1705c1e38035f1cf6170d37da587e0bb5d27f6b4bba801b8a45d9acb3a9c0cca4f36ab8ecfb3c2348eef70b1d598a34628d5b71e2e105dcfffbdceda55c8659efef1172852b37f4e076feadd183e07b72cd960c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he0bead6db100900c7ab6aac491729ab81a75314926b86c2bbb77250c2cd1c0f30216514c7dfe6de6372771346c1a6208bba275aa6e5f7feffe0fd97561e87ce18ede4a1469b8cf1db0e4de354290c220171b5f70e593e09e2c5339c65a11275cae6050ff8a80c3fe25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18db9431c5a05548ac40d88067c84cc2605e85aa282dbe85198481eca4c76877e247ad4483079a553d98e6f4483ddff62106c992433549853da20746d902eea5fd2e9f930c1a843fed615eb23205c81ceb0bdc0bf29e3b0844437df4a770ee6ee33524e2cb8f0089e3c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c6232185263a5ccb8687b34c531856fd90ee1aba764a4108f780a8281b87a3251b14d893baa81741718712f1fdf0652db82c2fb3ba68d17283b14d0e7e3c3b159f2f949948f84528395075abf11fab286c1c877cff9d00cb49cbf109653143f938f3f87ed9da5b63f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4aa15ec64cd3fd263ee435adb025bf5d6e4926aa68326d946738a96bfed0fbc5cb264bda2de4fd1672a418bfa12747d8c3e20063e51083b57ad0e5fb202c5e232b1929f144dbcf2a9f451312cb3792b856aee9593dec0574d65209d3fff180220cfa6021a99e0a511a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141f43f977cb361b64a729ade538eb320eb8bbb81fb6f6d07a73371f937d517b95160ac0102353644625224e4cdf081912ff0af1f4259d9d11420198bd54c83bd583be4a8624606aedac1c999ce590aa710f5a3dc898e664791ed5b36fdd6ee2dd44a6aa2daea13cf1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3ce6838d61dda42883f774f27f2b2f982b1fb58a2840c297527a2db8d8974ff8c80f5b5961da9532c11c4ad0e0f3518908334e8f3d3290ec77b51f7d34681259dab476a3dedda4072448242407bd2dd90330dec108d6d29819b3677050c38323856749d4975ce7b9d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bd2878282178ffa098e41d184803657fab49a0f49eaca9e0534a3f58eba96dc7353555dc10c0375381574e86e6a800a6619c9f867a5ab76977e1da00c7771f75cf3fdf54215adf0e4d132e86e9bb19f1cee5566cd7f016cf667231442916f5f471ea87ce89f64bfe2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc92c1d797c9a8f698524051a2f2054eb70925b24d811fd34f10fa0572029437b621431e6e7d5e68b20107e528b5aed3de95a1f2fcc84f6c5292c2ff7afd4817e0998bdd0992d275f46f2cf4ea5e79b3ddd0d12c8f50dc0766118055a93faf4a567a0ba454b7950b9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd6d978d2deda34ac694a9c2ca05b76e79a6670dbc0833e94d2d2b35820a598cb2ebe0b7e09bd4f2df88ad5c47ec80c5557277cef9c88561c1c3129442e891d2d76a325f38a0a3338a73d8627786e164bc0fc6ff4f5d6f0fa993744362f6cbd3eea79e0f9c33487029;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he25bf8ef6d6c875f3aad92cce6a0349ef686a59776d4e1906fc578ddeb9510a12ec66df14892bf783fb8dfd5df383db07b09e30fa0c33ddc71f3c9f83b63524c09b02809c9ebfb2a8c65efb0cb7dfe742b068966c7775de05810ef01efe7ca0279204ac097f83b858b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6d2f05fe681651f53492cc19fac97060ab87048a067570f73d3383c64439d5ab523ceedf74947c6f93902a97acd24d9943e394578397fba840258f11b1d839308565b78a809dc0328f9703a53f7a0fee2bd19d3385899f9e96d55860b567c7496984c14a852c99355;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8f96aeb7f39604786a25b3bfab1797484eaa603a2c64c3121a636724f2e15ac27165854734d33376008507afa176bbca5895e62b8ed13d281e980bd083b5f751320ce9bce985e0d69968f364646628db9fad267081e52e368ef5e5ab193b7b2d54c59ca83316c8fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he286e41868afdda9f05aab2d1ba29a6aae718c073df3a4819da82f2e9d8d348c386cc599421f878294b559792ceb4d547b8b610e55aa53e0e92244ae21439b99f005867d3086f510993c5472fc525a6f511558bfce654f6c03da77a14958d4e65422e0a173f25ceeff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc5d19fce2fc3a4b5adc9e80c3354226d0789d74f9ba0048dbfcf3ab74b180d8adc750d083a314486eb20c86bc56adbeea96787d637a96e05984ad50e8accbf70989e504716c60c7c84f5c699c41cbde9b4167d5dee81226a215ed5dcc802e619f3a99828d875b1598;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66aead8679b58dfcc7b05224ccb56362ada466e19484a1bc945910e8502184c6b6a294c96a3d27204001c21575f2a36ac1c0e8f7fcbe3efa49a45a266ef6454eceba5e85e027c9c521aa46b17f8df6e3d22ae27fa7d4cf53684d121e6d6279c06ba2d871ad31058537;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h281e374af4e59cb9211f5d61881b5011ea246e6810a8bea4854bf0a20ae2cea3c31c5b4aae7fd07958ae3e384272aa3643c86c51aa052c8878b5e711c05988eb3654d435cd234b1a673190e11bd7942fe06c01754efe4cfd44148e69d95358ee05d6fabc7574b18548;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec9e85f494f56e250d4bd1e2b096747f097afcf3beaac634c581907ca620935e990cb7ae92db3c4c73652c9427964f23196cb6156e5911cf6897dd7e1b9ce5ea1842a5ceeceeeca19b196644ad01ba7dd72b0630ae02f24bb6a9ce629f1932bace86b941b7149eb448;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14938f0c93b106a98a610f6fb03cd6c277e9847b0df6a459fffc5ed86645776620dcef40c194d7dc7c40764c6de3304726d71e9133879b0dfe561e71a6b2ae745faf29a1aad57285b6988597bfbb64c19a574949d663b8e072de799039b472b9c4ccc947dc047b03d57;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1ae15bc4ba569582c9002c30eef75a1e78f0aea57629f30449550803b4b5fb1bc320384c7ed547979583686b2d66b575eb0049751fa3963bd27a3e2038a57d45c4cea3e139a6e5e835caa97ad00ff836df085dacf480d0e599a1bd51c8b79053e9d3092fa9862dd74;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb060097676ef7dc15c73e43e9e151905db35666168929e3ae28741e683c123b7bf284f6bbb65db6024e344be7a5ceb60f3a17be9158654a21bd6878e25915b344d03aba8fb66430d8718e1ea162911faaaf7a2bba06444660472709436714844e8ca1fe978e669e0c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14dc0e7f5c553beaf36f60b25099dd89ce0a384e34d641b950d6ad307c1bbd0c0e27ef074375c4b3002abc478bc31a37c3c8e17662f47d1b281b99787ab01cfa5a273c05cb89ce642a5088457a2f10714eaaabe7ae7c17c0f2d5fced65eaadaf3e160f7e49ca351ae99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a9c23c18e9581327d8414f1249bdfcb4affa870376f0e8e7b375ece9dce790be7ff2f5edebfa24afc9a92297ce147ccd8563d625876cc7855b90f08c5bbd238cc88e3d867ff012e1cd9d8cec36d803e5d6ac024cf79906b82d2eef4d6b05ec6b7d0840374d537ac45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc65ae2e9d411f62f97e3fcb4ff1c20135143bf1d5af1870dc7a57d41bab6c17ce5e6c383e878d97e1ae9ecff4ac3c1b2ebd30bc9f4159c21ec93d33202600363ac7be2f7389f20e9224389b92a07589d0b087030cfd73c82d023f479986c5cd7ee5f333b99383ec18b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142b37ad77b0d7ef488d15c7c8af2eb8c8e7d90439b951a0dc0345f28d33635a67294338e3f2cba58e6ad703823187a61a7b528536de3ead72e2febfebfbf7acf4ce73dd7199a4e5adff4fd42cd03c678b22e90b55c5f06aed04aff4e5823ebfd265c7f5e929e723471;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16317a43722d7252b6d4e2319920984f0d9cd76f93bddc171a351b0c0b0302d0560ca1e17dc2c0709b13b30a4fa382b98d05488927a7ea7145b79ecafc2bcc8509a66aa21685f8b9352ced4ad1075b2bd48f932fbea3da558c7340016038b739984eed25e0b71f7c32c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6bb9780fea8d04d5fd304812a78ecc445f63fbaf76519203c6fb422cf5e53c2db23e1a5caf421a3a7c0bd34f454c800df5001021ec0dfeab0b29eb3f10157865151d856d3df832044c36467564350351cdeea2ed930830fc02bd9cf51a8be786ec57df67f0842e66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26574404d9fe9bb3e73dfcf7627c49d7b903b0392af749f28dfec8b30b4f9be46b9dddb84946f94566bfc4fe1673ab2cd5e6393b9c5319a574c4d5459271c36303f4b87e0138446fef6b6dc97f17c8587a7705d53277bce646e30d3a319666878848f4131e66803846;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac78ac2100e63a3f63fa70ac9122bb3868ca7ed387e8bcd5f268a5e2c6ea408b2f8d52c54010477c49c04d7478d7863c2029a2a9389daa1037e31512cd78f7d8f2fffa8b7cf60e4224c26a78772749ceae3224d8e4d59df2ddbe92faaf25976fd7adaa53a68d62318;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8c20e33b15bb1c1b28fe5c6f00ddcf755609c0172d33aa5b7facc2a040222c0a87ff1421ea3acb3742a934e7cec22b91b9778275f78983ee7f75ae293ec38208eded3d365cea8500d9966b67237e2442016f1fd8a07c8724a8486b560035c69623064d87236bee193;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h439391c5b2b152c1251b15b9542a6e900bd8d7b35ceef4c4d3585a75cf503471a9ac780bfbfdf859fbfe932e646a176e3b76b67a6dbd13982af42c029a1e2da9c67645e9827c2718a13b30f12284c4948a4a1e15cf4b754ad2a4c255f0fb256fe70f57131d1fd1c5b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17de16d92eab50a77199764eda27208bf0137626c91f55ea38b5e80dd46ee65b56294904fff30e56a5a47247186522c7f570521bbafbc1d11218e8e2290f1fe080fa26ccf44df8a67e041047c6bd340e1e18a43b650825976d1109860e7e41466c4883b9ecc9a2fafbf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f65f8a72f8d7ed45f578a2875a7304406524bf89830300517dba0d1b92b1a4fdd904da1e211254b95d6ff0ecdd964101f5e0f921a66a2902c0bec963b8ca0b09c734605ad6a15b0ca91c4f68725b2a28ab2f84f5d69fea0af803430e480d7ccc02aabf457aaf7799e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3823edca78462800a6d9171cceb0e045b5e513e5b0dd53405404b3dc93f77db3d7a6426fcaaf9e3a2f5112586fc09b87b192c8ab7b0b3232e38291ca063d432f80f48c261c461c6dbd50c2de7f9abdca52f43cf10ff71f4b0d8e2ff4fe7afe297e68ba79b80c4cf554;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1777876fb38a66f472421b10cceec21cca80512928f67dca3a80c87b6ea80e4b9722b1f77d2bb7009047ff5de12300091a7bfbd3d9f27d7c067d1a3a377aba968d6f243e6a2bc9679e0e1aaa72f010a692b18ed8c5c6d731d1d0b367695dd3d5fa99378f4579dea943c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b68fc18f53f6c2213afb3fe341f21506ef895cbdb9e3d721030e769ec3e3dd11030d19602c6d8b27260bff9d4c40bf7c2b390a76bf54166211f5281d957af0753f1749c4408252ce3be196bdd863a9485ab9495b13098000178dd08c825664eacb039bce444458f0fb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120bcf72038c4ca21ff2942d00b10d2b22249cd679a354fa116f8b28300293e5e8019ef46cb16f6d4a9e93fc8bae529989ba195450877aa84f28bed0da702cbc6f8183ec4839e0e7e161fbbce7e243fe571643d77da1912814cbe7bc884fb48584a6627c5beebac0e3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1436bb5615794ea3ae93d1300991a7d273027634cf64731f41055739cfdd8a3e61f5e599f3020fce91c796b299243c824e11ddc6c90bd0b1725b0ae6629ab225afcc2cae4e294809bfc1e4d022073c0320377aa0d3f7425d830f3492d93a3839f9d8799500972f9e949;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7826b6fdfad254ba3af74b4651b04126efcee8f946204862bde9b7f253590486a88188d3fde2fd5a2c5c722b86ce365dccd157df182337c4520814095d2d40045b8eb4201095fa79b461d2a9edce5aeaef6e0234a9676793a135cc494da902d044895dd6073b524f8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha913dcdf50c62ec8deca30e5cd6e06a8842924e547852e2693df59a83fee48c88892d84307ae714436879e41f49f98413b9a21f895cfd237ab2b0e682c0bd65638f0335a6b8b8b68e027dcfb9ccf94b16ed1e0a97e746b10262cbd75fa09e18ab2e3ca250ed7d123b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c276bef7581c7dc295ac55ada5f9093eb66355f8afee7391b16dc506bf4ec0eaf00869c952f7a18abda4f17ed4fdd69e0e4eae2d1a86830e7aaabe4a3116f848e4cf9e02b1fd9b0e124ef6ee5af14e4ad7a963add41ac25da5503450ddceb2b8e31a69e3af2ba3dc0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65b47985ec75923e6a27d7cc0cc340a9a6d6f10180f559384bafa00b3758ef05a44a41f5978ee2c272cd31799eee537186a79c2b3afcb10f137b1cce198703ef69d74eefccf7406c3dba15de403ed432407df38f76522bb4eec3369663ee59ffc85cc9a023b03919ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67ca671f4fcfebb2020101f43be6b951d47ba992bc166a7d90a587f2eb27e35e04fc1337002aaa04e9ee423911d134b2477ec41ff38397eae2da269f476a98bc42a8d5f1a8567515fab4070b76b6d780e0aab44117d1a8544bdc0bbb95c78b69789106782790ef0b75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8326da84ab1eb5db177c21227beccd0d5a173b859a7259270b480c09a4e61d8831729b510b99b0401a9b5984f0b9c7a23953050188596bd4ae49a2c904c30f41c6de0ce4cb4ad4f033e5b6b6848283c11b191b1e20cc8ae523a1a6ea82fc47b5996b42a2ddf6642ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c492bf23f4e1cbf4fbf792ca0c63a8559486cb069026f3949454e1943cf4bd19faea3537b8214d3b32afa59c37de78e09fb72811dbca8b05ecdec74e2fb11b8b82e786d011da1c23f8ca9080e12d7455e2e5294351786f3f9d92a7eef389d312d2982c40aa2653a7c0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167c0c604e749d4759fbab38ea53ca2e71636613da8b15551db735b77babab5ae38547af7dffbef581525c8aa6aae63f9e2e64cabe6bd8b5b57c0f4ef9adc5f7059ea0fe753909f1e2601b78488f260d713d67801b988e5c4f6964a021fed89181aaf41b97de85f7eeb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ab23ef7b43b452157677b15056d50797ffafa9e086126eab4b1bfc2d0acc9fcd1703a256ef481987eedeb05f20dbd5b2ce0dbda513a8bee7c28c998f1340fbe94622c15f8ca4bc812917c925496fd3b53ec415f37dc409b5b4713aaf9e1cb573552481c4810c7b26f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16204e6c569946e61a31f6ec161055ab1c5626004908d906a7feef521a1d9a014436165e495be9f68478da8058205fc8213a2bf9691521b5204761d79d8c427ec0f48507e2fac59ff8d6fcdac2cf7ddc3e9f980cff0b2f1fa6112436e6ca80516fc33ff185a3ea78954;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b5c53ecf4a4b0cead92bd6872f07eb55bee05c71a2c860f4b37c3af7b5ce095d2068294cfa04c08969b097ef0893fb915b7016981ac2723f64dc0a26537adc72eb014ef8be94e5c857f1aa3dcfb2d186fd58553eb081d2a19f966ab58f17891660ec3c44ca135af1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9bb23f71b2e093faad2ce99c31e577c2c8e28364c10741e0b3e743eae4086edc9557517d46922b72e62e48192a45dc48700670274b2f4bec7e13bfc45a6ec832b916f10d79aea4b6314b3e2fc711a2a0a41fe3dfe829b7bc6cd4e67bec9917fe6f3d1bb4d9d6153084;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174f774219d2fbbaf4d0c38f79c9a5993e8494db76e0da50103f1294dec6a10723098a6596a798a0c6bfa91bba10372a68441cf8fcace40e7f9543d89679ab112584beab2104b3bd554b55bf0891c3775a2aa7284e2ea51a4c4e595222aa005413871b51de6b74d95ac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63272c0603c8a407d57e526eeb049e5753ea422549943e7293730244033b9441f9c2d72a91bf105afcd5302c67b1af9b521cfcf96c47fd23b68eae30595984a6949c657cea4032017cabcd514b447170b3b6a4ef5b05aee4dad043197474b431ef2a8b82cff1e8100a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbf28bd697b6f6424cbfc53947f158aa9dbaf67c893fcab620a7a09f55da97ed497bf5cd0566d6123d7f37e4ea81f9a4583d7d9736e8cb8752c0f9c4b402f6cec8963bfa8eece8743bfe1ee41775fbf678a7dccd1f057b3bf28a40d9bbae1e7bde070ff577eee04fd3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5cf685581274ed52d6fcb9e3a8597ace7e816cc16849eb29d06df5b6e298fd6b9637dd1ff661c786dbf8a565311b5a7aa24eb20e712ae715bd24aff5f2a8d832e2b2740a53de596eb330241c4031832de4e47c298a059e3b9c398218caf30ea8d7827c46ea4bcca3a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7243f0119ef2e5948a7db637d3e508c8dda261a56acdcc4104cc23a4e68a9d0ed630798198ba85b6a690e7d83daa8f4dbb1b9c3821a873e87c95ed646e41289336d5ec4c8686f960e9630b5894928ed442fcdfd112f3410f4c710a3a39208c8f9809627040bde4c97a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0c96163b07c13b0ca99b09cf585e9fc15170b5ea98bcc632760a568454c8a4e689f6b676ec90a1b9032f3920bd393c1e3617636282dc7a289938d80d202ac0227854340d5c7869157b932cc0ffa99b5fdea1da6f02a3f0132092c7a2b5d5ca394d376efa991edb7e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b5b1c03d310b77b6ccf8c18d46e49c95def22a98ff521225b633a33673f1d1134e7291662343faad1d643c85be013a847abdf555b0bd7a341ae3a6a2fd0c7ebe6efe90776b1735e42293faea8f7d7e9bd7666afbf415dd6b72a5683b2fae4677cc8f8c9b056a0bea4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39328ee766f231c13dc9d56e25a1b8740acc659b92190825675510855a57e36f285c29ff36236181527f2fb886e1baf0ce316f83fdbdbdffa009796313c13ac3897280e835951fae811e4765eba9f4516e38e2f9372ab8b3bbbcbf13730332275c3fed900e0a3e582;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a225e32d2fbd5e3c7ba37a5c12c7cff064fb67f5c2f278c93dc070cdc790f35d4fa156dc4cff58ba2d6fca4dc16d8667e83cc98478c81f6715a11a5fd06d1417d0558bede9b531663acfa963939ddf84c956095bf6c96e50eafeea0fad2954ca04773020ff71717e27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35fe8540aa2c5473b75c2c1acf01217b1ef5f3ecd52462f0ad15ce04af0543957a1a719b6142cfbd567e14c8417015c893f8ff5ec2c6ef05fb2c8a5c9813908e9d091f043cf5e1775fd4fe61e0b57f365862f2270f576269cd4d8d0df2dbe01f08daac8519094232b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a508d22cb6700f1f2f281c12cb45508669bf466c8b39c0441a6cffe36e54c08b1aa0345443d0b72bf86e157d9fa11fc6fcff52ccc10726d90429bbedab2146dc41b9668901494e973e952b825e7a9f6c564bde396fded5977f6142f37da25b76bcac4279c72780d75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff932e0a66558f8c301762d44981c5839087b873b6be5e21e1101b48f0bd270601b96a7d8358b177cca5dac5d2b4d4ad39976e39d04a060f4c77ecb6529ffb48a1a5f6313444a1efd51936d0811552662ef44d106baf578f4fe355be7636b2c76e27addc75f3251856;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f0ad1a441d3ffbd6419af136f5ae63aed239a116428d40963ba9cb10e8223f551e096fd9eb50c619d9d3ce00d81f5e0c3b36c831fc5e056ddd76354c6dac206650d0e6c9cafa22dff7e8b04752a124adbde29d6a91561187d0927b3a5533142526d46e21fa1deeb9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5263a581a13cdd090aae0e74ecbdfacc4015991d7ab2fd72df4128f721ec6069d91933d9e094e859b9b2181a183c52e3feef82ff81f4e7a1834ce6bd459d20181516c757472ca9f9992248fa0b55a56e9399a8e32c33ca1d13c3a8ccb8874fe799139ad7d9abcceb8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h224e144b2af5e294c80f1515f4115024cfd12d753b2751f0adf8b79d83b37caa09cbd5649718686aac11a15d88d1fa96602ee40157e397806d719f84b57eca13728dbe00eb1f771d074f13839bbd029eccab5c50065bef6142d189c567af89e015607fedbaf9127e75;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d27830e71da3baea3d24d6689e3df94e4fcb5853972e9869063dc35ba3fa75ebc5bddb4d0e8fc720f2c4a4a1f2d377e5eb8bfd0f79a77fc1bf1160f08ab4e6f340c86bfc6ba6cc9b4a2b05cfa9f41cb630ff4acdcbec377472f39b6b84863c3c636366049959dd5a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc420147c6a9cf9b3a17a1bdf851391a06090ffd88cf1cb91defc2dff2e7d058db6f139f86ae4dec9c9932ffc4613bf69374ecaa2cad2bdf06881d7d51c0602c7d2e59415a9beb91a7a89efc52650c78cef1358fdc62cd7fa8f3542b6ade26bc6f7c802d50f009dcf1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a4d20b9ece05aebce6463c72e468eecb4b9b6a616c9bacac92e5abddcb8481ce4d7b95025c83aad15f0e9fea355bb7cc75cc37d54bfaf7cea51b55a23094286d982bda336dcf9442090d0b514bf7450291b2a2b05d9285c68e0abf84170b3f3dd2658ca150c187dac;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddf0c8b758fbcb52bbaac46378ce1f7f764f9d5695f4d6304c58aeb69ab3413168a27b4c3d37a3cbdd8f591269f48e5589764d5c53b99f2dbaafad26b890ab18769746a327db7ee4288cc318e76e541c8e04c4687a77feb2d2c251b7fe7a4f4529f099414dd5d48bff;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e604208d34d683f89dffdcefb1b896e07b29079049adfc2a5e137fff354d73f78504892ca013cfd51b68d6e4c62d253557b569ae1a5347694afad3be33ba4fbcdda357901f8392be009ecf803d996fa5aa29d1a030ad148cc60fc44e443dc4a81f97529088534893f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44b80fde192d36adb9d25310da5f7f38861fe7bc21f93ed1d43a3323a7e4c9c003bc32cddeb4d03975cc6ef2b9e45d78973d0e088d9495486a46ebd8f2dd33e5dce80337c11839b48d482417b2139fba1cff4f0dc0ecf59077e21f571d20e070c87c4618749af57ae3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8899e99c66972f57e70f81ed0cf5573ea266a2e925f3ae37ca7a8295c34ae2e8b42fbebaa68f9305fd1464ffcffd651561c0fbddba992fbb839815c2285f73336ccd65d9d8bc56aaf3d36b13439323eac9fd921df3afaf4b670112039347bb175fea24ac17e14b94d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d377886490bc92eb1869b80ef1d3d591311831400859d02e44a59a7d57ac879864cd966f5074304cfa6207215607578de13b41629a329feea76ab0fd2f7d0591c79aed47ff7645045313a713f8a007104fbf3fa3a673b757bf7926bf404457f2e3b5cb1fd0e756b136;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53f31c1ddce628fb0dd7367ce1489233eb4b56d39bddc11fa72854298486ce8a89f2458b4b238b4171f72192cb757f5d9e02c50452c6954d89a45ca883b1febc795ec51de916ad057f90da760de127180e10c3df24aff7eb7889d85bfcf5fcba6ce7d82c62c4d245b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc6b37af7f97e5249fde94c2cd9622deec0f52721cf354f29d0427974617db4e22f1658d562ded6d06adce478c3a05da386c63c8ebea86c8c4ace32ccc63bbc9cbd9d30aed7476ff83c4f2d975f9d42d482def77f903e4430ae949b09fb2a79270967af6c6241474eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc6fe6ebfa7187c69b6ea4c0c34960ee1c15572fba1b2d436c4b7242963a003b19202b65002d8a1f11320ad2840288dc65a3a41c957e86b6a751ea46801879ba9bf8e38ba8ef9a376f7774059cc0cf8bcc6441f36a422ef92a07acb9718ae7597a0e11cfe176c583ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha09c3c6bce250f4ce04b5705f6b83396a9dcbd4277b4a279bee35858f4f96bb9a6fd848d5ef5d23800a9f6bf7c213b8cf2a02e7f99fbfadba02d651628e5aaab9d903bc3aad727ef7ea9fe9ba9f4d984c09398bf3c9c7f2be37bb79009d8a9cfb09859c8336c889bf8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2524c38160fab9e88222013c107f9cce499331d12b8220b9ece7c90b5ce61521a500e602568974a10dc270b8f16033f9cf03e03bf7b52f41b61f74097c2ccf7586be675dae965930f7d23e4b4f498cfa0b867d9f6e41f00f49f08c713555c545f1a99170bb761847cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177e8bbdc6cdefd220a8b06c39edaf50fa182b03fcc9929a177d4035d61b5485081f428f46c75705ff45b083e739f7c9488fb7413134ed78409c6675e62b9ba62a82e12e2e04e1b74c45bf902f71216f8626b38b3f305f768c1375a954a7d7bd72a07662feadcbbec81;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18bedb95934d89124380c738a0ba368f3445826022da2841131024f1d3713df859ff145f9c04dc16e5ef89ce7af3f7164bd234d1957b6ef04c1513f322ead174399f2d47c925f049e9967d635c281ecb888a456d2f6b078347269f3c7073aa5386385f5ea76ea3210fa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5cb6f6b556639927e52271ae7d9f086785ba1514165551085640162a4cb3c75f7feaedcd4e06b6dc4832a72dd265200e4b9ec2cfd8e54d9d9aea387a13e094809797cd7c4ef90374088d6aefb3cdba8ae4d4f5a00705de77aeecde6848e68ab31bb9b5f111afc37462;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164333a736431912cb3e88f7e28c1af8e85b6f7fa7903d564de17e709b58c2a295a16a75b5f3e80311538e436fd1b7c98192124a3319838e136c96a900cac6c9ab0706ac33cb7802a83fc347cf4cf190f8f3939e690a41c4759623a08507b8210ab375bf03bf1b37ba8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac8e986e5f8d705cd276708cce45a6f918ddc05429c192a2a2a50716bf4320d6a43aa7ed624d92a3d32b5b8e537daeb642c708aac664ed19ed1f081f87b9d323040073a4eabaf430aba3d4a43b49612b428517fad0ee7b6e7fc9312acdc3010108133a7b81fd3f46d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1159d0bef6a01929db908c2b9ad22bc4cbd5faf581595bfbfd895c2b2b3784467885cee232378373613baf5e7cd1d33d0f5764da77c67d1fc18468f558e437391812680df56050728b6060a1aaadc10f26662f4f163e890f21781a460d237eac5db851d39b7d07f0b38;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116596158d547aa192c4f5598782fa5646678df9e3dd6dc6f48881a4915c4b4b88644b7c0951f5f5ee4c0c3b88f2be6813dbfff22835a6900c2d703c98ba8cf421b4db46e02a9a2cdff8cab73aae64ec3728c9ba0c9b2a4c79a0c37b4c78dcb0ba8a5468bd0fc73fd24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53f611f6f211794cef02f273041f45abcc78114b70b2a5e17438308913751d9e1480c155d293cc9d82461f8b176c2e7d70d00d6fada5469b1d0ca5031baeb12ec183bddd3d90575cc7dea981e67454ad1587eba948de83f6d1d84f22d0ba0008cff0081ff773115349;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h781f31163a96a0ff8b1328e072b68fb44d384283a17cfaa2d5a38a99992978b3d05f8399bbda8f885f1eee1da2cdff49a1703a080ce4b3daa9095beaec78948b8713c0526fae5922974e828ac5c728c872f517f6d5ff8bb5f02949a3c8088ad9d25036c86afe835159;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h242be2faafb69c809434da5794e0c9eb3144cede6e6c876977f1b9aa58319dc0f086bf468737f420d5531e6f093d41d949239fa93b4daebb586cba6c5c8e718318434c8abed9c633e8e516f2cfbc25eb560434e7e91862a0eb2fe1b2613b6c6f036c0eb178ffc98c10;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h245d6cde6b16b09ed1e9704d2b5a4f7d4bea315e60cc3faeb4b8317e060b6c49416f085c3c9e29ec96dea2264ca98e110cc9b8bd7880adeb8947c90bda74884cb590d42558c8c1838b48655a8cc2d5e8a98e5915deeb16e87aea323c7963f28cb2dbbe8d03224b6879;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb8c00e9afb2047c59d72767de1dc6da43681173997ba1a1230d7a9d491271299f58f1d172e8ddcc48c99d51e4968b71569de47075cc708fa46e4aeaf29c50451098afd438de23ec2c419514c32da8e96291bb4ef9e87a7150e19ca6ffdc70cc3ce97c09f48960f09bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h434c00aeef0cafb913b0197d1fdc77b37a13f3917a6fdc5ce0edceb3ab7c8e1a1c53c7fcd817db9e02fddc709eb2e1d1a932d334006b26c693e4d1ba3cb150812746bac92243675276cf5772f52f72785a1b76aefe52bc98ec4ed7bf712152c383ae60d3a406764454;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1548aa3415fc7af49d56208aad1c3a8856843b932199bab5296d17da6853c1fec33b1d84ae78f3cb36d5b3c388582a9c19432ef2e181895663ea4f4381888257c3971479c04384b63c8fb4b2bab469a460add09d59505f8a7afe551fc2b7e819f8c8a7fc8391f3fde13;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26ae5efce3f01a710d2475bf395c8b81dc5bd921c3d0dfecb0503bb078b322d3b38493fcc0a88d99aa8240c21c7458a24b4357c28ca6dd1154bcf3ebfcadf792d69da0f3f8095f21f1ae6bd680337ef63bbca79c5cf5f0045c1baa4498f3c1f961d162ca3e7df54107;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146f55e717109faf7cf4b67c9d95c6e525b0a8af11e7d3a9cdeeb718a414d23fb82cf2383ecec935b279cc58da6dfaf99043fe090bd52364ba285d03dc68328a3fb8e24b96a459a34951b1d9daa3f03a34534954e9e72591a1f1990d62fb147e27c6e70b18f9171015a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'habd18b5b0674bf5230abedc473fdd1f97c09e0ab7b0413b77102bd8eb3c296c7d32317a1f6e0acff83b896137019a8afa92b276f4f01a907bcb54e164590a89f2b90e8b2890f83de47b3c540d2743395b20a0d5641d3a4e861d3952e64917fa3a88be2b6f9c2c7e6ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a59fe492bc46251648665d35afc2235e8906c94046adef693cdc8c8f8a438226e6b511c0705c86779edebe6d4ca05b7973638b878f04f16bdd577f6050b5af73e40a7be3e624a113e53853cdaf7219f2ce39998cbe45b8428999bb8ca61482753f7968b13712813432;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9d4549250d0f1023a54332b280db2451dc76dc76e7f080b935a35f0613ef76f036bede9ecea1dbc27badc5f24c145787fcb6737e11646823ca9448a7b28eeb0f7126879086f9eaa658bec00cf5fdb81fb1c61fee46e81755bc7e84b2762fee32677ad4085d0f2c878;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h808c0c1232ce0259354f7d0c7ae3b77c67fe58385e51e8540c9ec2f4856ee5468de0bfe336ab69e7509ee86bb73a4f52547d165e91f9efdfdca0c08fddaae1aa5666392065abb0ad315695aaa7132cd1e8da3a9d00f9bf12c1fc2f264589b5914982c4a4701b0a0fbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e465e34ff6b244d6e0f407bd3a4c90f39e7c2940cd19da786c160f1b2db7d19f0d28a6357cde836e29c61b3a6d4be55ca749e14469bd0c0097cd0f706db8d915369592e3c495037ea35700885bacfb9c885005a8e4ab9c00895dc5b870673b81a901963f2ed41f0dd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190132a58fe496b4f79a5e24d0a33fa90c15e83f4542847bb855495264c81710712d4ffb33500a5a825feaffb0b7485f62a728b064a1720cb4eec1101ff80feea99bfe1368b51c653e5bea8711556d2c30da20caff0a789e7552748c66f9d69b8901868ff89cec4041d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7457508d9a85051d045b5a3f4e36d0373d9e4594872d9114c603d0e9d131ec8b72d7d57b18bf0823e82bd47abeadfbc788b33eac57ebb29f3da690ba6ce7f85da7385c6b7fece52ac0501bdbfb7d33e0ec4dea4bdeb827399631b07f1d138af03c6a6e2ab2c5f6b36;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3cc85b77deb51d0cfae8c9947006463d3b92dfb0d3c8a763b8262e5fe6209cc66bacb8b1696c333e2cf2f3d41190e9c57749964278b8ea0e5101a391d51a37d2e3ce7b6b675b34854b22e47c36ae4d55f38f1cae1b00285e8eee2330823967f45633fe62c6bf8153b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h800de0dd12f620627c745776fdc9b2ac451c919978bc4f8fedcd9325a8c57596504e951fef7ef5444b1d240f32eda48021e6ad5950d5b8754503906ca8d33b100ba539947f84f7d310f727cf8c71e77e5f745f113b8ab50208690565b3d0c990df0869050e59ce33a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79f27c8a78ea1270ecec01d251b263c7011c8fa1f213eeeb1d8a47916a5d855f5e56436d47559b08b488e00df961f7ae999ac2c9d264e0e1ddeed0d915a5106757ec9fc20b0124b91b9c6f3b5bc90a09ea6633e263873a6b0ab2cd924eae4f07af7092f06d6134cfab;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111e9d6113a300363e068e4edf3aeffe6020855bc17d5de2bc455f6a970111ffd3073fedf8e045d8f63f1d69ea77bcb4792ee3957539b990d754998f2bff837a7b90dcc2ef0ee9ed1b606f6a0db52114052347915a2ef4c9172cab0779d34ce453e862732c19f2201da;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb355c4fc379602ba8ab9e3ff5f10c8ca5c75354b5b3461390fecd6db0224464d3504c76fd6c1402ffaf3908b022e83b8b9b83485b7f8293dd7a59eb4c48a7a884f28989359307cd4f64656b24dbd07ada68d766a7f4c8dc495773678eaeace9f2ced7a9eb17f8a613;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaa23d292576e52fe30b19a2bf9525106c39ecc1f571c0f2421ae0a6b76317e48f4bb332bc56e56f14f337762e2f2270dcfd8e8a41884d34e13cd0315cc5ed55a560fb67a4b12ac9af99107fecc53f589d44227858d744f58bc2a61bba86da3d5dbe4fcce404a7459d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10dd19c808edf85eecea3f5311090fbf5ac9ff67ea9be21f09f78591f1db2a6ee7435de5d35a332024b05d74dbb70f381e38a2f56bc51fcc5f6139341d2758affd3a81e18ffab9a31ab0209029480abc0179b1c7c1b16b1c0a246cf57504c1bbda3e4458706e513db8f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heee655c1b83c2a8ccc139e08703de8637b4b6891fbf4439255a37f920e0fc20107d0beb6ba1d311ec1a55e4de254caf4184c7a84cca5962aa8fe50f97c68bcd433e11ef6f43bbb76eb174ecca77ece8419c6c07205bafd09df3c5f475376263c363555b34a76523bbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abc69c3fadea3239a59db5c0bce9adb3cba568b2cde4c79537b50b9d5ebb986ee14047857d5e6ee5230d29823d4da5ebca4c6f48bd8a500209f3142bbd000729ba947122f27c2335c4a896e2d12d9850bfb8921397ed60a913fb2a3b4adf3237b1065d8898dc3f6346;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a69a779867897f51a8c7d7449926c4ece5ae90a242bd59830da46adeda5d57c2820b396bc2c61ad0e3170d2f76fbd906ca8ed963f1bf2eefd0a659cb4ea96a8de1269659df46a85e2bb2aed474bd3609ee51e8f2b7c2d912ae30303a4f24dbc9b3abdb5d25896975d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff1095fe9c56b7c8d3966b57102d976f0f135fa60fd8f3a8b596f7ba89a7ad3d1ad2b59f5c0731546c661d840c3111c5619dba9dae629ae8690a8bf6b3f78322c1bd9f6ed23ad0bbab57d6993ee988f789e88be33455b7ab16327a69aac1f59e0f6a7b671d28089dc2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h660033866837df358883ec7fd5642c25520a66682ee917680fbec5d4255fb04de07b213fbeef492d995e756fc95fb7a1f53c221d66711714c4ca9721b7348997de8fb681dfa4ab0761f8f0c8ab3d1cc028f3acc8a7942a2efbfd2840bc4a1d3417c382bd7854afa084;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121f36d7143783d04ccabbfb15117df4a43d558f29795e324ad0ddf9269c1acb27fddf5cb610c2da3fbee2675023d0c4a40f9e9444ae5c88017e987f32fb0920e53f8fdba957271e8e4ae2b0b29cd64df3e0ad25a7048d4611c26bc84c08e455659ca72d5aee56af5d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7e1996f55e4a6bddc1199a5eaf20692ae1931d2b5df09dec2dc19b2f7a7670ef5aa6a642258ade2b73f07b7dfac5af6095c7e6ac84a4a44382f6aa26eedde6820cfd0730c05999ee54c068666c13d823de17bdd158c3758e488df822f9c005fcadd657647e2ebe919;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101367567c658ee8d16a6a4c1149f0a2b1dbcca34ee6ece8b96b8548b4975bf1d22a16b379310657c51a70fd357f04c35e35472083836d67ca700eb4aca9b8408d9a31f8f1d9b6842f6804c26427cbced64c88b4bbd45d3248390c139841e0a664c356d530515bb188c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187dd858a1c5ccaaec2af57fcd5a09638ae7f562f26b7de0ebef2f00f0fa0f10491c2239a0ee1db388a99965bf3b31557736bc5584dcd061f03b823cda6d307333ae27bce7c9063584b33b7d09be2d3e8f260869bc6dd3f8cdee5bc9eb25d71a2371567533740a85753;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19fd8086f1e3c4e255b4b6210a706c69f8719871295cd725ac51b6322afaf66715b8e69ca0b07e5a38a541861ffe6f00a0ad13edc5d4570be0517e851525a7681e96fe67fbc288d91d3df867c1c2d529809a07865051c62b86fd0d93ad9a94843b62f1628d054eeb25e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ed4039df18c41e5cdc4a8c385f692b4adda3f16c3854114d09fc041f47f6d0761c30fec4edaec1b8d4895ce8840d3d8b546644c933e2e486cb50897dfe8382aba4f52ca12d78e00b77da5cb570edf407e40aaaf0ba00ea9f3b353656551ce4b98bc982bccea5fef4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa907dc035816a7b169f60a27cdefce592b9d70ce593365fd922cc13187a4f3fe24ccbc9b8f5ea75f2dd185ebe018d1782126a7b64ebf6fc0c52e7cb1e594bb1b17009cbe84af70984cc12618349d6c043a2f4a4a0c16df52f9c3f50603dc193dce5cf1aebc1f25ab7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf557f3cace3b13d0e9e35a601475e62422ccbdd43fd68c5b8be6ba198886683f044b310ad4b589b9a10d3209d2bea362ba3e223532ee93d2bddd75946f52d3f360477720e78213ecd6e56d198a3ff10005cb6a216535f24caa192dfed93cf2aef0ddb0a870d52b8446;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75bd757bd795a39fc03344e583e7382b7c7b84bfd2fd13e227cb49a19abc103435da41438fff1986aceeda788758477b8ee5abbcb3be0e336a5cf71d84481f06de4b3d357491115c6f0e48b9880afaedca4d03bf731db28e01c41f0a908af850cf282bd464d0f34c6b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ae39c0857c0767ba38fac3b74147bf60df99431cffc10b64b2c95d4058e347cd74a2ce66d2a1edbff38ca35a72fdecde3eda48d7f1074bd870800f2f1dceb33cb0ae68456c4cecf20db393bbce1583ebae9f3c8840bb341780bbde207ca7e3345b87cdf1c26622f25;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c61adbdaa82f09e5ae7cf53b7416a33185c22fea7e536136b0b67e17334404982bf0ad845ff4999f19737cb654512673d34ef7f16a161d5ebd25e1b476a3bb2a5e16aef4f1fef9699056f8ac76ef1862a5f52b7e6672edf42a66a153c3f2189c66f0eb1d38154c6389;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56310414952298359754e4c4e6b7947426c8f2b5f65101afeb29427ae86944526ee5b0cda4db732b8f543775786e159463c7de6b0cee36b82c37937bc265ea1beb678984198664ec951f7992e85ab2e97755cb347ae6470f95ca91a1e92416391485b863c57b48cce2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21897b825d18a49a53c9b8b36fe25371c00119493489ba5dce991b156eb5cd9be48e7d8c594a8c3f575863453b190bb7e3caf9fe6d7a271ff42c55703109c44bb827c7f6b9f64e994cdaabb4dea814b446607ffb573bbeb18d181eb783288e82054d55949a98077b6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d90b6da70e77e25f2399b10e6731e996b59ba79cf2408ce3473e0fb74d417f3269be13b158fd548468a0194bb8480a28a0502b8082d72437adeddbdddf582ea9f0fa339278171acf732e5c3a29339e08ffadb075b61491e2765feea20b5beebdd3c24e43974696a41f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1affdd86019f56cc36fbaf15228dafc03f37bbe0a748ab738cdcfddf8d4def5e33f84dc5c8c3704ce4988c9b54d8254e69dd2ef5d3759b5402d37b315336967d26678e4a4a610a1a6d8620bd242c41fc56eb70622e6f0864cd6259236c4710e5ce35729dd783cdce982;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b70457c3247620145920029c8202005d1bcb9850e48b52a7bf1ad0de22b1ff8885244a85f057d7769a0d66416c941f3b3bec43549fa6a995f93d2d1c4d19b240ed85496f707370749e0e6f09f3b60c2e1f379630aba2128f9471a39041dd7d2ed879b78c533ce7146;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b4178fca8b4852d642bcf7ffb005221b88244fc08a39946e3b4e8443bda1fb17744838d706139237f71e7134a080c0425ce5c1fc489c3a7ffc3bfa90604a52893d89df856a50f42e25aa69bffba8a7e9571955975e332835bc6f6e5968c5115ea8dd704c59e34df8e9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ee10f72764bd0a2b87cba9c6c014b1c3b214050e0ba6cf7fb8d91d39ebd6545fcac501d535c4badc850f99d696900d58325f22f13d8f8b52920637588a5d584bcdd81173a0a68db3337d987f5ee2e6fd70131b222e048fa77e09f7abb72c602a44ad684e3c2f6585e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb96d9f263352439b0c71f8d8679882c99d147cb130d530f46d8eca89933cbd89f33dbdff3f12cf393be6446522647f8a365a22553ca4d7e30af072192385b6b97fb0474cf9f94e0fb3e6e1d1fefbfbf7d13cc19004e3075ba3f18704c445b4b4deee14d33ce03c77f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a7988f843cb90abf83394b3b574d893984b74960f05f2da3b94cc588c057a9ae295f69ccc64d2e51cbbd7c8ae1fa8fb379edbee0a6d8a4dfc272e3063bbc935c2c64ee9f54b48073aba1f24a435157e5fbe602449ebb37fbc516cfebfda692079b50757bf54eaa1c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e636705fc1e15803475dad5e605a9c13dcd7451ec5c8719a71bff96c1895dde4d08a2969b1bb4ea7a859e799d98e9e3fc5bc3a75059dd042586ebd3f1fdce978b459d41788cf9e77c1984bf89c71f150844ff1899c3745ed0ba8bfdc07efe006a04c6829cbbde67ba;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d2ea2cba01d9ea440cf2d4e4a3fddcd14204172a6362073c956123befa1cf94845e5b816de1b52b62391906d22ba97c0ded8acb89248e0a37deeedbac2467058405b498e3cfac7707990cc39dc540cc8115a332bd5b3693a2c98f06a2b1d5d9d77788f32b571882e1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd89f83081ebda4dd3819e0b2e0251be08a05da6d85d72ce1233cdccf6bac0f1bd496e179256b568b329b8690b32dbb6ad5331eadc11841c06030863fc751d4a16511f9b129c0dd951c559b730ac7e95430ee2267c622756b4864339aac82cf7f5003ef8ab832b72d00;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a139683ad880e6de88b2ccd9b9acd444b0a4033fe7812757ec1526e5f69a507294efd84f69679ec097a2387fe7b0415b699d120937572cf95d12e56aeb7e16023b47452a76f433f7b2afebb2b6194e1149b1d70e449c91447c2cf60530fa619a1b22a3d8feb66316cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122c4d7cc5450868f44d42c288d4e438a9ea6ae7c36790324169415a82e80688fb1ad6a1dccae165425e2085b54d71f631e807c50bc297fc27b46c6e63b283ade5bafa3f3bff88c54a43f24f727bfba280137506b859973539d050c67574d5e145c3a1b39c764f24d9c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5e1abbace17ee5331694661bb007394d912d64670aaa291be694245162a926a7639772a84fdc38604163b50f61fe754baeab8df0271632b31f620e4444eaf27db5830637f2f024b25dc53a61d7b3a94dd846a5c43ae8bf03e0a5dee35d31ab19f1995063928f02263;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5eb73f84d70becbb56b878cbea83e62ed3f78b41da112de69ba484b08e318b9f56c34ed264126994395377db3867a734ee5033646e7f9aafa9c40656ad61676754d029ae07ee88e85225860ce183b2477300ca38cbb217802a82bec904bf2b3a5dde22f096ba18dd4d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ffd0e4fd9d3bef6d4a1503b35c38237b6aec78f1591702d1984acaee343ff4a37e8753bf58d679d7fe35d71f5fc3298e751cf4411b00f20e45b33b3cc470fc7288beabbf5138919d8fb0bed9ab0f6c3b9d035a24e7cf670c5d7c1e6e9419a6f52a6971fe62efa3fd4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b4dc9cedd119bde61e720706319deb1e7099dbb921123263dafd45463820efe9012d11f92e9e56ccfa0d15bd6eb1c3642e64a7be006082d94b15151634ab4bd2b399def9fab7cf8d9333752ce580be3b3d7a63f1bf0617ab01f822ccb3e93a81cfa84d6100d561ae8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c6acf0a269a3db9fb3930b5bfe0e1122b8c725f501377ffadb56eabf46566ca3adaee13cdb3dfeb72ae50c7c6ec17408788ba5a7a06b1ab2dea79e64ab354a4eb0b63d3f9e76f9f749b8b5172aa8fac177efc49035eb17e1011a549833beef50cf0595b1f67d285fc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b00e13c5c68e9ec6a9b07af32608907d2b2d2a2fecd7e0ba06399f081be1490f99b413b7eab25fc2adaff240b087688598d58f79df1e7bbaf722e47860d4dc86288fdcc516d504e796e44b1c0a558a18b4054799a07a84e6a59d8df0ffc7b2ad3d28d4502e32405e84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c5670147d2d26d4fc762b73309c76aee5217d6f04ef9f2458a5cf0152470ed084b34cd84b247b7ee22337780424592925e756ca3564d10c56d2f511202835494337ff5d7dc0584c74d33a818ef986449a23b1c0094b083b85ea03d7ab19f891b6b307588b46749a72;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3aec5bb934ff30fed9dca36f74d18919214baa9bf28e065e7f2b3fc7fd7d13c66abb15ae98f30ba6831650a0d3ec4e0b9ab6a06723c0ccd97851a5090c9761d82775160eef4970107f896b63b202dfa221a9d72a962dc1b8d7cc2524b680930f1abb51644bb72dbfe;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he997e6c6bb77addbb14b0ee6b331520b1dacb2b078186206da066b76fc0e6024195a3fdf83430a9252f199832c1db8058531bf8baab0eec4eff4d788b58878301fc19daa885c3c0858d09c7c08b038fee6f807458e952d20cafd39f9584d111817032ca0e216754646;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127943ae7d98952600db20bca35811ab3a67012b8319ede260b4b92ad18887356328cf9b3eef8b631c4a465969ca8a5eecdd414839a26f2bb452df0aeb5d8ebfabf6aea4b434d64e33f11c06225ff5c37bb52ac5c827eb831c1f64e47939821b306acf10011e59d35e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ef8fd18251f015d71d38d6c3cc5186c7858f52696d741ebf18a3ee7174cd93735d62d8a46b28249b2849f88094135095c40e567dc0f2d65bf1fb9b97e75aab79716c352a133c593b10012a80d9a9982e1894b2bb0afba0395de6804cf52aaf0c6e6a1edb3597799f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22674b02f522c56de1b1e0759a16fb84abf43ae247df88747308c4a01242564d330fbc830de045d9cd69190078d147aa915fc8426d4ff2cc8be7ca1f5bc6428ab017c2a26c6cc4f46bd4f63ce5a78e544e7866164d665abf8b5a18a27370624ddaffcd2998553e61ca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ccefb914d718521f5303e524aefddfaddaf3ff6990e5cf8045b57ba1778589aca6fbe6532cc315ad000c064b309e7fa540414aaa84c865346172470fcd6c26a75af6686fb0989242ba5a84c03ff8fe9fb5ba3eefa38782b1f5bca9c298f62a05bfaf83a7375aca1a0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd977b7106a03b90fa4cb744bf6fd9737d0391b242c3d8b0afade4887a5c86f0ce09d5fca5369f9cef187ae6eebb67b72d8932aaa44e2abe9fc556aee71ed419042ce88dd6ac7dacfc43e4c886054d1e1de3e636416d339f7e7881195c123a794bd16adb6168f45184;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d98827f0ffb7fa154805997db59dddc46bc4097ee6c9a43e8997d6ea2a14d8a13191e9fe122ed4dd29cdfabc330567952acc308cf264ee3bcd377ca0f7254c2a4611189d7752531f7534e4c307d4f48b3ceefea4cbe393ea496dac621b4852007f977da7a17b9e7b1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1446af10c46f428f4e898162a3f8ecfd9517e79477d6feef80167b0fcc87b2e4c0cd51a614c56ba05590da28e1e3a2e4cf865cd93222bf91c653cd815c767aeea7c0c671bf83d9d997762aec48a8c394c9bf067c226eb8a2531cf8f836ebe53e09b84d276c79e368e45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188bb5fad32b6ffe51c6dfb88fc0b6a6640471747c0d27272d1f32c7e8d3b2a24cc544cb31a70f791e8646199ff0bc3f94a4e9021876decd69c3453277a6a54392a7479039b9bf5392b5a32c758b50350ffc4a9c3c72af190b8601b227bfb6f3321636a484ded487ac5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1194c067fa84723615b5d80e4692407d6a965322f7fced7a508e0b2b7f3b5ed3795a643b2c0e1dc93797e306f45749c7e985ed2b54f33005827c239003d544d3c9e52cb67c8e0dfdaf1389eeb80bea858ddd9338ddfcdcf3f9369bcc95de4b346ff6490b6a05eba72e6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8b597b79791e12515520f7ee5eba7ba9e484633751e858fa072b360405a4c5159a09b84e46fa20cffb3ce7612a19a5bcc79619a89a6cb318dafee2bc315ca70b75d8480172c1d5f96d50dfdcaa39e021bf618a771d5f900ad4cb09283d603c02ca367eda787feeebb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19783e49a91f339ea613ed94c39f86e4e9fc896b2aa47bb896eeeaf48bfd13d17adb627566148a58b79845b2e7a7f916b2529eb8eda0179d32a809dd5e7b4cbd59d3bc5afc7a2b76652bc1ba17b763374ed7d6b998b0a947657b4e45d7fdbf24b63e3ae2e738c2aae35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e52e861a685b64ff835e313d9303faebc285c3fe471e054e14c63d1646495220b76a933509c1b81f63b1639f1c33d8f3497e0b6b53cb900682c72b12f9004a6d01a4658e9a1996466e8e345d12d0e06abcc721fef6634a23066bf100950ffefe737c52651a96648b0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a9ab2ec5a3c9054c7b32f499d4bca25aa4dceefea0e028182eaafe2cb135c28a592d5d203601721606add67de411c01347364622dd6f15c1f9f27357dd3edb2f8456ac213a27b8e5605cb6b9e778431c3806370dfd53da229ed2b7d69181fac1ac6c354fa5a70462d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h650d6d846105bd766ade749a6404c8c336e588c4ce3a901d3ba6f2785cc91468465211545a0fbcd9612c0c600ad57549b5192d2d3724cc08e1878ca75099384e9f3f01a0c261f4efd5b48949cb5d457049c876b792007402f0e2cd8a8a20dd5ebbe902557841b90093;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78ac66675c8f1d0a1791e55ccaa15b9181a074f2e7ce138434d85017ac573488dd60f571eb6fdfee1b62de5b1ea30265e8b18d4b1bd3df1dd139d717b0666ddb6d06528fa61b7c4a4184949be9b2dc8aad69feaaf1dfac80cf841dce5c70fb165c42eae1b0853809a1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3e7100d168d9aff14d202aaf74682d718ce1992eb0a784d95e051a93f0a6173ab179e3d2ab4b75c47c1a42d31789f16aa10b2af08a2e6e442d36139cfab3ea64f630e67fcac516bf8c8535f7efd66f675b064c2fd0e81fbb1e1e50bd95828e1541b6f446b56f6a404;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3f24ab1a339eb6e12a8e09814023c6d69069c569c6af3eb14247da1e62c6b496e9faf939513dc903be3b653b1e2da296c9b6c049a1889245e75a073d95f3a7dad06eb6b79618675c4e1d4c728db08c79d168f0e90a5ae34d1b24e8ad31551b97b5646088963662cc3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e1d9794d3fb72c8480714ebbaf4f75b0e556659da5518db87eb85664d7d8837cdbc7dd75fdd9ea5befce11c43f0ea2c99a2adba7b411ff2fe4ea40a6a68fa05d72fb85b03bfabafcfa4dc6e642ef65c5b8bf21ec7dc6ae1aa555bfe92c8a83d822a5cde3f1200df14;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd5a9eafd47f7a111cba7ec92b9773dbc8ff58bade859a3d3d2ea81710dcbf78ca49276e471096bb864ea00cb0bf592723eb788965a81cab217b30244908ff8f92dcf42efa8ab73a01cffcbee13166d64a201a39cc5d904fe4d2d8037148e2c339f3cc7ba3ff07b211;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h922b50459832fa827f27f75ff2700a1826bb73880bd6a9712ec5f7940bdda2aacf10997df374186a5e1171cb9a75007f1a8f4a32daefcf794a16c4522cd597f58790ea08acc0a0d12e40543786e8d41df9a2e0e2d0016f09f67167d29abba0c73a880efecbbc412949;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb38a584c2b4e3a8759ad378abc8092e134af1ae8bbb303e31cf9f1d7e85e833492275030d2b3185581fffb4b6ebfca8c5da5b13a8cb22adcda071410e3fa667de1be6afa7c2ecedae40a57ef7cc04bd841ea28af0f9445b8de2d87f5bd43091c89db05d462a51cfec9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h68b1c4151271d8236f6bba1af0548cf126925f0f9fbb25da535690a21aece615c60599258667b85513a60e84503dbe3600c35b3d8564c5c8a18e4a1ff7f63a6ce7f3e36e6d558f27b17a0e255a5a7cedbf2fed4053965c50dc43180da918fa0fd0eb5ab51ce0fae157;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e779cc63edde21d5770bba6f2de3f9649e9f3a832c92542212014668620ed2fbb4e7027d9710478c9626ed3df97cb166068d716041df2f49e4057838c2db7dcfb01f31eba25dcfff4398582b493ffad0f4b71c9bb6ab17369440ba4b33eea7a02d309d50728fe4094d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c997806164c947bb548f53a98844fd41982f1469c4a582f63fbce128b41ec70faa2cb8f0c0596522ecc1477aadf9853cac65b86436e58b38002a01c4eab2396394c3892691fded7a62c7a80b0f75f58b6a23b9f0a1d711810efdd1ad6edc315bfa3d13d22b895dc0c9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h462b32833ab431a974952e706fed4065a4b72e007e02c08de4690d3cb33b68b6f5e53c7eb27261eced3c8e95d49234e4f12abadee2832173f976358f7d98e75d747e3ad63b8705d9412d1dc5824f45a456932947d2ca3d911f8e6c85ba88801b1c75fe7d98aabe0982;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e09e7131825ca687f31d36ca55586054012e3d1df30933966283070db2cc4bfb44f8fbecf4b2ffe2e28bbc593833f50b936286ff70767688ac76f1c9e7b62836ba76b926ede3d6a338f72ad2991d1c686c8c5c5b70b5694ce5337c0a2160a57b39bd9c63a711d1395d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19607615c40f9ac5ec197ae76a60687211b077046304b5a4a34d56a87c43659eb6be5089f2840e0a1c49ee8024f2d24d2f09a0bc8ab518cc81eb5636881f6adeaf9b5128ac290990d9c854f93b44b8ec5503ea18f9ec4091af572eb5924ffde8d588ae43a18f4e1cde2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f6e5c2a42fac6e275e56e61f55a718d692b9c74de4309347203cb04e2681b4a7570de2e40b3164f6c9bca1282aea98dab8d0031ac2a420171d3012f42a49b9664914cd3fea4b728230a38ba9d74f5f849425df8920405e289cfe0b60d063c24c68170735c73a86cca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e7d68e43ead743c8bf66f0a35cc69f313ebc951b123652046b692789bbcf15cf588919dabe5e56631c786830c6873002f65eacaa79a93c4b080ca736d5319c9a374fdfba5fbffaff393c29941771b65beaf25de17c09983cd0e3039522f7974d56475d23bd7cecc66;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134fb9b12203184159fcfa92be984e36cb18912c774f4c918c5f55b00bb8720f677fb9998b82f89c64a8cb75d68542ce8ab43fc8e71dee4690108bd948db9b4716c32b0d374e9f7383108ec2c426393f5c86711a989f5c465fa9ce7cbc3f7656c48d4290cf88d53cf7c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a8fd17eab422c6ccedb07ae76e2754a66c69462af15e7fc08ebe7977b4b471367bbdc2ce61e845c4913236454576fba3e291bf4e445bb6c21e026d7f3b3cea877a09a1d33b9076cfaac94c700f5d0275d642831acfbe43427ac6618c271c84ef04422f3ff7afe7be9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he979c82360ae9173e771a13f9fc1bdee4bb3e18af30e8ec21d72089b2b76520fbeb9565c187c4278278b82631729aaeb2fa3f8e2455f94d25540e6dce34ff180b4710ee24687a4f55c2ef6b9c7cacb06cdf858ede0e5e0c31cfdd5e63a932deae077f5747ed109b05c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d70be1940c8af44cb85b6d0b7cae3974dc2a9f0b987e406bf7fde55a9bd1f812c1fe0355bc6bd7ee63c8fed453e144062c7102d0c835b3bf86c174b825809efaf23b0869e551ec5bd01c6972990f1d775ba25a5b53ddc774aca30857805c454f1e1b8768780d81376;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c5472afcc4aab56aff92366af14dc779d19196feb6ac2833e084c9b6e3efa29878096665ebd5b9328b109b21864b31baa084415b5a65deaf2b0782b4ce8bb08e123a73d3446c7d913d1142cb6be02a87c23c942f4e1f38cb03e73032784e0797d33e9b8bed2e0da33;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eed8f6bf40ddfd3482b212ca5dc2299ce117cdb91bd4dfd690e0f0114b9e1c5970f1d1dda65c8bbbc402002f66792e25464a43241310c83060151408cb7e8233fb328b4dc224c5210986f18013a2f7a372f5fa566414e8ae66d21e114a7acac9045874174579d33755;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12065e45a76f6c5a69dfccb024ce9de80d8a4b7867283ff49585c9b79fd78796a3060a5b361c91b770e9b27145e4fedfa9e377479c0a94d93637d55d035c111ffb361ce1e8ecd0cb53c8b2921c596fb40349b599430d02abdccd8f439f10cad516666a4cbe5ad40b307;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb323f19ec3d56860afccb5f193b501014b9cb946167e8643a9eb0e16c4c01edb64b923d39cd86b3090e57a1c19ef9974c7e53103b3907085225670b37cea24fc8209fcef1eebfb7814eae1f30961ecd98ae45811b57fe5e40474cda222741e32ebf593634448b2372;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43417634fa63f8b07607b2ceae61eecfd76afb9ad5d93d81cdaf1046a33925875416710128fc14f1cbe01ba80e2d38b746a527b618e2bcfb115d7302c76c8f0a0effda31cb65bdc5b4049c40e34c2cf25b6cb642842ab0b9ac16103c153b19e7ae116b159461d9c5d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4f634033f5027e7650ca14d801178ba3ea7d516cba612b69f1f996cc5c73f47a5e4f9f5f22845800cc5fbd1518cecd15dbfa7bc01166c2931bd986eac5c5062880ed67e5e364c4b7d85cd6b88daea207c90d7df7f3cc6d053a12ebe3dd4afb944ec376af36eac12aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15cc7581488bb066987e9c5708466480ee4c91df624f5b8ef4f932eaad21dcd5a277bc7064003b266a11780e5bb6cadcf76898ff78a40e38e994964d44c2d19bbd6097d81153130b78506bf862fae58062722ab9c3607bfe0a571d158c57cc94b307cb55c8ddcdd9fef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7bd14ad11974445ed5d1bbe314e83b331283ce00d08423ff8a8fc329b9db54cbf5540ecd9f0a60ee98dabc2ccf018936e0e2276eb95f2951bbe157eab2c9bddda52bb3ba248b1b1bac2ceb608b9c1b9e7369f89f54b47f5b3dcae8546a9cb15e3479c47d04ab90def;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he575b078401a4cc331ed1be978115f86a69ebf062da0a7c9e15cba0f2d58c88012079208072358fa05130a89a6a576d4db4aeb52512de37a6983f073ae22232386b4eff2bd520e14387a692366122ede5c94596cb6962a128ad8c11a8dc6fa53e170b4d25b95c01eef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ac3b0c6d2cf47b306dd4cc2590b77d68af0cbeaaf58c45b2f62df25761c5aca02f17108a63e612604ae78be19b22961ae5ecc785d12988cfaac3a07a9c9dfd4c66b0048e216c1861c4bd0169dd60010c13e9641158fe6ab10536a321d6e67663f003838c7960d4573;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1faeaeeeaae08a292a4f884d255bdfeb62e59eff2656dfe84d83fe0881d32bb821fe7daa908b17bf23a792c0cc1f2b26999cbdd72c92c3092777228042e45ea55eef72942de1a35bec0d4f732a498b395712185188fc760f7a4776baa7590adc412c258acd3edb8b205;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167693fd7907d57dceba7a278d2edb6a0129a1e0c8a0c6ee038913007adcab61a81a1d397a6eb44562cd467abb6bf60b38b1a4cdaf8e9d5c4c012b0dbea024c2eeb417f1ee49203a68edad74c5e2f6bb33356a90c5d885b02c3434aa884d99b22fde2c9042afa0ad598;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13eb098e57562d3bbbbedb3f51559e66b72eb808d91d48fccceb366e3975b900a69dc40854781d98ee157cd98134f1f7d5fae85b6dcc53e4cac070b045311bb7ab93dc9ad771f8299337861fd89b31795b426abccf09223b34663ba7369e728409ed0fcd966e2fc801c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d41d57675f1239bbbee6f51dede44238725351aa928e1ec4bb6417495fd326e5c388c258afb5ea02dd70aabc5f87002e9747a1a253f3ee87e8c99f51e561471aea8ac3ba2b550372824ae85cb3a9c8bbef61462efc018fa752f1702e4c3303ccfc09f6dbb1b49eb941;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6c2f2912aeb38567da539cd2df01423e7a52e632c2cfb855109138002b61e2b22ec8d69c70817008d236bc3913d468baef5cbca97bcfa05bcc6542c2f1de52854f88aefc0c1b34370dd4353c535d4d58f5137c1d0424588b7d84d9ad4e7826af8ef4e74da3dc82a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a45021e8b7c251262760fb6f11baca303c54d3788a9403d65778e2a335001094ac8f7501eae0e8bfe3221e50452908474dc08f963802bc7cfe96d29bec916850f41a00e418bd0cc0ef901fa2cb249bcd7a400a26f1b2ac2ac1aae08f9503fb69290f7e14a1e20355b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f748ca644420f0037e7962336f2c6e18ceee264d940132febb1c5a50f59b23e95caea57f88d0fb4b83df51817b8656340cde6a218a3ad442c6df47c2e0ca6f6ade368752231f18bdbc0cd4f97e29e5c2ca731137cc3aeb0fbd22202a126a1463d747a83ddcd89bacd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1fc418fb26a330d5a4d43c105c2a65635e1c052d128a9abee5948c20fec80a5f321d7b6c3c727f92753ae7442d4a7bc80d2bb2c3b36c1aac4b70bff77686b52d3037c87d24a9fb353ad93f60a5ec9bafc81cbfc5ebb7ebd4c427be86382e20ffe0ebf16b69547bbcd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba92e23b3c079688b42c8e3ef91a923e0c7b9074fff4e780a55d38fb9b8083d14b9d5d6ec59b98187382f68066e275dd53df0c1072c7f2ab45a8b97ec88027218331bf87cb8b37b6e531c20b13a99868a9e32896d7256b7e4bb6f811acfa2db22125d15f9e5b48dfe2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee871fb1337cfd376612f058ee6cbcaf5bebd683430137edc4a8c94e8cebd29d28fbdfc6de67c5629c192c242152ccb136dbcf95c01a4fcc9c51e1957df2ab90660b5a7b94042756fa8a58b3e36e831e6d930e5949adeb4387d0631f51c1e61816bb208f6d8b6ab17e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbcf0083bc6800faa22c53b5fc1fe50f45fd0504a249a5c91bff0d91369639a811e13d87352117c10db85847bb85714276052c4558159b30a484b60e58fab4459628f6cf85e752ea6a8adaa8c5937878f30411eca7f3c68f1c71f81d0fc98445cee87b018ec39de3cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16db1d9f01b052b504699d53a823b83a10e329e18fa3b3f34df34d320cf9a2f92c3c27a179f1d6cccf01b4ed816c5ff1f67592fa91373f924299aaf4cff7ed58a0db2ef6317bdfc441792356b21cd7c28dc83b51eef23e48be68c1bcf67685fe0b9ef9bd833c2c7a82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27226c7dda1864139f851438fcbf58790af7e7b250154ebe6662960970d948c068204e9e9e121aa4dd35009631875b5ac0711c1263792c26c21f9066863793252a0e74828eb3888bff38731f97febfbea67f219743f15401a05f6447ca6b0f6b0b90f38e2688cece5e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15aa5d18b640981b8c563056520e449aa0ba33622e40063e1b6e04a5c97c2913c4bc54f09695a6f1ba0e04b3f3dd36f821ba94cc57348dc23e87f70888a45acb94f7a655010acca43cc8f4a24eae75c8da34360297a7c32c9b8e24002b5fa56491f503c7236f1556e82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9f84b860dfff84ebd0affd9250d12b538f7686c6ac3cb4ba525b2748c5ee73742ae8b9817ca2c0c66a39fc7aea0d1ab52c058205c712d7759cbb850b552c560aa45ef00c5a10e57b4a4a839fe87ec367ffeb07f833b7d5aa6bb694d8433f77cdad757fb4175fd98db;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ed6cf92dafd59a18772488f3d36155831a86f3fe9eef918f0b258b1b47db7e80fc05b673f7efcacdfcdf8f005bc85177a4ee59cc9df2c3fcea3aa3b7e22245f5f4411dabea164be7e40242c1547c513e23e063cb644033848908cb5ebb7e4d4c799ec5a0b2ef6ce2a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16dc6d73d96dabf2e8da29aba6fbc70b6f9723f93f3c0550176a879928103431090521887c2689d288e29bf2300460bf46f7e0450be5e145f51ee17a998c6825c4b752b943e555442f75c9f6b638031ff546f6a96dc5f4b80a4ba34147047195c804577a454e1c062bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb43afcffd0309ef35657830a8ad052fc06429d7b07d32059e0eb5e58bcf8d9b00f6f7bfffb17bc550cc53381d19e5c78512ff7163d134f1fc953787bd51c0566261fcd4938d782f08d02f8dce7653b2811c0b46d047aa5cb855315e3ca5e10f8d4b80e695729c3a1d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec3b3e3bcdb03aeca54b4b27727285bba5a3cd332f9c5dd0190c871b33eedbd302c0bc21aff3f079084051a13fe813147c94d8cde8ecef2de0b3e2c849159ac8119c615a7addde2dcd7b829706c6d18446dcfd4bc904d695fbc98556d8afeb305ad5001e574a446378;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda2e33d6d384684277a43ae9212379b85a86ce45e6f4477b5a3dba605bf072d216c3da88f7888d3947735ec47b51ec229011bb1056bf976021d3d9512465a84d8bd75a1880a0ced856f34ea8f2a419fdac1fa69f2083f1c6d1cdab661ee7e9b52d28f9e7d5367b8909;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1285b56389ea76bd9a77733c8eef342f9ff432ff9f56216cfd9f8815ed37872b6310b644b4eb5d4324c29667e9c5742f68f8324d7c02171b07515432f2ce62e33d1ad526495adc0e6b8a8c992b2e6489f079da47efbccfb3cdc094d7a3e62d681cec2b96d0a2425b606;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'head689d193df847b96f4fe082abb7049e305a509d151885138c1c781c4a87ccbf426a233af19486cb804667412855eeb6c68f407193363c48cdd79d00fc3e095eb091f484e9a6d22e041b10150a2c6af0d68ee6f6621a5e75cf0429807face4e2c6fbd02b5196caabb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaf31ee7d368b0ab4851ccf5762aa69fe77d760c9bbd732d9226286980a0baa3a6aff6b49f75ef3978bcb4f99d61ed1e28b80d07308af1d6e5cff44a2a5de04bbd72c831ae29e14e84c5bcdbe6ada13148ca8132bd0320ea6c06478805e4a872e59031c0506fb196f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1609ad7858bd13a3e1867eed9ab1b568694a94e2318c815bd878eff4c95012025cd91afc139b3dc4c3501eb3d0c568089995a71f27ae3cb70fe82358053356669d87e7837d0174ab0f41e0623ed2c00efbe4d3b045b33ede6589a18ef19d18046eba0abdbf7ac25cb9e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38b865febfc63c6b4a737089a12abbb985f225d098a8e62f0652a949ffc8b7b5b963bc542d358bbf9034673d6b31d9ec7d1f9455fc92d3f14b0c2d1b00ccb57c78248d4ea99c7cd601966744ae25722acb14628056338411ef353fa86faf3aac26e07bca58fcbb6eaa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7d532759f140b0e5695f699d08dcf016f9b0b3d32e74138a5c5899a82cf3fcb9fc38005db35a2aad009eacb657bf93bb670ec8cf518aa21a408dcaf049299e2d39f1ddc93e454339273c73830b91faf1530fc625f113b3b51642c86b3e4fe5674ad5e2cde6aa2fc03;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cc68db300bb471ee0ff51ff1c83cf314dc805dec8a88d8925871ff2ec730a9f3954814483398d0a0fa48e90d005ffe26ee523e17381c248d4c5b11588e932f92f994841165e2ee6707d9993f9742445f8c68814bf21bd283c781fb6be26a9df28e3d4cfccd9ce6377;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2718b32363cfaeeb7219267b1cc2e3acb23f6347f67b0355b664c8a2bbec9aaec4656c9a192bbedf4581e46aca53e6a53700d53b52d0d3697c2192ba3e3dc3078faf4eb5e414e0d39a54ec2e341c0ff044b631cd334614aa8e6d4ecded8a93340609ba58de02d7d0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h435d2c5791efa1f3aafc1b33b10f12d43e23f18c886ca020c432684983767e5d23a69bd4b21cc7da41c17122b2964c0638450c1a849ec77b2ea8227983d5f803b1f82694c48085140137269fb7c76cc182468728c7ceae14fe0ea2e439266cb22941b45eadea542393;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17aa1da7a4b8222856fa117582ce9e1a57fec4f9eaba96c3fb1a5470b0c543e4983c2e6f1773324a8e9fa6025ffcbf2bad2920b568ac221e8d5897c2de78e0127f3922f98021a346ab07bff589276c19166fcdda959478b157f67b8028e1ab002d2f8ee5cb8fac4f434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd5225e6c3e8e95814429a18ad4a2489071bf855e5ec5588befe4fb91b0a3acc776cc1acacd5b8bcb125e83bf849ce1ca7b5d025e8a60bba762130945bac6fdb699752a1dd59899b09847072b506b4c39b9b75a99891721142bfd330d1e57fe727b2fa501a2ec50c543;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a940abd6d80f46ddf1a60b9c3d9f2d0d4b3c725f054fda7af2ef1ca2b8cea2bc3dc84b77cf61a149b82520d40bf6f1d9747b562cd4617132c68ff46e73903e052d8973a8447f6d6d3cae1bffa8bac1b26a2e1067ced821ef82249e5b9dbedc0a7cc200efe38d1805a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f58ee23279754857eb018c45605d715cf6d120aaebcb35599af1d77007b844fd742d7ce3fb4898694e4509a5b7be13cdd91d537a8752f6f8ff32a4bf9c8aae725b92d4a139667720547c3c0fc2d12c7a83f0753d886a7a1c9466d17f9432c8081f961cc2a44ebee324;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e747a2bf46aad8ad8ec7c223efb070d4c5f387ea96e4cbaa6b868f43a316d873ab6411ff229b883038849c88ad35733071c1b753e0dd3c0ecd3e38d000c3fc253bdf7a6dc81c7270e51583d6e9ec2355cee6373724516abd69678f9a887d8f9a06509e7c484890790;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f6c0572306b84150cac0a63eda3ede4a7aa325b4664155dd3e110866925dd8b57adf385a6f370d15aaa3d6867d1706a22afb2597124838460728cae8275c8e6df0824a72d1b4e382b5c7abdbc439267d5b6d69ad7980adbb07c59a74067186d48984877255a71ee99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h583ca02ca678077606535d6e1d3fb7e3d2f547e3c67e5036f1a8e7fa26afc61472a86d81c74f4b8aff9fdafa3722152bc2c860ad6fbdeb2daef9bae38e3c8c5fbaf105f8a567d8eb4ef163cce3ecd3df85e0a63d15e3e8232dbbd66155b24a61c35861449871d2b249;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127449a0fee6b64353ec062d2ffb38e4836a0a3bf344f6c140a4747a1534f453a7f8551faefe0a2aecfb04bfb414ded8a2f0d2f4e8831de9789c3dbff8751423fa8c329c6c872bd592527e11d7b11d83b1ff4f97049e8abc08bc26a1632c00f9a88ff8e796ec3b5e433;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed7a72d471c8c02cd753485cb2f73793e49a5f928e542ba67be9b7bbe9db197f82f82436da3b3b77e1a94f910d944ffd0b3fbdae7076f8a957e0ad63e1b2983b9ac3602a2fd092f40b7b1360449cd5910e46e47b5ca88d78f1c21fd05b250b2facd75dc962b3d4005f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fbaf55508739e5893e173952a55b7edc20838667420445f0345b177802667679aa0d88d08770a0540c4e141bf03776238de04a57d7c9087f064652942903cdf9f9c8cb1b0c7d39aa9ca59ec569bf04d4bd1d07a4e3e10a8dbc367bdc58d53ec307af8ed3545c6005e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ea44b9285aa4757ac7a5e13d31ecbc8f1e0029f4cc601810e059d176ac7ab79378007d1512af71688e8b5fed88369b925511495658dbcd7a3b0f35c07bd4dfd3ad6a9961793cc92e70fef229308a04465430e2c9b9c0b9e6a2b6bcc7f99ed5ca0dfe641630181e53c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1699db709c4f73022f4acb535a668ed9e11b5e8402b5c5c3caaca8f6e279345f7872320d2316f00e89ce64b8a945038990d6c9405a02ee54345875986b238be7376dc77add08b5373c258bd2ae7d9907f230247d931c2bd21747e7bff3f8902882208276423bd457fed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4af015fbea89d44f7ba67a44e8dd6e799d1aa054ddc499599b29cf5392430c9012cfc1369c316d1ad0aab7ff4ed9268bae0d373405a83d29531ef90924cc4ae6c8df7d1d1358f8290fbfd9792c29ef2b15d11db71eb5fa242c8360701dda6be24ba1885ab9c523d91c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h199b6c2c128d3c528131a59d4d03eb6d9e397f0578c9b86e20aee0342b2bc4c981d96dc407d93528677cc7e9342ab00a4b5ea273ee19d37f8f8fb392740cb9938e8d13d15aea4e772a6e4c6338b6cab5367c6431625061caeb61c85f5e4aada06694f89e401b292f135;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179f2bd1d8d68e68dbdc61d906e8548cfaea53f978b0a7f773035d8dc2620472d5e5b330a045a576e560c1a4f4a0d7ff81e3363686982bf94aed966d3f106677e5e960ce328a561a9bae01008caa9a704f30170181c820797de49e49002e7c596dee52b06de4128a1bb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc571a0575de711cea2fca0792b62df4362c3390c34d1a7c43911d46c0740547943a71745ac5175cfdb2c99cc55757da85daccebcbd622115155a39a979600dd5d2e4c877d5287d746ef5bec9806537af0f1e74f31abeb086059df8b684d88aaebe057677ad2e6c60e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2804c88c7eb68d5aaa952a07dbbf2d5e933e2c11305beab95ad3c7bceecc742ccb6add2d3f0b7b14b1327a391570a058ca5335f9a52c9161e4fd02ff1a982196f725ed76f867f4643af833e6981375cb8e42813c90e4a7e97b97e7d26d75d9d651a0e5338d8b32b31;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9936b34edbbe2b3fb3ced2405452a9c9cfde560791b9353bc684ccc921bc19f6166c984cbc092fb5d07d038447fee9d44a0cff2c08e5ed9f1f95df921dc3ff038487bdacdf873ea059a411626c616be8b1abb9967f7071d1b419b6f276717ae9e32829ac98d00447f0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3969d98c9ed1ebf2a1e512d209d1368260b2d9e07f5aaae940966757b815afbc0dcaf3412244d48686a35c999fd4f31d8e888e2862226fc758cdc524a7ed5dea22929e1a10141749d6ecae4a4ff494d729d348002848b31e995908830f508f0529c580c0027129a35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hddbcf8d0c2a5b5d60b965e0bc88018a406055c4d5dc43245a0b1262e7bf4954178f9a2ea980bcf3872de36ad229cf72b4983239781b24569d28a90234514e5089fafba6feef217a2f64e4517af1f7dc3c87ab3a577dff43d9846622df124c8b63734b7425ba4fc655d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha30f24a0247157a33b2cc355ba2bca57e152f1a6b42b05936baedfdef28b9962b75fd807cccfb41e8763df489a5bac20faf09285fbf9592dcec83c8dc51c68a458273f3ad6e32d8ff9585b4f231b986ca12e3ac5d07ec41e5499965213ea9a3158568e265f83b9e1a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h949f28556086bedbfd23dea2a0e1ae3575be7b2f829c0a83f226796b6443cb950f309ae82b6d36f1af3d110eb6d6784db73d54f86d96d7c66fef0232f6ffc3a17a5dba69846c8f3e1a69b9b5b5c418ffa30dba86fe4b2d67a80ca6f07f73473338ef727dee47e1cc35;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8b3bc009111128dc6c55acdb63fee434f165742119e5ecc845a94b4994cd5d3eba277dc476db9d9a16dd1f37e3f95cbe1ce69464da24f3bb6b26c213daa324404e531b6bf0a6fde305e8b37f0139095f9772e962370f90c8566ac8836d80a870b1aa93c0cbbe07c24;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d3fb76f2695682ab332a58470de363aa71c916b60a6dbe60e56a85e6aca6e553227f595dcc32cf121fff15363fee9b2cb171c5c970a39bdd44d062f39035df6b906fda3429fe7b09201e4a1cdbd18277565fe571aa8ac3e63978f992ebaf53617cb32e1fa131df597;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb595a3e5d05a699a722be40e46a52c87a369c3e5008b3356d2db92afd300a709433236ddb787492e5df659462a7a7097d315cb65c782a467aed31387f0e317f3fbf53715e5dedc06dd644991404918dbc65ed1624e6bd858977dbea29cbec4c45955fa8432e624c99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd5e8ce577fff45d1ea073525b97c5648696f25570a59ea26097b80dfcf620a3cabb67fd7c50797a8ef8d51f2ed56794ec32f35894838b16a2aeff0ef4b155bb6025058c089297007f4d3a577710762e8eebbc7f5245d3123a2682d98a976429ec78ed580219ec474d6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b54289c100f14d0ceef0d0c6aff579f2eef90b7aa970aca498d8d7318b10936072e8e87be9ba8d1f066858c4d2b38042482d1bc8ab6ed3619208422fa06e5c9a4d65721407697f08aeeab28cc0d8d8d24d6a7db03c8591e5d1d600277615cae1b460b8940906869d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106d7e364ad21f047a83ca79898deece1889e8665c234f57839118b5cc476a13f2949c016745664494a8eb13a445bc096433ab2c0552b1fe90d1db7f80396cd42967f5a15ce7e27c29123ff73c55aa61c9c7087866db84ddb4c7b49bd1e6432ffc1fd09ad09bc7238ee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be11fa1d14128a36c11dcf09682bf266412bd1c7a8016852ea9945329bc84f0628013b6360184dc1a107c909e458f778d998360a44d8e41885dc90ad9bd87d757362d9d4b64ae8d16ea128a7230029634b4ad8ea9c516e0b5177882211887fbfb43aae155a90745c6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11348e5ead6bd1bbb95474cea4ff14216045b0e24825da441909db85e8cd5223e651ed79511083eddad58817b4ba8b787f3c9d362dcae05f55f48deda93724fa0fe5efb0658c67ccbe6aa73b58259220b6c826429561f003475198a78d7d1e371c2714f1b24068f226c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a949b21ca2dec4ff82e446490374bf4e18b309218347320f33a554e5eedddab87837dc5cc62cffed54417110032b43b5411021d695d015ba55464972dafe6943197e0cec424947b62cc9d3da0a63aff08b9fc53c4e8f4b7262a4b836656ace5a0c574639cb4a3af993;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0630b9d144cfc469a8adbb31742c3b14b56bb276b1c4aa3d7c778dfdf50bea229bf2196728a5ad76bf34a646ce2acc503bba81f52804185a547961f60705a2af3690720e76d468e19676be00a2f0679f3c444e2b3d503a8ebe34780327568f49b929522020d815b60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1250f1271cf35631b6b27a51f39c1971367d33718f2e1cfb378fd6caa66a5a936a94963c038865ce2167e5d66eb4c647197f0d4f9ffb55bbb399ed312bff292edd330c20a67f5a690f1cd9983f19d4ef3ba2c29320f36f3bf2eef8be0ce85184007db51cd8e4947ee27;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a3426d1f88904eaefb9d2ab22ff3ea06c2e5936b8f221a8aedb956e14796e264411dd2d36dc997ac50584a3768d6b12b270c68bd2e2de9b8b00614728ab6f9de4ec135a2a7fc186372aa391b6d1071244fd53520e41b9ed9a9fc4e1c6f70de698da1174d4eba05d40;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc22495b64a1bb17eda897a5c678163ffd457dd9a3278b079106b8662aff9d7b500810075426fd093756c29284c80e2cc0e3fa77e7d2c9ebb9e25dbeaa2987053cd6890d6ce9462a3484863f927d1c4d1047290fe3cacffa4222864c885511a73ac8242dc4896bbb9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddbf2f42908340393f2e5ad4d877cbdb2c56f6546ff1020eb9304f0dc79a146b7eec7bf03e5bc569860e68a61fefc506b99c6a15bd72b156030d9fb1f70d6f0970be3e6c8975987f5f449e6f8e9f03c5270c06b24912e549a42fc2646e0bbe5c47e8a03f175ca70171;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4ea3a25bb74879322ed4d79f33e36eea0450b06a85ee9e4bc481b5c0a726ee2c70097286354d20624a2d9daaebf611badc5d2f70db2c96bd7700cb4f0d358e44a2845296d8b78011a6b8ddb57e2afac3f1e4630e0b7f6b8a7202a9bfe47faac22a69a3c17e1e48a8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h658a707639375c44a9813b204925b9fa690f5d6f2a9e13cfda3a03bbc3b25446a81a2472e07b1aa9474b03a3371035bba872d7f3da7e2f3a0fab29f40499e9df6091e4e7b5b0c21e8ab7b5bdc50ade8ceacad51347b872bd09074d5a6062422bab320df03180c9a20a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13bc4c5d34db13ea258a7ea08281ba1a3944f7ae555398cd32f2d39f1c71803a213e0c3788ab0b57e82d6b60bc6dc57c13a0ebe0c1064d34f6333b12127e02ea05d7680af48183933340b842d27ce45074e9b5175214be15442f9433a6c2a943afd03b84e01d90de0e7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha02aaa15dc910d5ad13786b20561f0c59a0908ff6378ec7c014159a7fa950b10434db750421340c83a71f9820dd0ebbacfbdc91e2fff47e15e5557e235b5777fb29bb7490890e0e669bf36a32a7bdb5a3f2119e28b953707a2a7e2730069d4a14ef5e5c88d287c92b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2383da12bb9b9db1c75b96199752bc1cc0825c10d0c5b2f1ab488aabf28986cb9cb1ccbbd9ecd0d8e0dcf55f210a4f3304edf79e42246b83a549f061bc4f18baa61a60a4730c7714c461e89ef60255ae025fc87fe890034855cbd379dc8f50101a29aca9f3c113bb3b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3849fbe2b1f7440f5ca4319f8aad79aef260d1566eb634025dbf62adb3224b716a41013cd2eb8228c7e3acf5a2f187891081cde6c038ab392a9923c163b667c5a6ac960ebf461db333db7627e9c40a507e866459e5ce69b194fd845c9a5322c6f00e253085259c7f7f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb31649300908d59ae7af6023ab8be4b10f7e75eff16113ec786caefbdd869560be897f223dd9592bfb8d1b77322300fad1869a9f5bec27ef9e00cffe7721b76db992bca17f139ad1773c203f9f6355867e8ae37b0a48ef27f9bb471dc1f4c06de24208af59aaecb07b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a555d433287d2df8908b1d14868c003085a1d85004dead6b14e2865e8a5227295f53b06fc72f2a6c6317773461ffe5a2d5ce910ec104b46211adfad2f8d15c04aca2cc401af7d9ca581c0a2cf4d3736b8ff05574e03ec0b2bbc7e739eebd4d467880d29074e14ca84;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6608592bcecbcd1ac90367de3ef2ce4d82fcaee340a0e9ae0c5332a0d0f7ba34aa7b18ab58e45758c1ef304c0f97dfac43128940c4052339fb4c3ad3df68fb8b45b38c889d3c281ac06a054f79a2b1ff734b1ab0efe159ae00516821017f85696766eba5b8338a1a8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc933d408157cde9b8df9f357a7fc3fa5bd9191d2ffbd6c69dadb98ceaabc75e8a15887f63459c6fa98a74ef5d5d6116a306a7e12c29bf7e8cad6314f49e89a0bad40677d69d5a6c5d20e4b68cc124bef33869378a754a5bc89f721ae33e4e43db5725e5fe5b52f868;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147f55722de223b67773c193896434463bd8e12a8799f944965acbb168becd49ab6d65d599b3369df8f0fba6fbaaa3619436869f752f4fa84a0ddbf5cbc0d8e84d03b53e11271352c10e091ca940511f4e2bdbd6ef70ba15786855c31aa6bda10b05f4a36561f1f8631;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dbf734eeb6c1f7dcd13680eed70951205f41b73ebb69512cb5bba4adde4cce2a4fea52c6892091bc5b2a6ffe12db2cea88ff9d847390fde1cb728da8546925755d520691afd83edd4067a00c3857925431688cf32818c777b60f7b87f5383066bc1464a1c1b65bca3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47e5fd13844af570e46eaa74f31c65330df28fb8a92aea29e43e35646ad0bd2739566dda6f6db0f0e2321a9e67c7d684b46794dbb2981b18f3b83a002435ad7f23296c513dbf3ad356591ed1e8a9e7957495cb34f02f011b5f29652788c6c52be0657c7d1803538a43;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a88f4b1aa06af211ac540dccbb80f78160dc8e31d3817f3ce41d8e90a9f6923f92eaee215b4f45435203eb51c8d495b6a365a5fc9c0f27f3d3418a33c63b5d4f63b5f6697fae6233079d5774ff821e61a605a4fba0172f58bc737be1cf4662c0779159d5ef450b14b8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h189d5e838934a492935e06dd5ec369a63493c1c7d5ee1b078dea2bab56391a3c1ea16bb36c3fd5db06bb1e2bccc00e86919481e304072b845b6b3d1cd01a87a3ccc405f9604da9d225f7f3c15f66b21e9e44e88bfcd7da3e05406231c1a8d10c8130cae47af68377649;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132a450150538b100e47ff1073505a8420a79ac1f6c53e425b10525ad3b796c41358928b5025c66a1e1004c4ff0dc00c023521293251fd52efc19e3951870ec7ea6172f3c6ff04a60dbefdf56386d1dde03660cb6dd4d68d293b85b34bd29ed411cd90b203dda5610bd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc6c46ec1d358fa59cdbbe6dcb62eb0ff87e3b21125b4c9fc60de7ccdb1c5a4f3c155ac14c8b2a9bd8f3303a858942f9cadbb539e5f3db7542b1f03960c64f5a7b7a07f46eacb2ee52aebca88f74e105e601576546601f4e042b7db3e1396a05190372755039328718;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2be22deb7599a4d9ba5bd3af8dca6fdd07538dd62fa77e0a01c9a29fba3704d1fc4c4844855f66403f0e03562ca8708612f5e1e25ebf639285ac81f3ccb7f3e7a7af241ad332a5d3c9907de0ab0630298cf356f6a5031049b2eb6779923821dcd1f9da81620dbaeee;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c99d7d9de03cf7fff32944f5b34bac97b3817a1c627eda6c7720336418442de9c082cc5bbc4bba78e09feeee5c7f622f7431e544ad222eeeb4d1735b5b4ea4a9efca22a6237e1bf1b91248002fbdcde4b23be4aa4e2d8c6ae22e909936e14f7d1adb2e19f42c8a1be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h367723eb26268b5257ae557dc9badcf93cd6484920f40da28aa188859b823dc189f1285c6ab0a03fb17a0462dd72510b75bf634ecae68c211197eb3b605d5314855a8efa068c6dd063e4c62600f756854be61ed68f8752386feb9b3997db907b8059da98ab30c6e789;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbb63e6b263bb3877d8886c8949af5a4a0a83b4529db43a576656bbf6b34b3f28f61d5fdbdef60e406108ec1cf32fecaad04f6a47624e5412bfe1ff0c76dfe0b120d0cc1eb668ea2a2732def41f8cad3f0c54d20ff27a3d7a5f1a5ec866d2554d071063e32fbe9a096;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c5a4267d8e746e5b0e38d16251085d98244c76954abc4efc35082f1ff8b97063974608bb7a345e616f2a28e876e137f0441f97119b17c558853ede6628d2834a1139514877ea1e39a6865e2fe371d8949e6a4433183b47cb64b6f5172b658603d952b37f876eeae69;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1511559d38a18f01cae6d7de2ea665609ee3064197d5b4233c4c249eff54a9912511c638943fc4e11a062b408f4e8a965d297bb30972c6b3ff8c0c797db2d4a32eae413823b90d5eac9da4fd75a6cf13bf3cf89eb31c3361bc3f4320513c453db1ebbaaacb84b18be;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123752376609ddb68e2ab9ceb50164af7e2b7036599feb678a56fd92fd1812be2d7fb03281a0ed1e987661eb9efa59c1d80e30c5705070e3141eafb3d66d1e6132ddf62921feb87fb93f79f45e052fff37e332923cd86df967f1db7bad4a84c79bdf935c3244ab8e8eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9af7f44686aae04108eda2300113d7930067cf0dab5d2872f3d592e055e20618df8001977d94059333f5197a959e0ee006852ee7fffb0e21f902cdc30d1c9c6982ccc7619dc057e004b869254404779e8a992f55b01372da5d140d81271a74d709945cdb8aa8d01c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149a3a1a40a123a1df1fe2f135c3416308d579b42941824f3056091b60774c29bf5d60c2e63842a96a880c3f67b96a6744804e4a61f6e190ef6758c14afc798d46c07c974d4a1b2a9e7240a43de3ba9bb1f2e7b396b4f7fa2832381ee0e395dfe35a443af4b4c2c7732;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57e9c81d1eac5900320adbb9e449c2718f0ed62d249c86fb481507b6c0f2fed01f7498c89836f75dc5158cd89a2c5a1fcc181881719fe59c6f8c0be4e3efe53c4e3e6063262a6ce885269b0b52d81839941aafab24daa8c92d1094a1f7f2d5039d713845795c141580;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db3fa63f3a60a1de9ca1fd9b269945d0aa822024d9527bd16c38f2401b210ee12573ed257ef72b111d5462bf0fc408c626d59390a01fa6d252d4a7a27ad17da8e80ebf01130cd65ce2bf68fd7a1b89e5ed905efffdaca5fb7cf700dfe75af79e04a224b0d2cb993350;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h24dd03c790efefa66b1e11ab1f5b1d422798d615c8297ebba8a086007123b9c5a91c3946e835fd38a2c3624e58554174ae5b9ae721a0b35c0f1eb4505a61f21cb971bba6dd89649c81092d98fad54b282b39ee80683c466522e4c20103997c45e2f78f07ebaf588d1e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d03c60e67732223d169224247d839bd8beb20a44007c999ef49750e7d9d46d8ca5d0d34b176bbc0c77acc936036b45eca25985a78409129a417f705abad7a76f46089c0444b455aa3413ec65001ecf6caa4fe5db99ba7b5d61d9d22219666c29c36c4ee07f44e12ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a9738682a1990be065a74693514dcb0b2480a471cd885aad3888eb0ecbde7d069454640670e876c043e10a0b4fc0b2f40d7aca4b9c55bafc113d97de207026c0370eaf0924f923c270d20a55692c27cd6cb40079c102e3f8760946298ba7f69f04b4682ec448fada7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ea30ae46f40dd05be4d6db92bd7c4c25549f3e9e1fca7e7c249862e5d784d4b848f1af0001bfa3a2d4ec55be7b0eeb481e65e38c3dbe93d8453492e07293fb9a914e779e6919931fa21625ad7d43f1d9232abf94c3948fd653b3ab85982d91fe614535f95ce0db09e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e747c902d1e911869443541766c289c54eccffb7f4440c5acdbfe6fc67443026b9182575d22e2be3446a4caec9788a054f5375f27aaa93a3ed3b0580150a686e4e5bef5b0e4f1e4a02d4b268be7fee4647e7b5057f9f28430a8722bb4225ef2911f6613588640de7ce;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0ddeb82f80e1526dba88ce34e59590b5657cdae5c5ebedd5dfa2b13ac512575c2e13d4d0c27a8b5d7169b3f848bff2730a79ef6480bb8b623b6b144bfddd9e1d27a840b9c06a489874832ebd34a91e34c5c4448838fc2792e4e686cd47e4b367817b420f938b5a6f1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183f72c437718499673668e29c16177acafc38a89216f0f0caeed8fc82374435137fee4ed3fce302736ae6efa51b78cefd58716961d496830194d724a94cb937f03090600f517981983b3bcf4268dd8f865af9dcb24183e8302a328774287ed62e9cc489b911c27c434;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19560409445d99c3037fc63e7a7277bbaccf72b055ca51c86463aeb4a41695ca05e041e5d8c9c0f677ac90ff631e22080a300d188aaececc64672b513df438860fbd77068af6d36246084a2916c8372ff0291027eacb46af1c2c7aae333ed77af9c3bf1435d2382081d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a4569de5ebb3fa1b7c1222abacc71a23cb1fe2584791f00e170674e7b22fd186714921d97de6be4564dab5d548160a98394e3ba0510458d4dab3819609bedb0786362e5f424eca35f9d68b47a4022fc713ac4932f2cb53c8bfb40149556a709bb7b7af19975b348d6e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ca7eebe3514def465b728913bf99dceef400bf9a39a1783d55a6f73ef5a6f06fa69d648708266ed73a30d97f991693b253460a6f10ec7d7a145d23466386a792f491344f53382e0b3b95cf9ec49770f7ec8b78411180a7efdd3127cfb3b177b420781284499ab95ae;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166bd608c08b51cca188c900f9fe91599ab7b9c2ab620294b9464b45d7a0a0a99146e0ed70081423f6d43e10a287412ba73ca7de066fbeb4a486d6a0d2d8219df17f19fe8ddc5ee25d238492983494a5dfebf85001bff980149d67d1b89c67f4092540183af8c957a7d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1775f9c15a262ab6f3275a808000ced8b29f54f72c061c43a624a628180c139a87b6d3e0d239bfed9add9e705e741892d3d1f0089778d49b3cfd80ec5ca2d592718b7f3523cb45287f62d9452d8ca099503bb3541702d5625e49f8266986029212664d7fc4d05f11945;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd42097caae368ef4b2a7945000f83482523903b232b4c5db17e5497ad25aaa4936b0921311d7f072b0862d19f64c8f8f9b34474897c1e061b3ea83dd43b829319ea13fbc5d06cf0fa9f1605dbcc39bf4045e11d8eabe955dda9792a74e0b3d70fa875e20f26a1c4ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e05345d34dbb3c6c465502a1031182997ea4af7a5ebf37b6a771eb3bdbfe5db71b2623f4f2fced11344f5241cdfb84fd0522e5fc2be8a19df190f824d185c90eb95c0464255547723b8dd8f6af9b28b594d0d480f8af69df321c96d4f894486d52769b8e7cf85a519;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1ffd898f967dac1fe1b6991ab1563a2f686670198abc603ab9c3460c2fc42a34a57dc2992adeb3031612a1921e671cc00e3b4f3ab0a5331cf12b9e72d2c109109f2d7d5ac81db53bee33caebd1a3e72482ed752211c891940c88af67dc78091195ccf283eacd7f964;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39728e682a1c83b2f894373a29da8e498e85dabe71f2cb5bb273c51bde368a3c5c48dad90a1064cd0d5b690a56db1e0bb7c785c3bf11675ffdfbc0c455a35dea7ae1c5c6521c7c253a557b9e3469745fe972203d3cc48c2a0ceab5fe3f0e7c7ac40f3327290e4a1d91;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6a4b26e2556773bcd71ba717fcb7a0625ab785e0c2df72c4d964f2ba8cc8eb688bb30dd80a424bd119a114c376503ed8f7a75e4b0c157eb6243686fb888f41241cef0644782aa03738c91995863f53c278bb891ec7ce0726764c0ee064e2c80f89709ce58fcfde4d2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5531fb32af0470c554dc93f8e498784cf310a1c518177ebed95abe5613708898dc257605a027b60547cb1f60fab261a801708ab97f2a46354bfdb9bec194386d285831ea76f16c06f99af32db2f9a50c66d41ed4ad0dfbdfe2ab553f42f3b3e609c1ba263a67aaab0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3afc817f2988016ead2721837d997e820e69db527a0ddc8d441f5a8c6f5b8942ee9798d73f1c826633d9d885065f4cc77bfaa6b6b9953a8c66c0263c00e2dba8bf38949d69e64c38d0437b07860b544690ce79a37514094e1adf820b39791e3bd87c3c0622309c1c3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1825b033caa109b4d5006b55466ea5c70b1cdeb5ca051989b5f3f7b243097764ef061ba78d85ce4fd1539c8bb5ea1065841bf9a696b1ef0e87ec7c0cd5577305ad23e9cb42cb56cd69e169e84f58ca558d41e60ab0259cb85e5f65bb8b930b71b410275a2343c4eec08;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11516bbb0393b6d603044a201dd363847003eacff1aaeefad9f61a610588ede8ab6cfb12143291b1b11dcdf590b1082dee64f1a63eaa7428ba82c3ce0d9c2ac0c011440722126c4fc7f6747c58da9e7d0a983a277bbf3e44423e38cf3f1628cfe01012009032e355db2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114d53bece99cd8609d2f42781595dd44b210ce6523cc1e9a0b2bf5b9467be8f85c83d214c80cea9aa5b6404652d9e77456973acb9d74049cd5712b51d8a9d2663f80033555d285a20a8accaf70f5890e1c82e18f3253e32204074a59e590dd2ce67457d3a55e95011a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1614daa889b4d50a895f517c664507056f4f7b9c26a30471312cbd34f990e75da80edeaad29672500f49d38225c5e6b23f99aa0c3e17d3c24320015fc3b17276602afe61dcabbd0cafe94f122e85dc6354f73e815b18b9cbeda4d2bc07a961a7d562178f37596d7f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93ba11c4b45d340f0b52799c95294a9fd73027c47a8ae3199fc5b86111bbf165c418c331c535cb80981ba1158776208177fdbe23690f6b41655f7e0faadb92e48e4af95ae75241404206d008abd6c5098ba4df56fcbc7f2c9abaab69497a83e770fbd8ef81e913ea6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1add31c0c6065f6536a8d9814f54f4d79511f70156005eca8764428447896c09da2a32fb0676d794934607ecae700a916a30013ef67fc7f874a6cfbb20f184a48d14bc1d3ffbba1530b1220aaeffe74170e39830d3530a2ab91f18cc5cc8b3c71fc44f661bd9272db9b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac43625afc40fada04c43e1c785e3c4cb659b45c11f60717e5370f09ff80c468bc5575021d2564b004f88797db4bdf69e77d7834cff6fc849300eaf81fa65de76f9458feda71bf228e1f8a4d34b60c2e827de639a8a20a9ca6dc7e6ddea45d4d4f1b61c9902c321c65;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b46cf1463061eb1dfc9602686102ce5cc302c3922c20fdaea22bbb041d9e2044fbcba499cf627fe2e88a9bf50706218c133f70918b98a327fb3f4de71b4f067a9d39f4aea02576acb941da9493cf117e936736e67d7ab455ef3149bf31b5c493dd8384f3662811cdd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9682122287f31795fec1b3cd973ca24ac51cb53b026ccd5b2bcff6bd77e8497470e96f5a28e6ef3f5f7b30cc7ab6b7970904080e1e9e58aa2c3e23de70534515ea36c7a7070210f7f66e0942831630f0edf89a87da5aed99a937ded0f767ab221257ec54a071828852;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc3d3a5c6167db3c8a7697f3b8cb35753f1c5528db7fc3dad4fe882a1994a7308258f9a4d8b84777ee5c0ecee5ebe7b7b5d2fa9d6c8e1da4ede47cfc5a3426d371e9d3b141b5b4e545077b23d66c2c4beee2ec03bd9f34abece2ec2fcf8cb2d44ae2690dde63103daf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f928faaddcd2a73cd6dc4333ed3acaee7f80423e8b128f0628248088eaf875dac1a912933890e48974202034398ea0baf6cb94a4bc2d7c249d05f09ea35968b3af1fc51b583b402d133807307302cc60b984046e98fbced09a29e382ad4d65dd8be6cee91b2e5eb53;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e4ec2d403617e3c36149ca8a784c76189246e7a35f34eb43851ab6737879f965cd7fd53627ff09a430b79f9b47978f2a6450934c5b81ea4b2503033deae9fe728885ccf9ee4847e711488e080df0ef843892e3d330d52080f3494d1ad9d4579b9dc9a1c6425a0ecc5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93ae2153cc19bf8e9de55a3cbc8e8db1e5c4bed7d8ba58d721f3576948314b32e5043a2f170716db8c34d3b0d1eae046288edb9c926a698f3a64d60208837940f3543de1880159b144154171eb73d0f31be731faf834a7a6e8d33e1e546a71df9f492a93b90e75674c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2fab2e228bcd64d517116afe1da8c4af10e7fc06b855106c2a14e9ef073df24ad99ef54bc08a448053dc54c95337c958ad2423461dc3ff4b2659f4e1102317396b70f3cdeec639948605cbdf089abafe4086adb28dd7970056a72841d9cb6757faf8cffdfaba589d9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c97247f62998eb84bb07283550be0c9e33075c0345d3df56ccb572c4ebca2399adad8fec15ed1d412482ffa048c3b0a1ad5b222dfab2bd8e8c41c8d59745c797a1e4c4711391e90405fb14b635e28c4339973b73a82ebdb30c04d6a211f11aea2c8646b4453cd316df;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb09821ea2a4aab9efa2ed7e1b4c82006614b4df015ae7091b0122a0faa3f915084e8533d70afc2dc7098b9558060872986441027cb11a534996bf718a402db1adcc8e045a815e8d5162a2ab6397ee09216e8ff6818ea4a0bba76ad18ea6382cb4a8cd01ba4b0a243b5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9313cf967bc32a32e21f37494e857942f54d8f5c3f12ed1264eebda6ec77b5b8d05a4a852e0f97cf92e9ff9f9551ef9f9db1bf28152225af65b3582f98241827fa8475dd78d12bbea07652f52ce17589624c8a4cf35fe1493e05100971cf4694923694218ca694295;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd1852d51a02669f1b0c355e88ea75bbc3c1d7004ba86ad71e8207be22129ad3bfa83b9283bc19167191087bc8c92f3eff68be8ee9e8222612035850bdec77c63954d6265a96094814666e2920dbafb91da3848cbbb3aa7014743463d73582bb1cdeabfbc8d0dd7b60;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6eee4d5e6edf39c78c801d81faab7de31f30cdf1f2585c5f1e4e48646530417cdef1b16387539581ed23f8457d7e2f6b53291a1a090579bdd6d2bb6b05d66d6cb4ecff2e782a8fc139fbf774ed26aac87fdce99f87618a9bf65986f7e0d90049491d122e512727a28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h535b5a9ce92d37d551a855aebcc11342d3944b5101d547eb37646a0821c5000a34dd4f71dce147c35a5636d92d90d8c25e650db712f224146d24f456f5e915dba0bbc636131766d142774377fef5d8050e86e9c48c0e2b63d6aea982d124a858f77f98ced49a349c73;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f64d2f7760696779bed6a05f4d95143b119f251aa83eb3d9089ff22bf55bcbe7dafeb58182d9abfb252175dd625945cb1a35baf50755048ae4b334424f7d849a6b0ee88187194c954a1a1dbcc698f17c5cb3508d103b39a6254bf2849fbc01cab073da9a94c598fba6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15be37f1d636e14bb0736b1a0dc4d1b574e1fe9d09eafad352f2e66a3b66b9caa847bfb93af3656ed879756d1bc027f187b01b0633ebda3f3b5e4645bddaeeb632ec254a7ef6f8b48acd701a755a68e8074271f71feecea5bbb883432910ee8f27a45e2c47113565fb1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c86484c989f3ca1eff705d91ad509117590cdafb7404c58ece1e3ab0525761a5a0561e88ca92cc5eb052cea7ec1ebe33874453f2e9919bc79a21088438e0c1a251b67f0cd860f6b8f95b8f7a09ec576bad6a44b7094c9a9d8b93fc0be86ecd23298d7842b513844915;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f68f9d77c9d6b0d5316e759814aa0b4e0d9fab19fb4428d26479a1443640b578e0548ae5363a6524c03d2da74bcdb2d611b86328fae7b36dd2c96cbcd355fceee6c09ab6ab8e8ff1b10e8704488bd4068a31a70c6319e35a5bba6210e35f343ccfff89f1a8972cf82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1693cd1efa2d36a5dd988bb44097d006f59a1b91a70207b21230837c63da003b5316bf63e4f183694b54c02ab45d31ef1ed70d28ff1e3b332531bfb37d5b9f680d011fd58b6489b7b5b4c40ca9e2f79c9acc81a48fff9197e8bb03a7fce4bbfac97ad02ed7e4c3c5127;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4199dfee69b2d9e867a063505adf63ac6d1ed81a25034a4dc118f8386109c409fca9d5ad7de3d7be07a7d18bab6dd2ac544bbd3efdc883e9077d85ca321117fac88754473f289d9096e3288f7986756dfb3571b97c06ce572b5fff9c52fc8adf254f65d902b3cc20d9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7a90ba0f67328166aa92aaeac0f5652c4f7a6c7b64467c795c106f71e27bd6f61464ca8cc5229523756d45a6b242cd113ea3c679813c975a75adb2f3254fdc8cf02aee272cb24a877bcb6d7aabe5ff1036210c11124543911a3cd82e7e6a1e2c2bb6b43fbd7fb7183;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6ffa3e59f5cae3865a752bda2b9a3e9f03a1fc4776ae5d3830e521d27299e9be586e8ad98ffd1fb700fa9a04fdb1b4874187832cb3a99612aa7b28a7cecf6452befdf88f3693834e376fbc22ba105532e3e6c93a29afe2ac52a2b586f755569a2d74d5aeda80262d3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c519e136f0b2fecc4a119a5c6f6fde27483f4b7b467a9cc1dab0a1152f1e629040cba7eb2106f290c8d585a76b200443f3f23c1d2b668091486dc6e2f64a4fe847ebd9c028cad71b5bc4f77536b39813d2d11b612b42bad98bd99bf2fe717aca020394e3ea6f5190f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he75e0bd0956d11b3e860948a249cd8328d5665910db19e21c204f751f732e6f0b079d9cebdb395665f8b626b5639167ccc67701a4de2864e375e103899bf00633a1fad072e423763fba790c417f53f8daf5261100a339d417fc4f12c2f180b1a749964aeefb5dfe206;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cfb38c990990f8b83878ccbc301bcb6feaa3f0364edf0756d704842769791e0805150e86f3b643bc56fdf6a2cab90e2ff50e690fb4ce366459546088fdf524de90e8a1c80495867305c81062a08fb8c4df24e34c22dfef9129407e8c0890bef82a01084904ce36e5a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cdf9b0a1f532481444f95d3c0617436c92a1aae55be262c66b4b951068742e706e7b4213911baabb1a2ad0e0596686d387661d1548ed9fac8189075a392c6db08d0a303d8b55f20e096734c96cd95c7e5b1b2b594142371f1c4cbcc943fdfdc826a6fd6540dd45694;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde5f152ad6fe6bf50e7917f45cca2d3101aaa7884b6c12b919fa307323c3886d04948df8a18f1e0d40dbeab6899b5066112a2ee6a80e1cd527201b7953a6eecba3403b9cbf09a048d1f51e42cf1f2551433ba490909c4092a309fac783f038e7c3d9feda8f35339552;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hece73dde9a29b004e08e98334017584f55e1b84f02b69e172dffd6b06b020504f85321549738a623a38ac798feda55821361e179ab18cfc8a42512dcd6a6ea9ee437abdd94cdeff586a1fdb2c8afe32918537af765c221f4ce7a50affff9685f0d987e48e033b8939f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7952961ca1d3f1b64da81c73b7f379b9388fea27407d94e9ca9d411e4528f087eb01894b3fe0e4606d610e20b22e9f20d1cf899ed765b7a092448ad89ab6ba157e64351497134b0fd181d6247e523f3d9a79b342c8cbc2960e35563bd468e2735a736be070107d8a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100a49ef577e8820cbd39426bc44f282e79f90e3fe3d66862b63869920520ce4d975206d43a9f805092562a99673c9523ea4155a158e9690a271b6dab6cbd02e67b896092c68cae3221d2f14d0043378cf79fddf9c487210ff99df80a2b808aee93f60b81d2e275ee2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc73da7fffe035e184cf12ffe6226a253c49d9c89719e468b5b031d7c8da8cbb8c97f5aa20fef388f0037ceeba6066576d98a145a381ad80936762cc8258b7da5f37f40f18eee8ba5c1dcbc72cbba639afabb26a58e635b4bae0f1e9df53a52496fede01320330c184;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h765c37676a66e9d8a9ba4f4951303547e883441c5fe23649c9044f22029dc12da1e1a375879c6d27802b04f225c24cac0fe4f8f18e8f40be5d7f76d7c906eb97b2e1c60b0938d2859291f188d837dc421c87a80b44d6be62f1d8c7fd4271ba9f9f483d4c8c2b20f4b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h281d5450a5897c00d258c7a26319a0c9ed030aab9541eaf20304a3597cb353c75cd3e08d5d2cd310e9e4b9d450a8bf3872935f491a1a7eb35f68b24c20ae54d08800fc87a09e93f019259bd918456cf0ce58a7a17456994798240bb0e80aec10642985d9aeb02efa6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hecd057dc19a639e5bbf55cb5b4aa3f5b6fe5eb5c213ef05f4b803082d21758304f2d850632921509b07b822ac70992977674d70b5b6723949b6170c5a1f24c5e0d51f206f034177334369ce86d3063153f2969b6450cd4d10037f85166f055ba98835b6c98c0cded56;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd66b3894f45a46a2577dc359135d82afb5eef68606ab7968aec96111806fe0a5b16064591ae72077b7f1f476ebea8cc8966f03d081984202a15fbd7a8ee4b48e793cd47eaf4a6bd85369acc71bd99cc2c2ff163f00d46b5107a06785042cd7026447a8ab7e3b7541e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde373292b1c1d3d9221419f85ada961946062983aa03296b584e1c5535a1f1b437da951c2fcd27510309ade7ba0ebe249a31dbc3249c176753d19e380d764651c589025d96db1d594a0c4d0f1bc4917cd7335e8264d736b892510d6bd3a13008b2017480279c9a8f5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h291a1ca823e4d50227aabda705223cb022942fc7f486c8d80f7a32a4f6a460b07eac8d31c5340248c87c9c737b654bd92614d9cb91870e846fa53c89e31e43f6102ca0f10814a9a4c060aed2543378a89b46c86db527ac3a2fb68940a0226f517d2542f39a1b8ce2ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdfed27b4939cd773eeece95c86b66744cfb1ff4915ecb3a2acb16dc76e8929d01dbb959921e708c7ff3689e3f99f36d2945285a8fa9772e046495c924128e04dc989a8c458ff5d6add9d9d62b34daf9ee64acd00709eade86c112afaeb854df11585cdab13a1cc4c80;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc2839256bf727f6826f1cf0e9a1b6cf24f5cc5f56e6d13c4167cd13820492301e997c2361e0b528e20420821251e1b3d1a973017a2f3fe01a228a306d4768de22bd967b1bda3adb4e3672540a6f80d43ca8edaa53795b92d3e43eea0822bdcaf611ed0ae585573dd8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3c76362baf03922adae756a5788d2949350c5430c06a544d1c3e617135faa5e170cb89b948505786afa23be26406ece58053051b94c57b4f39defc50e708d89b1e416308d1238f1686c3d69eb1b3e27ed8085b39ca506a6014d1c6d255b771b511160f94272a4403a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f182e104768c07c827c4c3f62ae789a48bbce829bcdf21a6ddd8ebd7760507bd7b5b778b36a4b3aee89bb724496a399507eeb5b94bfb4d1f7fddac269ae912020079322daad0777db2c17c9fb9c8f08e1e087c76fdc743fd53ee03bd35b185561a2865c8923a558d6c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef5b2a5f9e27fb620a4df5a60266e2669b54240b7001d7a820c0c1e169b4b6c03285f686f746e6f3e11f9f9389ad6df6bce0b26bae36f3035a8053e4cbeec6ad41850a2dc6ef4d3480058a72adab39a6840c9f146c44ed03042dee5f2d16a7bc355e0c375648260462;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18445782758f40026963da68d825464eaea30c1c50ad0cca4215eab1374a88895e9f015d9e399dd4c3c6f3e5a454f35750fb4bca0a9117470e980b937f814ddb5fc915ebb3d6aa1365018a95affa99b8692d010de795344d6ab41c0dd2e2bbf6769077639c912b8d7e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1750aa04d24dc59d454338381b880df00c14f2bcc9242e4286a017d2013af4ecd7778e0b003f1b5ff2a1645749cf213028914bab0da716b184d0f13b9c41bd989eadec1dae9769e37f95d4c79e1a0f36e80e4667f8afdffddbb93454cbb8fc8769d7f4e40c72721082f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112f777640152984ce2bb4674ccc6406f3605998315984207158b67ebe3c6ab279d2318c1ea9bb42e1ab4f3f79c5fb3abdfd019873433170b08b92b5a5b6b4f64b424b739d54339aba525880a204ce072b8d2ac2b69ea1e6a5b1897ce8df2d97e6e902a55385282a3cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6e9a184ae803b472d854fae0a695fb36a7463fc51c06045873d360858626bc7aa2d00144f441c4bc669dc0187ba460236da01cd6168d244f38ceec99308170fa38982839000f1c19e8f73134086ddc88885ec7c38da200f8563ccc18beff3ed7822bb63c501917cd3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132c0fe7cd7a60b829fcf03f8e21f2e7f9816a1c82478fcbcf1f4ca5ee371b9e24cd979cf0e10d2ced15cae46b90ba08bdb4c890853002fdccd06a512a55c36e6e23c91ee12ddd73efd4e8b37b5856eae1920fb8b07eb628a3f883816d7208fb107a04a6c0213b7eb1f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfcdb39ebe542d0e27a38caafafa01f4d282ee9a4e1869df5b413995fb5e736ae9a1fbb5e1e85db06323535e1a4211afccb79d56dc291a590945efc84bccc68910342307d08026e8943e0d8e776f958900893785899c4a7eb978e0cd25fcf01d583b20a94bd61f6cb03;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f9e42a5626a83611e2010ba7cb395f7d3cd77aa0f26d1bd778ccc56620245b7a053130b9c436365e88117f7dbe64d0e749beb5c61131af76db46cf1f53cd3713f2b5f873691f69b09bda46348a28dc211ea97f7ced82e7d80ccf84d79fc6b1bc8275cf604588500ed;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fb1a97074de32aa82f6f961eb93cb2ed97e99dd150bb9c4bc7ea7eb7c1040d044b27c93e608499ff6aa6d471d5f760379af78f23fa9ee3146de130c60a5f2025079e1c92942a3d7347829f20caeda51fa7a67220f7d72abf1df8ec8c3f0e7c86f6bd87d7769846ad;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1d4742f2861dede80b17d3ad055ea53ac9803884d8a5bc1c118f2d22adf300f68670b635531e8b614eb2759d9d67a0c8ef994b8ceec91c0aae72886ac25359f47ceb9abf9d120465826c31353b132d2ae9726b40448efa116e3f771a883d0c3a971f9dd3e97e3f1a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92ff6e684bb3ea669aa2db3920e0293f05c847608b5dc6679fd49022d6c93fbe05d17a38d3053ebd51d2fdc32491a66b959799a323d6000d8ad75add258c1a1bd7ffb573a653683c27c27e59b613b7a6f29f1b9e90ad2400b10a8f42497c8525bb1e569bb40bcefe8c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb73a3555f5f57c22ef43bb12916e0dbc97dd910eea81563b2ec5867fd5b52fc4817a12656fa41ae511f1271acc08e7892790823438a67f1962e1de4dbccf859bbcf60ff6fbf2e3c03a510351ccac619901fcbe7f4a8608d7d1166d14cc40503f1b2266f293c34b6cd2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b27c684a60773b9e419ce36ce1ab076368dea2c423bb462d150c11fa50642b3e51145028799feec920772d098f17aa93e1c20bd78a66943aa8223d0cf6ebfa43e9055965fc5cf53c0f226d1bc2f60b37ecbbe7c9a1dd77aef366a68e223d0a834c3f9a5b86ce7a92e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1733aee70dadfdb2e5ce52c7bb2f66407b44d8290f830ce4b8460340dad8ea2de95dea960e342317226603eadfecb09c6599581e6a56186e8c55aaeb9cb1b946cb2801a038282b2cabbc84d6967891a8075a2877fd1a1cab6cefb601649c5448b586e457934c41c0b47;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h569588e483f7230db64253ff9f56a54f6abc2103f6381f8467a93e3faf38827347b903bb5f1b5134b012023029c7d460537a02a5f1c77d4a0c1b90f68acde77d931e6fd49ec47a7d57704aa303c044c9247ae48981483433a0a6b8eed0f09b5d6c58a1d94b7d6b8779;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66369b7e835d0d188f70e0c30c367455139023f03770c6db42a0f72595e06dd3bbcfba4338f4d12c383858e201f692b9cdd30b7aa8b67b17feef925467b298160d7606db06c99ecc0e1743044b5b969bfd6a472265e9392976b32087ffb170464010f2481cfae84ccc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118ea1004285a0a08921848b413b1c6d427b6bf75ccb94be6062af68f31f5717dd3dff76328ac92f160f9c87d568822f134b4ae14d1d8aa69750a2ae477bdfc1fc530b440631c38e82cd2767dd068c6c0bc7eacf5c3393b420757255ebd906fcec76deec5140fbb4af;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f86da25e1f7a0ed8e85b53666a499a415d5834f265c359891e563af6cc729c9aa825910e75539405ca2b96c7ffdc7cd72c4aa0580490efcad4e01d756e6cfb000d99ecf64a1518aaa08f0f40b1cbf919da66d047b59447e9ac8d0e7a57ab48432f0492feac0f61759;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a52de490aba5cf625561aeb21214356de01e8a708586be3b710977888ff3b7e57d7c07bde00bf6753e7d12b260b84483d9ac83e985d93a463453e759ed2c315a545f11b7008e8286cdee30403dad0561cd20772d440af4506d70666d71734c2fd2770c81951d6e7c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4013f3ff9e73dd01eb2d79040ac52c85163ace5bcbace4c3ee608930ade91af7994b4fef04aee8ce993c3368a7763262bee8e5edb355ae9b18732cfb8ca34afb2e136c3deb18b133f01aa9d960d73a3ef7f6ec805e94108d044a4849fbee66d0778d701e361cac48b6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h704a2c47551c86955fe377513881109bb0ea52154d993a6125fd5fa02b15beeedbed5080757da55b9ed65083c42f1836e7ac8dc058d097c71e30a697648f5bc479d5a3ba38d67b94af280103798b4219cbd5b8cca3be1735e6b62e84b6a563801793fd2e5aa5592ee8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1822278096bf6b47d4a120e72d5e3fe40ad58909b85a8158a96f26128fded516306df83f66e0641f4334a5f30042d4a2c4755d92b3004a7da6f728833158f87efbe19449ca876d6616b14e5b31bdd3a3f0e733e98308d44ae0a4e101b02c00f0721e2a921b2d3f08be6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e16d3f55b1da150ed0758d4371b0faa52a8ed5346cecc1a6f73a33f68a06f1a038570571e1cec469ebe07ad3213eacc0ff75483afd9f0695023048c54af54dfa22e06c81823fa8b477aacd7e11e04aefd07fca518e9739f8d68569c47b917bd3d19f8fc1ba815bd0a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a81c44783cf732be5fdaf86e7a5e9c84935eeb57ac3821c62bd190ef53cb3f6ecd5feb3ef5c73b8950a4a812b167ee59eff9daf68e107344054bcf9d8f07b6b3fecbeb982486c0da79c85fe9a757cba4854cab0163b9f905ddfdfcca258e3cac52b0008fb796b968c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2258b49ac7faa00509c736d94fd6aa40f33bda44c2b0f54319fb733fa7c5d3efbf13625eaab9d0be37c792d4c3a92b2bbce357c301791ddca6394b2da62eeffab962e424c255e7fbae4a977afd22640dac2ce7f6855a45a561af7e339e92672dda297369f81f797b99;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d599fff1c2d060d6fee9f123967a2eb64a51119cec4fe23d93d38219351625ee8cce39897fb8c45b74de8134731732556b19ebe8fde13ae25c8b610f68434c4f3f1085ab5b3e2baa3279f3cd2a2458d566519f5d5340fd009bf478f39321c0d9cf18d0aac4642618e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h258298f3fa7d6b5ea932716d88bd666d063a57bf590029da1746975459318b7e6b578debc312bf5f43dc770fa8cb5f516fa60ff7eac553460eaec9076de9fe33377952fe1cfa39d4c1038d5f95e3292ab72f52cb7f464e008e636285da5ec1fc75e2e38b050e3795de;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8b8a6d0366073533e86a8e56537e09924c75a359ae7bfba2ec04c494be42422eaf5e3e9f4d11d44b574db674e4ebddd379d4b5ac07bfc134353255a757b165c71289b6a427275bbe0aa66208bc79bdd4dd9f09642e2b90e6ff8e39884f0bae13853909bac91db1104;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ad069da6ddc4e810e6aa083362fdde5b3f77108290e0f3d6213f8fe386f0de9927d115fed37fe8d311e7f006e91f9f1a765285072e1b5d4a2432bdb180e9f527bd7d203f8a72c7a64605650a283df5e3d011ced09dc68e4785b216cbc7d4ca90bcaabffb984538695;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ede78914bcb1683849fd680cea83b72702403fe3c7e6b3645e7a3af56c5fe201eeb7617c8f94f6e2bcc82ae2fb0e933cd4b2b59130b22bf770cd8de13ef28ebb01051014fa3eb5fe1d8c303cf1e714a770d72cad66e9cb2601e04536ad5e2c09ebd938f2cdf619bbb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e4ca32466d5f0695cca74d94a670e112b5a4329f9b5038200e6fe7375947c082b23a34969b5a827f1367edaa7d6c7223a689a96df58f75019acd56fb1bfa4eec4c80b854591a29642c2aab995a145d34a28431397d2e13b5102cba9e227b95f084c77307ad739e6d1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb2030bd1a4a24317ab3b65e839382469df07b86e69d096a559d7b68f12bb397fc764b6818f0454c29a50ee85a51a046cbd65d8154b1c3e21b96bad47d41caeaa067222f563a6cac6a3857c4883932e9d9706b066633266877043ddc3f4934f09cd6f842e12ab7e05b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cacc0608bbff0e91b576f2c6e6c37aec2982fabb575685b9e4d4f0eb1be6d607d4a5629d541522006f5e228adda8c9ba0566b995d93de511449b50ef0e3d079880a6b8a0c56d72518027c2d193592109b50708cec21df9aa3161cf94cc42cf49146f68ead2711da4f2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb049579935b003df033fc11e4bf7f16e0869e52415f55753a581869e84cee379d9ad67528176cf4a162135554e755dd5ab8555dc4d43a5efc6860b7b143c8e5db50e6969790332c56b54ffdbedb5054cfe74637796de12ed7c8b9a86093ddaa4727212c93eec4f3f78;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db14aeba787215e1e21f4ba31c459cb5af6ab2fa1e35d7c7e73d28d4d48baba846c51212e665d2a1c768f2266a18663be74cca55215de4be533e9ca0c71a702125e5d04e324f50f59d5dbdbbbd848830fa6ead9f99066687db4c44cb56b10768faaeb36428e8d56ca8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd99a96291d441fdebac3e922ff6c8ae3454a1d1f111ba0e17afa0f83e45c05c646416021a7a39f93bf331ba0bcff05bfd639379b7ba27c8be68a83df936351ad8f6426a7953f9c5c4421bd55de1c15e0d66a0ef1071e301608f5143d37beb436fb569feeb6f8a32bdb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a395e529c95f8ea5ffc878741a55a712c45c94d85fadc1e05b62fcd1c6cc39ad4b901b6255e00409b04f3c57b031f236dcd1f865877e8461dc2f8582f59ce2c0753208956c45a69f55dd9a80a49536ffb5b86f7ee0a050dd35f9f5963cc9a898a7c9bce6fbaa41ebca;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148d1dc294a18bc54d3e2563859acaf4c05af0106ce9e021ccbc033f41cbb4156f4a014a8c731a655878ecb7284b1a6ce4a260cce9725c61251ab53c9244355c5690e59af84361d9fb3c12f9c2c664327aaafbe1b82eb2cf099e1edc749fa935e6550019234a1266eb5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f999b9ca8cfee1d567fed920a3c49abc677f8b9e7247e9c4f27af0ece0621e073031678a456f4465a36075afc9de971dc73a633e42bd8df9c669d25928fbca33c61753bb0e279ddf5c1049280a64e836d2db5e283b44e225e8c25529e6091d9b9bcb098e741fab83f7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c515560fbd8e5450ddb16ce672e9f92d1413471059dd712a6e2a640dfc03d62ba1d01a0e07e62b625cc5bd9bd7d6c889c1b03e48b6701179ffb63a3a3348aeb7d01d257df83748de7f558cc1b16b5fbb4afbb4ba9b33be4472e8c16f13319ae6203eb873f0ac6c0bfd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed01b46186daa7cd5fda4ffc2ebca82da386b89b72b7ab946f2405ea62d722fadfa67f60b3a3b32ffcbbf4866d03c18e22bd2c00b402adbfa024ae3cab6b4e8a6d160baf6110d696f644e3f97f8640f6ce644394244139166b5b288f1533639f30b3c83589b7862a28;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb4995c0c5b38db36f7d5f230b18b206bd82a89cd80a05425b07128da2197fa1842a6ff37bdcfe4b8c211327ba83d128b2ce839bac28d6ec7716449373694a2799899714433268ebeb3901a2e3cad997268fd8d0f526a45786a5720d45ae9aeeaf8a843b096687f70f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11cd0a25994ab8d5feb552277195197ee7c3c1497b4bea29df2ba40c750912657b6b0fa2e5a8c953d841b2135a733eef5f513001f7c351c10b38ee7b9212677b08c3fc5de5320d3cabecfc12a977e5690680c53a1fe9496440fa954c5de47a67b46d4ec298a8402e308;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3164128cc7c5c1bf55a4dcec5ba3834e6ea2e63a794d2988dec40f9334387506827286a8fb0b17553cd34170c989470a8133a465113fbdb1e529de1269bd09ab0d1276daf92a47d5dd4b5c4e5d5de3ca2247494ae96cd0eb428e1d6192e68f4857a391eabf99af415;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc7ec0683cd5541b11d7236de2ea7508b553e976c309abd4206c42a589fe40dda99360ebb620ef5f61e780f7dbd13c0d5a10039a058a6470f70beb5b82fb5875cc75fcef8ea59edea6594749c49a96fe2d470ebc0f6a8fff94c468b8c666b4260ec5c8f5b0efaf21def;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94796ee3e61db46315cbe573f7b5c821c68b7be2c28f8029611535747e7eec92fd16fa7d4d40a6a3ff843721b0cde39a9a9d2b22924fbd664335997c17f8819ca39268fddafdda0229bf396dc0afd1ee2b46edef2cd565bc1d22e1423afbbe7e5eb8dff5aa4d6c2cc9;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h400db6aa6f1959445a9de82e6f2a4b5e51742c1168ce894041e6cbe5b754dc471bdbf5faf22bc98430c46496c8655d8b1d74a436482399224172ec1f08e7039c61cd6a3f073237ac9e853ce39bf156af29483385849f89f9dacde13f86a08c7d3a6d8525d00110ec07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd35f22e0e6974178a888d8ee993a61c234527b581fdf17fba75a7514a1295d76b4a8f4a80f15cfa94df1900fd15c394bf0925475c1a7a16cd0558cf4d3329fc1fc7850c79f90095c7052df1916bd8b7c81e06d6a0eae85398071dae34a6d907535940ad8ab0c2946b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h543bb8dcd12c801e126776b39cf82f792ad5da3adbf1764fe186c45385191481ee418c03472e6d930567b93f7cdc96d9a1e8e7f3a9c12ca382d935760ebcbae26c93af3fc27b9d9bf8a6d06f625894ad6bd0290f85b5e5e174bbb783f863f4bbbf6b9f7a3af0287ebf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3c0e33311e094f9dc58394306a7e44e92a1376237b0fa946c4b892020c157f07815a89f960a24c822b80fe7f5b29fff9fc3997f92a701c70967ec2ff213218e7dfb313bf4c498b434c183f64d4de035798bc13d40cf7d06374451b6510d933220b24b2ba5d699fa07;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1002ea1cd8f48abdb7a582f02dc889abffb1f4f36be08880678f20568df9392b4d69af6c54ba86f407d929596c4a4ef76a112839891e926b9dac5c9b51ed5bca530209f9c6a983ed22b760978ad97c3acaa4b830ab2e20f8d67046a02d5ed27e034afae6f33a32ca1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bea5adaa1eebf61eee3131c6bd36ece3cc322a7664b7d48d4ee20623ea54cc570b448d5cf094752054ec4e648a0eaf06e4a67e55dcb20f93be4b0c8f672c0ca5db22dee2495bbb2117194300ced4785d972aef69ea92337d1c0653c20612693f7b309cfac84ea0754;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5dc1178d6ad87c001419f41e5d9110b86f0eb5c550f0509c57fd2621e68d983ab9919104947f653df7e6c14dcd87c14166890421bf9c359b408f39466c6ce43dabec2f376a02ec5307bd0ce1a47a4e0908cf16fa1e401372f9b8e59d322b54036a10a6e0fb3c4351c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb69532db9e9deed4bf557ac4c2ddbd63e9963ffbd5a8165334aec35c2e6c0d8745e986f0dd336a8c74cc09b2ed3a81c64e3fe03a2952c0ad21caaaadd5969a26e6343a199df4be1a9956e8af7942cc90f11fe4fa1f429f572d0bdc81566ac799efb0e4f1da360c919;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11556b0c896c4a354a726e3cc09a482228a8a7d9da3fbfcf545f6d94df76d6f5b0aec668df9c62f080f776a6f5f4dd429efe5a450b27870297cd899cfd0e08da66b8c086b457df2d1305db3faab208b7920faed2c5624e419e76918a42576065eaaf3d4534c70021ebf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1527749d732129468d6b1760e4a3f08926c74f5a301c44f41d5e3ce6b811bde62c0a8c260cbfca764b86e5dd9d13e5b9b9d81e12856afbf26be319cd635d9356b9c87e513fb84d176ebf12e15d7c23309ac1d0a7a5254a0c27d61684b09b4c3d5e800780cf736578786;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e9afed49799f5a70e4b50e041564ece64d47396dc94a49dd01e4d27d35327967e95f2e13b7cfd6ea5dfbe591ebd3723879ac7522f341826ca1d6e9ee72b4e1ac2b74e82763236da6d6052c14b090b108122502d84a445400cdd458e1d2c2b80326d26c6373675c3c4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2337175ece849bccb48c86e0cbddf7749f55b02fe72cdd0374b575a021dd0ebddcc8fe4a2b5f2119cde495ec50070ce1d9a49b14053a69653948dcd60d4d6bf1be974e1b94eeba0915ef3ea0f990486c23c7bd57e8a5b76ae0f1289465ed6dbff6da9f0ffe2a195522;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb15bb3a07520ac734c04ef64a12ec37e4d906cfaac05bcf669bc824a6bbb93c2f9c9faed09565af56cb46ec2f1c1d00a5cef009ee99992132f2f50d59269284e486f56aabcbb8219d73775d0cd591499017d2dfb28b28677c0716420e1132ba9ca2a990d4803afffe0;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe76e9ec3cebe0da51e40286a6df90645657cb751205c7a022508280ab753321a0048128d179616e42a0674e2e24919c0330c39469e5b2d3d8cdf78ff3e5b72710f3177bfd58db7cac68f48826cf38b900ba135107f5c105a544bb256d4e2ca7e34cf08f8b5d5aabaf;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e0fbc0098382bb5cb1eef6d76840e56fcfe472a39b7c59c4cc7bb3412a5f174b5fda1ab0856db32109f85d62a8dbb55e084a69cc050556ff21d42bb44d2becb5e7ebeca50ac7c742c693f0ec93e8e70f922ec1465e4078065cc3e8e26af1f352969bc47f20e81c9a7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d8f44e0988e263ffb39f6d439f892ed1d53f6cba7e3b9ac3906f5774fbe5d2a59f1ac595aa013019d6ad7ff59444b540b48a36ccef288658f9192c41be4fbc7c7d6735a6ff43b8d10cc74a40df3a29bc54489dbc302a1e09523bba80cf1f1cbe6b4335cc8167917e3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb0a442dfa84219c93661e0f05f73cd7e05586b0ae2b995fb715229906eac55320ad7b832e34fc56d832055f7e955e620071a28f9db3d94f9dfcaf7c6f975a5a209493f2027ab5ebf9c94fbf4ce84b41dcf88851747bcc4fb568edcba4ce3ef0d5de8c2e3913ecd1c1;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18683be3121268849000e4decfc58033ead04b202963befdb8d00c720b4ad9d12478f87ed11b7285f40ffdf3d24efcc405b0ed015805cb358058367cf7b9fcfb23520ffc6bd6912c2ed160dbb31ebb5d24b1f81e02610161eea646b44bbec68791bbfc8453d3b5c022;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99769533be2994789ac442f46611869cf310c48d132b275c655b143295d4d66ca264f6a5ebef679dae9cb06b989e1ea832b52b39143008a9025756e974d4211ca53f9d504ca6aa6d4a934387d919e8530fce9746f49f8ab56a0f99ba9ab7974b897fe68c77d96476a2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc89a6e7069c0f54d87044bb111e7ae6069836c11c9bbdb0563e9ebdcab1a72e117bc2ceb116b6d7251ceaa745d8cb11d7c2fd2aa60ac4c8f98db5df28831ca88fc7c0459c9166936189b0599ace9671bd063394ba6e0da26bd3146c6aeddcf21d2f4a8524a18dfd253;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cec75ce75fdfed13ca82faddb75377c105d711feaf7b3aa7809f90b30571ac20ef542fcb21637ab4684012c318deb28328fea68b92ddc5dd73c59006ab10e3a633ec1dd84a5844322bf7a5a8aaf48ed38bcc071b6865bd10eb66d9638e00466fa598aa0c368a73cddc;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1116c1387d4e12e6714c8d7743c573502d1a7f029487acd5df23212f1d8c21dcec931ccbd42379ce01ac3e3294c0f08e92f29a941da54775500bc82ef1029c1bbeec3996324c8bfdfc3f7a7abc2ded7ada24fb5f6d19906d64b7a5692738e30ba2c8a75d4cced92b2a3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea9c3428a117debff031bb83a0478920bace58a9ea88aaa6a8dd4899f717a83443ca993708183db7eef226af0b71d93e34c64856cf32c44324e7f9a81c7ecfe63b8197081dd6f3f66264d547904f911a9d8ac92574f3a7a18b449d49310c51205c2a713969b9500906;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fe2fc4604b00b6383258159803ba40c02c47323e6e6a14c458b1ad33f21dba29597035abbce5dcd949e5fb21bcd8a5b157aad2cb22ff69709f59db475a1b9ec05935acbc1b809888a7d95f15d17589b8aeb66c317ca5d4800887e2b0b8623e9bf9a9910a39c16db1c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d89d7559749726915c206e915ef3130e1f102a8a25d7b94648954ece5ca015117731ed55474b95572e30d0115a36765d8a4c2095210d3dea79a8ec40c583d6ee180701d6a5e49434be88d73507d50f569cb864293c51da8ccfd25b96835ea7a83c14420d66f4feac4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc612f1c27e7e14cb9670c4a53cba2171a35c73cca4841be20f6c99ab52bc68a24e690dc1651bbdc51bc612af66f8f6c9a5674c7da311952d17cb22264cbb4d9dcb860dff3196d917ac40dbfc3e3aefc1516c33e996bd6f6ffc86e24f0dafcb80a8116a40381817cb0d;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6d78e3fe0099ab31ddd7d8aa5a70eff1089fdcee9f43a2190387bbef89cd5de940e488f3fdd045fa213e5131e1e06e9a3f43637530f50aae9f340a1615594224122ec73a5923c47b094b413c7b33ef63b267dd20f10058592e255e82bcb67ad73a9bf345ca9d6fb9a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e30d90b6049c0b80e109e1a8193fab54191cc3ee4a8ec8fb5bc3ca92a623f022b762474efb16ce19e428d0da4eb861d3c6ec7800e2fb4c07232be007fb687e1543d11bdfbd78ddb872cb1d623449116e85753132c09d80c7a23ef13618fe8b7cde4a2e85419a97e9aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haed711b1cad58935917c43f8d3df361b9e6a064cdde34cdfb804b0290138c9717cc8128ad5d2e8e2b9bb7381267f78bb5824a1e108b738a1d27545eee034f2d13a35f346710bd898634711d68e7702dc7a238415eaa3efd069be26babba0c773f208bdc777464c895c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h528cbd3ec5ff59336f6b9d3f8424874abad5cb80429899919fdaeaba0222950a563190c8d4ef2416806837c50534ce71065cf2ca767bc6524c9a34d9d906385318fdc6f9572d8b27d1ee5ef9a24bfba5de687eda0a10292d061476e3ea40589a7538fbefa12650d34a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19c0d4e26fc21019cf29eb213e494a960f5465c7483460955de514e45b014419d68e282cedae9224fd35f3d35c884cd040c9ecef23e7c3ef0f99366a099ef10762ef7a551369f9281ac65c9791e9f20604cbd0845f337e7ecce3a4e9dac542f8ff0a089ca68884580e2;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae53aa49c6e9e3bf1f3ac404501ae54b573be2238bdd22b9b1c466d41e2df259078e5272fb176be720a638dea8b8a32c33b5b20cbb16f569abed3ef3e706a13433e256b003b529f975c856ca48f359c32a2b9d45d0609dbc53b90d5e606f33691ad1e3bb471dce1957;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f377ea2ba3334076b089f18921c1c70747cd16b9e7976519f908b94317009319a6124c2d547176c4f5310195b7d00f15c2ad4bf1ba6b99de946d9d211012314e131bb7ecd448cce5608c5acec5929c3fed7663867063388e12469ba4b4addaf100517be5bc0c294b8e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h396c3e5e1041a6f239b9794014a98f29ce3edae093ef5d4e20aa52146573169157ed3a26ee50b4c73e752aea1ee11ee1f8b3c519a3e6d8b1d4c49f07425903950666c2d8c588464e8ab136eca89252ee3dd246311e1abf8d49fda20becd3f63261bf0bfb19d0efa30;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb86e502d592515077ae49fb50fbe4b1160af04063c3dc3c0dd159729bfb9baa2700ef399ff328fdb685927fad88753050f4d574cefd3ae3c92f344f54730275a4e5a9f978722613473a56bc71ddaf01e1638ec1ccab31ac748098bdcee3366f8f7144098e5a8c8317;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1efdc23c4645122bc1a6f4989d9d595d0b415045e8fc1bf69ce7b2f4282cb3b881b8917ab2fb1b31791163cf8ca1820df39208fbd1740ebb3903e414f1a9e418278fc6fac0cea07c45da82bf1ebbca18c7f59fe7287ec9587846ba6669c0aa4b59e32264a81cb6060a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c18d44117360035e2bf30f6277b5735cb22b81989737959f90866155b5d8de5b69ce773031a9740692d48c7231ef6d1ad8b0c0555a2c8a831831bf9e0eaae2bac44f8774db8ca6ad3123286c6fdb7a166403d4a9bdec2e51c46797d8f173effcd1c47fce6ea48795b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26118b2c69bcc0190eb5574e9f0e5b61b57802ca8e54ca0b00af0229d39086ad95d165c67879c596105d0e5c679b2c7a502c44a9f0ba0e5a967f56146aa526f4d75da2923de5f3310c48db3c6eb3b6384f78df0d5d4cfc2f339d3a1e83f1b8f35e995614143b6bdfbd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfac9827504726044c7f06a12603b7df273df566fede807ae8ce03a63bb505bb854e229ccf3a4f5a626d5eb1d304311c4dbe16869e72fab303274d9c7956655f5d5935d6106d622b04c8b391f5701e57eb97d0954cf4668014f24b9253c7b55ba26726371940750bc4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha122edc69ff07e94fd37773b685aeac8adb59409ca7cff2a6c001c56215b6d305227947d80ebb438bb1a58d5c5100b929319b76fd48134fb0e2c2f303e9a6766564fa95972956f65071722f657456ab6ffa438839b63676698bd0a9080c3a9af28b6b2e3a0cabc306b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5dd24b711ba0155ea140bb7ca937a6180f008010c62024d230d2cee711cd483be490d3e727244f88ff7f6e325c149dba5594262a200863b4289d0768538a43667f6e8bed90c2b89b6e16f054ed6417d5297b1718c7a0df5715e618fb80ed33cf40ff5c3179d172707;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3b175cd55ac3bba4aee7c3008e7370d73d59601eec752526fed6ba37a470c24801d2205eb8b16181b8409281448a1dbec9091201bff9e2b41bba400e311b51f236a178d508b742d57ecea1d3e0bfb18b9c22c52cf0704f185f6019561833b324806d0fdd6271e9966;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a66b423023c101b048d7987fdd2a980a6c6965fa9125956217aee3bea925c76ce8b04e4685893242e5bf013a95b816818f4e99bc4744d44cf7ff86ff0965f394994624e58e92dac5c089a895c4cef915209a4f31addde08f7eb40c8ced37e8a288260ea199d77c53b4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43ee3819f74aa95ebc9e2ccbe7d20536b70311f515d11369a00b31a9819a33e3b1cd28026bbba75842b0edaf139a1fa358800fb5afdcc0c06247f0b5ffba11600ea1014c11990256a780cd06b356db775a59737920d703834a303d6e5a657e1d4dc9139a57d7247e2f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155a700a8937c79b02e956ea5a6cae8fa88705933200972257fd87deffa601b482ea4585f0a951ab7f6d714973ef0ea7386b90efb7fb0a090ad431efa50185d97cd458a35087a03df9ba4eff2d64e6587b2d3725959506be5057071f1b9c746e60081474778876b835e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18b1446d426a8a8f0625a80e51d315394e431e104c5351b8a0b80c778c7106fc0343852b684dfde2f0b5ec3a217b10e34fc624bb54b7f582cc83751052cd231a69e71eb7d87f3181ea0ccb010a549beea44ecb755f587884cfdc7661001eb2eb5794bcc1acc75226c8b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h249c3815afeaf0bd9c2482059922bfa735e0c32f9ea678cf4f73b7450fd955a63daf862a58f8b9925cc16267d48674abd0af183408be3bd7f757944a0936a360774765da315806e73522e244f92211bda2f7df9ea0d4226f86a933108f4e1d3de1c577a26a7180e901;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38dfe9e30e9c172904a92681df332cacb4da6f3e96b32aaee225945798f49bd6dfa29600f1e33e2a0f2f30bea3732c07a1702642db3cec2d546e7d3fbcf40cc0ad46370df28d3d0f92f7824573a011a2600d517bc26fe917fb2fbd99c384b0a3b52ad7fd81d5cda9b7;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2d69d17e596103d716dc9ae6b32ddeb50a98bcd9a8df44529d5082db72a121eaa4a4a6389a131ec5a2e34e4a2545e1c8ec8fc92fd0ed9107af61b2e7b11a9ed453192c4bd2441364bee736796c855f722698fac92184243d8f32c385ca1a75257ae52cc371943d982;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132d62f4f0c033ea96e880a697e8b9485546f6e4236d0bb6f215b23a8f75079cc624771b30d852ee2c3986f4ea7e81e3461ff84954a598a64516f00868f7ea61615ea60bb669d41c5936ca2c9685f8a0d4249eb6146d79b2d3f8e6d7079e852ed507ccc61856d08e2a6;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e10daac5c82c777497e48c6b698cd9f9cef660c96906d532e216edebdaa515b1c680c8baa5852a37eed8ebf016e922804b3988cdcdf2ce5107e671f0f54af524f4876903470f008394699c40494518d174242046625a747881c1acdde7da0f3ddf81670b094df63ef;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a491040e83da90e935ea10e37c39380bcbfa12558e6202840885df3b8204b79edd4fd6a7429f4114c933e867cace2ab311bb30e86f5fa16b25320052022240f2accf482786010acc0d8acc0c1cb4090758bb71ca4bf50d3b82a9fd83736ab3b16204fb0d4344eed59;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f7a79e488f642b34db576bb28b788c29235687e9cefe4cbac3f0550c808f73d81c30c35967d09dd95698db560020e0767cc59c1d500c64b0f75f58e40137babd8bec521d18ca48b5ec7299fa5dd7553817710a7861cb6ed213a183c06dd96e14e74007c8646554c70;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f652997ae35cc890784ddf2790b9a5091b5f471390f88a955edafa079322575cc078c2ee5c310f38fd4638cfef5f71baf4e4d4d9b7ffc9000fa911f2a5d6c7bc7efe12d91478ed21e07b5e42f74c133567d38db75569f7742cf7fcced924e7aa887449fca6c4f2c82;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha1bedf657d58f9297e0e720bc7bbb8d37a42fedb03ac93a5b05c15fe6594e46d982f1dd399730e653a47b079f1cddc2a81db2fbc2fc10fb30ebeb17132137d98f17e7da1524eed41fd3ebf87cc30e0357b965c80553c20dcf620e9a195cb2cb4d5190458569b7b4467;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a007b5def6bdc8103ebac87117a37c1a6adca6ddd12561e428303bf39dcaa518836bbca26e4ecc928545426e0568959659e3208b9a01423d117bd331d3bcf2bd445f73823b5f107f9768a62394d328edb0ad3c3886c9db5e348e4f948d604c29fcfcfa5be9494a5d4f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192ff5729c457568de9f491ed8ece94bb494838c75d5d7d5f09f61848b6076eb996279c205776cd1909ebc12a90b3ff5198b3821abeafc8b3fae1d1d0701ecd429f8e30ddd0ba53e51b085404ba04a594e4fa4e92f9e9be87f39a2efc0ae3a106c75df14fdc2777b06f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h497281c72f2cd41687ca543ca08c3f75dd02bb843b79ca6a6f14fc39245a378173455b848c7f1fb8606a8e3ca39830dab9cc13c4b3c331bc1db4770f0f1ae29a5dbf6332d05c4b2f00720399a3061bb37565a096908776dab19b7bfc1323093c8ba0fb17fb66aa93aa;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf330c87bae9c944d0a341bd90886901dc91f966492b093b4a1372ff3820f0c92fdd777e4be5cf8c2a3352b96660ce613faf122402bccbb038bbc73bcfe2385b378baaeee44f798318bab67b71c21e92b2162935a48639c541042d71f9b3d24fe88dac5b9d2f857fbb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f42d1ac83025c0b7301714d1223ee6ec85b9063eb393fe75d364bb1a2be1efa139f5e0893c57fa2eaf92e49e040688ff30e2288b6adbf58ef218ef48129ddcedf454040b4a0f88b497a72f39c1ca007d830ac24caad1548c04ac17fff0d0e7d4480e4440f35f230e5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180f30eeceb9066bd3a144cad1f8c26b88ce11607c43fcb22ece361cbccbbcee9bfaa562ddff629aa7f0918da68394c9a354301afee1c145322ad034e6b2ff43c14a84b881c6cc17ab94805b86563cfb68f8bb3f07cf257fcec8b1bfa5a35eb1659d01eb9bdbd3d7903;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0e6bcdec3c8fb79f5f2eda8b2b744e9054c1eba92938865307a9576ae8711974b859a6debc814f6f2a61dee6a3c0037aa08eaaa3eee4ddd3ad4664d9e9db07befc4df7275d27e4ae5a5ed7a8dd386655140aa9f16320b8fba0835f01ea712491d99a81c2ef1d2206c;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e5d289959a025144db372bb10a4e88d71b4f82009e8cef15f59ad60ab8e5753d4e145bb7ef084140d313fc4c5cd1ab31066faafde8d3a51da95e223797e98e46a79a4fbe45a7de15ce9973ae5f0478708c491282f09c5a1642903abb643194363f524e35fe4fceb8a;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f221d96544d70bc622cff21cea498ed0f9afd2a684fafd061a5c2427198d97a7d7f1cebadb29f276efd7ac60e75f17527f443b85b9dfc935ec2eec136eccbe3f5cce2f5a194e8e6cfe9b854c36626563f43d3680410b0b4a6eb687c880cfaac200d7ef4fcff6a6c45;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ac16e5511cf77f03732253adb8d709bcfaed03c5350e5e84176da875c66cdf8fed44dcabfd5e065127bb5b3dea2fce9e299e5e0d8afd61812fece620b3714bbea19c45cae8d78edd1bf3e8a8522118f7b75136abe66e7fcd03515869afd64d92a55780965ce80c2c8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab1ffc4b5608507ad87d66d1934b1aa9bcd67bd6ab2190dd469e5c1373f4cd2d595923368e785687b5969c752a9e38bff9f55cba23cc22c9b7e4ad9ce3f18b9b558edaeda495bb1d6d67a8e68927fead51ac806de4ffe80674430dd8f089ccafafed20ff64bef94ff8;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18183c9c1fdcbdcc95456941545e4f035aaa44cb38f4a9fe029c1d0525ceeeb3fb4b994eeacb6c60288d7970c138a597c2b539f121529a172f59983fa89c88787f15d8484234ad56fe463c2254f957fe1502a76811cd9ad97f527ba44af3fcd282bdf427a56b73446f3;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17528885fe62b7d6369bea4f622727ae9cbb31e2c04ebceb453c564cc69c79aa63c26f328363da527bc10372831d88cde0f19bc42b850a6e86a9b3289a0ed7438c62b038dc0bd4d38c3472b225226d83a016a57960d0dbdf8e5472a4c5a1cdacabb492246a701ce35eb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1405e1da2cacf493b02122826b45f33765ed922fad962732e035e98e8a6c636e9cd2f4258bd3b95a3991e105bfa19fbaa109468ec8c620f7638186dba3a4bf69f43984d2e594d1babb291d1c6132b9d8d87441f4a4e2091ae6f533656450c1419e0e37f104e462ec915;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f87e1acbf57d0b71dc73f35318fa7423386ab8803c51e7de5453d3342dd50bd0f815b055cd4723ae480332432fdca0b8da9d8f9a35e9599bf1cbd4c330a1983137498d19fd14a68730c05c23ebefd5374b44027949b62c366b188ae6597844719e32ef7b5174a53a5;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125fa52f053f36ef9a442d77d52ed276d4cf31a152b87dc6f9aa6a309fdae8035a2a23f4f5dd71d3cfe7dbffcdca180f254782ff5d765a9e92cd1bb8742f3b24a62c07a86bc6fe659d3700a41e23bb7ce134126d420f13117affb419ec51c0985ae6b3395d47200f343;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6108724d86931b3fe7b529b529c48c58ce888dcebf3a258adbd21cb6577cea1730cfba9f21ca871837632dbda3a0a1c88b221a3d4c4b66ae7c1ade19bd03fd2ff08508fbc22c5cf414be2d95cb9e6e346e060128a3ccb3321c18178af5881b2f42da92690fb69443f;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65e956eda52d0290676159ecc4ccee4a13af1f407985c05c9bc4c61996575f6e052b4ffd226c94eb2c53d74962fc78cb6da068240cc8fd1a14619a399e7ffb7a3d917c1bb59f6c8618127db736df76b5e820cf95126e908cfcd829c8f181a85687659b9a406bcebc37;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3aadbb1848bda32b705a7c9087a2d9b7795c3430976e1dbbc0f3ba68b9390efad20ededac224977a47b1290b2144f3f8c3bf046e70617d1dc701bd4a6078f1c9e782a3b92a49aa602ce0f0b5544b8eaa7706dd716794e42312153ce599c5780514d46f3563cf765cd;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3aa42652d3eb966e7acd639c098adee173b4d3e84bc0338e0034d6ef69cb4a64878ed21bd819948eaa0fedaafa90b44facb1f6cd054cff3787fa53a0ff3975604eedf019a0817417d0d8a0a19a49937a0eb3da8f59087c29a3bd5c3ceea5b6b5594aff0321ed7f4316;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8badcab3ca94c2383ab495ac867c4e257f70c4d7dbd7133a2315c8df9060e69430aea6dda1ce77acf9986fb292df6d723dba777b150ff4dc750ec0d76ada594772a9e0faf97224fc79c1af03d221fed9591cf7a45a16a69ee5a5676ae8f0e53301005a57a9d06c737e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84257e28ef8ecdab4c582df2abb4e42903627eb83bb58d2eea03d708084d6187500f016b084bf297526f4a50bdf7c8aefc257d2d7d6cec8cf3e2b4a65cbabfbf1e6e4a29241efa95bedbb6b4fd06f145ae2651c6c78e065a817f842240635b880e54961b763781164b;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3f42063562b71863880f3f51aa8a03085d8dbe18df6fa8cee25caf54f80572542bb981c912ec6a9968541fd36fb59c986357fb335edde67d82e587c96066d8326bd4cf8f1230c721b8fc5ec2673fc3f8584b8cc31cdcaef8039f3fc4a796c8d2882491e371fde7ceb;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c2b41c3560299bb1ed6bd79b342070be7fbd9f203123ff266c33e9ca81dc5a85b793d1f43de916657cf2ee211e3b5fd4aae0d431bb9a0ced7a62bc8d1148694fba1667a2be56d87bab4e1992b3170b2212e42e7dc69217779b8a1f743638e166319f039d79b6bc616e;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c153603dd4ad0cfd574d5ce9dce66c7de47e4b6bcec129965e584a562e099ee3693e807bf7d61194c79e1ad61c4300a0be567a89e8818eb91944b90b8dce1665dd60147b55792681030358b129479cc3935a633e3184ccb6d2bddd7a17d60e036cea12030a14f34808;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109aad67a2174b156255da69d540f8077333cd735afb9c140ca05c7f1c795bdd32ec31041d3e4e0cf309c7697dd0e321cacd893e73b762881cf03e8eb12b5eb99746e5fdc5aa8217eac8ee66aea008267402d7fc3c3033ba12cc9b9ea417d280eee32d49bd71ae6e9d4;
        #1
        {src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f3340ca36157b349cb576fb9598241b6bbbb078111a7bdb1ff6e0f26b8e3c9e9828e68610a15597b6cdeeadfdb6ba54748e85255fe7a281f909d1a3b5cb46e056da294e3efc6993ee1afc537ca37c0fe813ec060e247a16d44b833d3f6bcd268362892af59f606570;
        #1
        $finish();
    end
endmodule
