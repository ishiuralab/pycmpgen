module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [12:0] src14;
    reg [11:0] src15;
    reg [10:0] src16;
    reg [9:0] src17;
    reg [8:0] src18;
    reg [7:0] src19;
    reg [6:0] src20;
    reg [5:0] src21;
    reg [4:0] src22;
    reg [3:0] src23;
    reg [2:0] src24;
    reg [1:0] src25;
    reg [0:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3])<<23) + ((src24[0] + src24[1] + src24[2])<<24) + ((src25[0] + src25[1])<<25) + ((src26[0])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd775732f8edc12473d0ec4d1ea8cceb7ca3042ba05becb83f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5e0bb87ae87a292483d22929c7736f399ab8122e5b791a87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51b186b2c0dbec58689dcf727326f197bc0297e1a73512b96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc59599a71464dc9239daf219d59394f12ea194f3bae52a381;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ce8efc7219bd0cc6a2b2cb1b24d7ae35b5b3df3fa0e38d06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd227673bd34ee5c325141b7eb7ca903fc77492feb711424f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7f5af446d5b18fa1011b9d44141d38a307373da3aadac1ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h313170633a93874f7cd1172030acec142e8b201ce1c509711;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a8d0093c00802078b6a264913e6efdac3db8800dabd19ac6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4048f85493a6293a0b9b0082a123a262b417b38b306d4c280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3678900d13cd2d09d9b5276f2a24e58a49242f5d7f50e2a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedf2911536f6ba859d07f94b7c792d91a810b1d1c5dde8f51;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d4ec0eef5b1ea2b41f750ddd91b3c5dd3b0dce0863c45ce7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc648df8585f0ffb1dbee49c63acefbb1acacbfda98ca1d6f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36f2cf3e7291afe7f6e2d1b93213909b59d9fa7595131dcdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7a82f7f078ab17b0b859ca93bb6d4a39a1018f36e3c96733;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4068deeaf5a1c8d13988402ef1bd62447902987a97dcabad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd721c257c21bb622ec43599052a64be7f881947d01b718fec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a35ccef095ad2355b4a82d1ffc3f2e6163664d096ce7a525;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd412ac7f89b9207037ac59fe2b680ced704c1c6900767dc83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59bf084fdb28fe134d6240a238e0232b6548b63df95bb0d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ead1e0dc71a309a2cecd8e7006b1c672aeb1ecca4104282a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec2eb69be28683c03cebfc5d31366aac81a02ccd8874d1811;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb061328afe2ce0c1d8983d084fe2cf6e18a0da9476d428874;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9945262b2a1e99edc511926fd50374da9347bb58bdcc2d29a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51adcd0331f31a7d08a748d84c7f7f53821538047956321be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3555d93d4721118e7975477a0f6e3a82aab8681e9bba1ad72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h159f85df9042f2d8416b84498a13aa787cdceef67bca2813a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c7675cfe8ce37b0b970b4bf9546c5b57d592b09d625abb9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd32970b7e221e1bc14fb813b4672d0d6fe856d051283cd11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6ae3769c91a90b0257cde285817506d7f9adeda51bfd6b7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c6a16a2b3c6cb4b0934a2590699432ae092c6481598af14a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99e847ad95bb2c1479cfd8c1fc9ba44bb9e594e3fdec2daaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h812448401c75a849e7cc4c41523d0c957b2abf163cfd4ab65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h637630e1beb83efe229c96cf92f808db6fc540943bf69fb0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1da1b12ca18e598b056995ab5d66f038845009954ca716034;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac4e54a5aeb583596e495c7b2d0fb860748d2738ec28e3833;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a9839e4c046df710548e1fff38dd718f562aa34cb40e843d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf48a108d31ca5acc1f293fc4fccf4c986ff00d5b8d58bc91d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h780959d97aad271726d5073ef2deaf267d0afc10e90e477f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec9acc0334f1d3b06778ca9e7bb9bf9e1dfce38e6c37d01f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5abe97fb31da0a875301caba95aeaabb80f7680d6e2157871;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dd95769d72a5170851b9e22da9d7390232194be4000b4d26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cacb7f1cb40e64c2b83d7615130c52cd4e5e6172273c7921;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89a0a049813be4b57069caaef956e16e3967a1348f1d1d11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he73bdc2548474ba776c80cc89f4abe527fd9462858c4789dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2f883a1e45458dad9e0004787cc7f77aabaeed12378f51ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb941e41fde37b0adf122753874d9218177d47773189fac2ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ca963ef3f538da505fed868918d558a8fb3fa9bf6810679f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a647515eb2256b18b7688dad83b53295767b1d16bcd7ffea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a7b1bf846c416eb35ce6c15b68004de36ce1e7327bec6803;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4e0e365ac6d1e568f00f381bb63bb140626e7b09295783b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdda0da55f75f85abb5bd50181cfa82e040be7f8453242dbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha13066ddf58ff0cd435df97369ea3f7452dbd105229fe9526;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fcfd90c9c10ca5bffec4b6766ae4b3f486665214fa46400b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67241bf1f91480dc52eaddab95114c7e20f9105ebc39b7eb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h998db4514e91657ce5be7b4476cc62a12254a4273ad5002c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2b7138c35d26a81c403660ec1ae5419e07d93d75f4807501;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b969aac6707ea0bfb8926fffa76167117f891757aa0dfc39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4129888d2814f39223ccdfe143f61f4637f8bee2b096adc68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb711855e27a82d75d62ddad8085a5f04d405515031725baec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heedc2bf6eb176178ba12aeccdf76304576dfdd157d8e087b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6061924ce289c027111afbf786a973a45426feae0058faad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc59d2c181210ec5134abdf46625fb816de9c532fe1ac87f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef79ca01ac95a5d279928e45790e3fae08f000f52500f9a11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45632d0cd0c0961a65c03e6dacead73baa631a49917d8e1b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdc4f39c1d02a1058830f3200a7dac812ff35e54abeefc183;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6a0ceee4a5cf3458f98f4a84e6aaa0f0e38872afa89bf390;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6188c23c07152f9a1300466792f2a6c59904aba211958b1da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa1d68d36325a2c38c9920c91337ede8aa79c74eb630dc016;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc64493233944b2d61e4e10d89a02023f26dc0c8bea7101798;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h790b053b259c7af91f389b7a0694d6b8e317501c779a7f32e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd22e3487758a17245270bd4b2b398b7104760b94e05e36e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8eb6f3e2587395da832c13948233534decf12899030bf522e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h241d4d3860ef7e76184987a7c73a193601b77ea230a29b44e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50b667408885c041425712be986cf1952e18e488304d02a48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2395d53900567149c06b994b0460609137a403cd967e16d04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habca3d961a394337bdfeded0073ccf023a030324f3397311d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cb73b906084f4bfef5c4adc1323f7d937c445928db7defda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h446c26c5993bc5ab1cee3b753829d6cb0db8009aabfb02e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46099b97ea952352e996b07e7a2df17160fc387cda2ad2255;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b10c8be88587c639346edaa7fca53323a2df3e778fdd4f4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h507479f0a162206a114b8542d5dfa471c1c636ca1094bbcc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he36025da9ac97f190935aef52c2712fab6a11db24bca36011;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he952aa9a631d00a6b95958378b53c2f486658489390b86e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6ae353be4d8ff21efbb96552e23af556fd63ad386bbd0e49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e10fd662f5faba28827eac7d50fa7bb60c874c925924764;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb91b0cb05734af00f91aed360ea10e08133a43098b2095f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26373886ed9525ccdab9dcec582bef5464db8376067fa856;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a522238fb4428271a7e7546c0829cda704ce57cf8ca51840;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb52436f024443fe958310d353435586b2502c2f498175c35d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ee85601252b1112f8912d1746ed048ee4a42e7e44a9c7253;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2c81b3ac021cb8f383815caedf6d256a41d0edf7f9460372;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb693c25ab90f71926aa8bb1a27c48b0d235316046cc0c2769;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd46cd3b7be1839cba75781d6d2ed3ffb74390a6b9c6513fa8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d31ab962aeb7f5345a89a90ed31b36bb0865224c3f4dd71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h353ce9d799445caf72be9e7e3479da62a0e03c48d842d55cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6561520b29ed8c701d44774460d055ceee49382f8c0bc3a4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaedf5aa03747b55b8e1e17117333f79adfb07ca7ad15300c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc034e15434af038633be9d6c5e6473ca905aca13971c6d10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcca6469facf2e4de922f1ea6beffe1c3730c28facd138277;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19c0788190a949a38786cb8ef72c03ae8eec81584ee32919e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a33e3748c2064e365329c972f48007779f6a967a72ca60f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf48c47729a0a4a708c491221289597fbd7adbd37c05446176;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9a256f6489c85fec340321263f7d1f9a289310cf9132e7f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf90c4a313076b4809e3ca9016f010aaef31ca015f46813a7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c319c21e7c043b3979a07ee7052da7092d6a12cedd07ccd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fb3db51f409be29eb1d3c39752af1cf23435c01cd46a70c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8ec7e14fec7e292f5b4ea5c6299af2222818dafe3a181523;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd79db1ca2adbe967f0feced62a3c207c70542ec804ab54a9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he93b88cb52225f3a7244321a7257c692e50a571de4f7fd346;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8940421d8f5793f59f048b43d099d74d5b8494c54a5f5545c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49980fa1314b915a62a3eeba7d7c7c026692fb85fd01ac349;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93521117448f28cbf7ee4e4e522da3ba0feaf5de2ca69d129;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h705785f2de2f674ab0b341ad5a87666182229a8cefd96ff73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc891211c012df61cfdef0583cc2b9d60de1488e66cb3ddcf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddbb33dbc18ecbb7c3b88cb8484071049f64ea1a35ad09a28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54eef30a4aa0ab48cea2e46529f76d437201eb51ef1f9d457;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc191c88d0edbcbcfb289469ff736b86854ed274280cfa263;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36a5312c03987f675a41e10adf9d8dd3d39bcc67ec9cc2c1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0e26e47604a939a909583bc928773088c6abf1cdb6f61c75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c07ee28d13a47da194fbb87c649d62275809ba7982e4a28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdccc699d068c3c20ac07d11df44fe8c7e3fa34650666fd9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e8545de575609e519e2768aea0d5a7e0ce9cfda7b306aa3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf68cb919fb7133965c0b2102615fe51f4d5868afba5f62970;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21effe2270b588a7f4a23c66d5b0fd63b678b34a8ce8360f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8d249b8f9f3fc0abde66251d46bfabf2208326a0cc45fbaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdaa89e4f20111f67ee765a0848a9b59fda0c4ae0c770cabb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h976194f121848c7bc712830ab8a103315a9ae7466a8692852;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf5859b10f59cadc962b1fd81c1b72b11582bc1b33a7a2201;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7277742269eeecec03c6624fd17db862eadd226ec1a3a735a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd73f8c177233ab958617c8098e673140c9a18c656da50e18d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5c2b8e59eadaed29f33298e72e118327c33d86985a1a0fc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h193eb91c687500d71acea7423499ac96c1b7d25026622c6e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9be798a8d5fe21d43f6d559c1c173378003e777b3d4ed3bfa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fc89fa809a26089cd9c88f3a8573bc880cf04c2de8e43ec8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69a9e4a5aa27fc77c7c7807f01e84c7b1ff959fa9aca2a558;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he390a8e47d170913c069901f4e7c8c58f4a715ba352d94533;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bbc38449cd5311fb8bf0944cff5762b53850d0b4bf19e00b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb1bc7f0389ece6e569e4b619b532425eb98e58aea8cf1606;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed0853f1c988968936560ee2327c0bae22c1fb219cfac5761;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8c2c63443400356222c9143e500af9c38cf6baf417ffb280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ce1dfc4604ed5973ac6ca9ca723e7fcb730c0f008aba5e34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82e6726ee8516e77e0a44e48082dcd0d551f3dcfd3af803cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62f56e0c2e488181912a7088d6bd0d5e66d6fd4dabb509172;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb13f92f4ba732684ced23115d9ec461793a8d7a61f88feb7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69a09b420a09f88a1a718aba7cfaacdb77ee82019e9f42f02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4ea7deec6fe707c79dc80ef6485ac2ced8220e2176ef0b43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3965b17a6fe84322c7101c6a54cf877dd5db933d79cc315f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62a2f8284efca4f6256a80859fd6caba8a77e085fb36dac4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda1b76f8a63f84d8d9ec05728950edb4b946779a5f7821dad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc41dc095aef73c52e26865eef89a993b83c0ac52e0bb29d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb9df47769c8b6bf651b639afacece561598ce95fb906da0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8f35d893a34370e0f870931d8ee9831feb31ee2514701cbe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8b99f4845fc3103971d2db2ff4bc366711403c4e2e4b91b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6475bb42200a03060b0b18df38c0c399bc7a6ff3bb3c95e18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46734c754097e3519635aa765360d8261c034b92c49247b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcadd1398e2bbad715dbc2ec3623594cafd4db99abf8b6c330;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ea014e4249a4931fd6192afb52f6fa31c5fe5827208adff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1e0b36c4963452bf60e7f5a274c86ed05a25d8e26d2a8143;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf17ca002b1d950aa65a90e267453b5846daa344d0bfefc04b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c5800f477967cf605f9184caab23ac8a506d6aad0a0321f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68da2c68d0b73550ecc04146a3256ddcba09463785a3b2b19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb08aee2ab7b6f1bfab41c425ee892f9af1015fbe375cca011;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha61f71534e96d957978168ea2949a76a047abefc693c8d32b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a797f0db878606d198f196829fade82600749d14eec9fa1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4397e526cab9c678eab56513f90e7cafda520ead81b6c385e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbee2b853a474172e3d05471ad729500fcc1d944d6cea59a52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h884678da3b1f414ae9fc005d9e83904ebf533eb3d4e9eeced;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24f319b3fd7203a37befa8631cb4cac85770caec8a8d27ba8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73b175be4c5c43f9ddb20dc6b7e581440316492cfdbf1e7a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc692f2bf5f7dd29fc47c1518bf16be404a4cd9b5a237db56e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6c967b9c446e114598048b383689203f775bac2afc74c197;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hace77ab8a8090c3dbe5ed05eeab547f78b241fe1135be5463;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96d44cdd92b6d655af49ff4fb322ccca5a6161876ee4db287;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e4e1a67585cf87f5556a7fae25e6d4e3cbef601ad8b2fe25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8dacd2fc69d1f00ee956582c4538e4366311bdbbfa9d79ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4ab8c0658d095e806a1fa0cb3b563e4d7dd555b2a0d5de21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d390eecf14d5fd6f37718f099b2597c039e5e042d40ba675;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d115bdb842cda0bfd777f513f46b2ff4e82196e3c7e0e369;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecc01af931799c84a2d0aba8465d79773964b56f648ba8e8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2904478ae888604f42c6d9e253b3c13d10b249d533750aa61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7623124026d9b195d7f2baec9721ffedf76f43249429c1661;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ceba2281fb76c65a04ef5ccdd510544e8df141e6fa81a6f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6beb74a03e1eb7881f744aad904c53858590da9c5d3505fa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68dd34a4b7e083d307e5c4eac9f74e1abcfd7e2271c9b1214;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h480bd828d3c012eb2fc32bcad07cc44f2c67480bce7fe6d2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc17421cd58652b4e2dd5f65e413e56693393168e3bd724c28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16d92c3ec9d4331e17580011d56e10d7342d0a02db48d63bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4f808ec0a264aa37822e0afc99c55553b277ebab27f4634f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ec0e8e2a13e73349f1995a45e018f6bf97c8c5a64f02a2a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91e986c9c05870c065ca753a25f2023dcb1a3ad3f753a12ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c22327f23719da188ccc8697b7de900e02a822d2fbf61957;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2c1ae67c5c25f0d56ebd06021f8bab19f69554f6fe37637b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fc992c412fc33471dfc18300e38c9e3d7cfe22c35aae8454;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h572e567d211cded2b6e683df3baba66d0e093da1498a669cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0ebf50b24247280ff3cad4c89a19de542cc9ce94d5362a93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b03fb05f586ec886f324a86461bc40fd90be94843a80b2ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef81a7dcfac5233b556c116141e3bc728d30325333babe003;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h193b03cb44e2cdd2dec5e95f55119f28ce0ba4aa652321383;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he654c282299786451299a095baf120a015e16cb7089c99968;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb24a94552b6edf5f2a5d77a107ecc457c6f1ab3d6375e1e64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2e1eafece0d3b44d9f872c4cacbe2fff9c34380273b8c866;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd84785a4d58a20f96b3d006e7f2719abc034dbfb2b7be36b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32afe25306f1e923006277e48d1088821ab6a1d5ccf09fb44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd0effa5c535957b79ca2cf729da8effc2a5e1b99ab08176d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he179693aefff5c2ec853bb8d8b82190eda43910b1102e79d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72ec322423aba8d2d113f1b55de9db607ee62aa91bf9dfe08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf43d8899713982569e9aea61975fa023ea14226a43077ece;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c17e5e28c94ef98e71fccb771c3e8842c1e02313687acd2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8c969b4ef77f453c716cc746e9763e135e5697f4ec5eb716;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c9f35fb1090a1b77e8f60ebb5afeb63c5a9c1b52347c90ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b3f65c2c35adf92ee36bf92b15535b2f4c445cc998cb92f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a86d3ecd164307a9bbd777e9ab27121198042a8ed146c3ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c8c98af863592f7c71d6e31c9bb9d3a638e8f0fadd772b9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45c848e450742c64697971aa8329f9f71bfe4ef0aab3e089c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6e73ec5c4f6cc00c3302078d7499186e305e74419b58add;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29344bab141ad0eb427562410d5fdfa0344bdb29f36f56374;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5fd0e4d0784d9df86008a2019689df425c10c7a5a388ef80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30215bb0c15d0fd8105a4e0605b36e606a0acf9efc9ee1e0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28658ab48b985462da20ae25a4256c9c1203e75ea53d5c0a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47f64585963d4e6ea83d5005ba96e0db464f8ad638e9c2b4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4133778c84e5e7087e8b94002b917587ff946e9439e78a11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cdbae48fe409acb95b3906efd9de230d987f7e2e5214a9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha28c22dae22b37d1eb286220af6da9a06ce8774ed29c736c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5cd184ca423e9db2e259e3a66e1169ae70b40f9441838d4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c84991c1ce9263435c6ad8d72d312a483003684fb61ba42d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c0f87cc83c176286f4f46107ccd2c156d35a0eff857944ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19004897825032c087a2a90cedd33b678cdd0e5dfdd3999cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd556c372e36b6b84bb2000b94dbdc6fcc2a3d1365c148493e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd63a74a4fbaf56a2c7469ec3764d1997301cd78d012a5a0f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha03991c16f1e6c67960c84a5fa459da380ce32ba12bb15b29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f034df7f93ce63c8d5eeb42b684bead4b1388f6dc3c076e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81e33d91e064d626e0c4e30a8c69eb313f36786013e9e5677;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h711946130de55979c9bfdbece156c9e5f6b708d9c74e4122c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h639d3ce69bb1de779db661b06dd22213e6163752a5e73e0c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4223c13ca10233bc52ac87bd9a7e9e306c102923ad08bbc34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32db130d8c1ee9f473b88bab2bf6f15c6dd1e2abd2f526a2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd34ff8ebe7fa06e87909cdfdfa0f133a97ef2a0fa921ed7a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36249bee0045f18891e6729f83b80461faa3933c17e968804;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25b7cb57c2268c844972fd31438fb6f3317051bee4bcc074d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45ee7d25ece7d8dbff00b7cbec0b557a9b6acb5c1ad349932;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33cd9f291943a101a0683f52050be3594656f054fcc147514;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d6f7706ee4bd1cf5fdbb704a0f3a4712ab5251fead802eca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc34bd7e188287945557c2b571c04f04d29055846fe36636ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h835651d91d0146cd9dddd0115194f8a0f4aef3b0615e54ad7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc41f992b3afb5c488e1fe740235cbdff85d83844011b100b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc87b3379439f63feb6cd96a75357a7449916ff855c9ae5eac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he70ac335fa800b98de19180b820b52c98e06bc801f110ce11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c44868ae8eccc688affcd413cdd02ec1b8bc54bc799a1088;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb21ab90569a2b0cf38732eb8dcf0f09f423db0a0786254057;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8df253be1cd902d2a9dcce455af0f7db039e4bc7e1e71a07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d8eab85cce3c22367c3a9b76fdf234fcffd8f4bd72baf970;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he070d21ec6fbb441f91658660d8ff5f7cd99fefe8dd7e7e35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h226684257a61bb7f5a479ff6f7cd5f87189b4ffb4160b80d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56ba335e499f4772f8c82a2dd867ef3e639da99e49e586431;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc99bfbd96a7e9dc40b4f531cf340f6209f58b466cf715c8f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0eb0fa6bc385fba809b47928bef4ca01483c852437ab5870;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ffd8daf7bdaafbe3460a287e691f1951c2a77956423d88c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ce2a61f7472913a74790eef0a39197d3191f50c63ba37302;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dff883922c59f27befa2e301c09b1940e3213a72ef007ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc0787954070290dca4eca630a21011611f37e595c8269297;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12933c0e483445fde255e94a1cb35a2293b43c54be1530717;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54699e23a1b73a1f18a3a837699ae9da4fd5425b772051721;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2f83fd91215b7544bdff5d4190020297c1b85ed3c79bbca5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55e490487dc6b68a862e6f15ec88d06484985dfb44c07d8b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52871b7f61d58fd6e89a113d75a822c66376cee04e4bf5410;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ac0b32eb4c0f0c43abbd99d5cb6312cc8c7bc8591085ca7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1e64c0a7eae605bbad83c16a335dc3e6943b217d3280c3f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa05edfd984c8a54aeb70b5f33d93b9b61bfa1f7322e72dbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he636b07d69cb5fdb2ed48a8e4927fb934c7384d0ed471b6bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c2c57b01fbf73484657f7d27da3e83c70d7b66ed110609ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3a6f92cd253f1b0270162ed714ae4c9f6cd897f9f47560f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97c819d39d26292b94afe67be3b1c7cb26e678d6149f987f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7b546401fb7f568337a66644f4d20a1acb3d5cd15d739028;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ac87d51091e3032ca8b325e5b2a2912303d8d914c8cde18f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70bade0262f23b9f3ec0279eff1a611085634dbb0852990b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h599d503989b2db77f3de8064e7c8647ffe5915341f96deaa5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ad3cc1e2a9c60fb1eebed793564e284dcb0ffb22417fab01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5daa3a1ee688c805c0d7aa1c72b73a97e46fdd3ce78c0e5ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b36399c4ad4c21322f0122c72b0f61b91f0b898fda438513;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he45ea4a57b4c7df5db50f92545713c47e06c274df72ebd54e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ba10af5f3d6c1902876293b8c9e7233353f60d582f69d612;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73ce20c3d82e4e631f1c83e945ac8cae7fb71ffb343fe416a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb571435136e38e25ace83c4a1e9507f70cb49be0a7402a18a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dcfed0fa23fd84225934dd0387962a5f3b1c1608f2184c5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c80346dd787561643dc5c0d71d1759dbd75d6f0aa6bd4311;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda672c32cac5bbae0dac51bdf8ca325d7cef5458faeb01e62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53191f2c3c840e1558723732a287cd1ea210245a2acea4b23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde9689da939dbe58cb36fa2de9803abf3de773da7e265c1f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0d779f77d4b0c88aa23ff6ba79776274a5ea7201c114fbea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e2203d67a2f5e831cffcb6bb08b25f909362c74191ac3861;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6575a55830076229863eef100296f79feb32b9fff30474ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0c29fea31eba01b8870483afa4bf567017ef7d3a743f759a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he38ea13f2c5515eaf44e75147bed451f6f186601a1b106970;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea8c7416d32c309f634ce8a55747f9ccf4a924297782988cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1860ec5b216e05477fc211129366d06cd5d0640c4f1aaf966;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb178f06b85941f56dd315efc911c82f3b98d6be3af4919d06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea4b08d39ec3ab0050aecea43c8d2b7bb32c8d446fd7371a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a8571815f3a140c4b63bba6cd53efcbc579989f94869a477;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfacca93f1ddecbb4cdcc53badfdd706d305d679f29bcbc37b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4863c9a58d0371680489cbe927202a681f0b9c2004090745;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3077661179eb33b17b2514fdbf80fdd6d392410f9c203f636;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcab93cbda70387aa3d005d151e3ccc86b7ba6e2c9ac40c27e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h302e90399502084b458deb52d5ae08d7165ff60d682cee4e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce2b08843c7bf510e30f4f58a053607dc183bfc1bafe14851;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8d7ef6b1ac619ccf97c74680b7452f73fc74f5a2aeb9d4ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h583a511e88eb76abbfb9ddf3b246a860fbb30a18e82692fa8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cd6bd95015ddf0473d98a58e849970a855364722b7ecddba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h742dc392e354ee344ce3fdd89a3091e3914587c1010e15918;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcebb77cc13d3dbf4a2860458169689f65a8d2efb2589ca131;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd55c6a2511a97ff47a5a113a69c836d0b35ac400e4039cfe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5653cb10a69d3a88f4fa53a508f26534ce99ed6c94cc9a796;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1224f88befe886578c59332becab3f9eee4c62d36426b5d4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6dc8eac8ad8a37b75ca423664cb8d34017c50909574c65f97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3900023756603b8599e90b5929d4aaddac20e9af61e95d077;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbffdf073299b555f295631b4e69d2c0da7044900b4a4bb68f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38c418461c8524c494ee896425cc98969e9c5bc891cb32a72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7a350324141d3aec94d55e97b5fe207ead941c13f9eef761;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbceb4b69be3eb31c02b3d8706fb95e38db867b296f72b7a3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf4fda5be014dba13db1749c31cc912bd0eea6e2d0d8c4fa5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e29c5a693578fc97a4cbe6d68ad57fd88fa7bee93cbaac3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77d82635ca07bb9216a32b2effbf31a788c553f79e8ab8352;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23694c52cada967765b97b2eb84cbc5ae35243c5dd0074461;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h433566bdaea2870180352801e309c2468c38df6e6797cdd02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc26abda10649251404986894990bbfd2d2537accdac2271e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27541be08169ff8823320a7cb4f9ea978237457dab7647540;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9863096c15351c6eec289c4dd6357c36543d1252bfc0ee4dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f9adaf2d63915adaff5416440a92479beb89082752cfe327;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8dd7dc263c46f461618b85d1d6e86eb28ca498550b0ab7478;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc1fd68d7de3d1b5c491d78b1761450c5679f5a19e1b79539;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c05488ffa4b7acc668f34ee3b74d7416b9c8bb7a750ad62b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3358f6c188ea2119ffca1d645f3efd007831e2ba299700137;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1759cf6816a99d82a0e33884f07e37babf8e10a8de59ff312;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9c056369185c2811ce9c472492c5cec4f6bc13431d5addbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd43deb84f5463b544124b62a8259fdb75ec63383b61cf16fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dc4c09a38437ba867d59f4f1c45f94e7efb00f4dcd7aed5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he171b1c5fc152a496d927d2688cc449e085995155d5df9e64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h139e6f8a298c235c77731028d7a3035c7d3d0c46f4e3bbd7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb33728ffea130dfa8d1e9c5d38b117b2a3d717a7494f596d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h225f310ddec7194cc591e52bf7754959bbba68ce226cd6629;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6ff5902c19064d62c0f890483d840dd84b8436400e9c1f48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6ead1ced96d02c16a1d28b57a9bcf8eb1944ccad7c78c212;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cb3c13d8308009754543d322003b89e2d7461d7e8cae9e44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72e2644bdf4081b7b33ef1b676fc635525d4da06b1e228833;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd72593ee6b607868f19f218eb3593be6b4eb98d3652ed87bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69450b2900da98fd9ef93aad74a416cc34f931e0472cedea2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5978a33bee3d4faf85c34e09a48a797c354c894e4c68a57c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfaddfa9e9c4b4b58ce6b414eadbfe9520242b159322d42e8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdcd0f5b9f3a571d8953e4205bb195843f8beee9ab1b8010e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf92fce8352fd32006aed71a1ebeb3fbdd854eb0d7e870a74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa8bf2ac03ae1c2e421358db57b5f0241583d885f952677ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5edec5d3d95ac11923002b55d1237b8efad9209781f3877f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f48c30679ce25d811510d1860c8899fd7627e45a460c3c5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65703b520924ff61e6ec662c3d5f19b2fa4dca18db82015f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34b1e8c5f0793a8a0bf698b20ba11ca8ad7581e8943d87ed2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf75eff0dd87ffa246cbf40e7d56f78124adc62516f022ba2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cafb1cb5cfe09e5f25d70362a9a5d2e884f0c2bd7410042e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadf54ac9aad65c544a14a82ec033c025582eee21bf3bb816d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc08c1f7488a78eca19c4cbbf7cee992e14e56a7de5aece614;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54e0778cfaa477ea03d312ce05a38a1d20f398ad470f3f78b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c87e435708a0c7d5a6cda84f0787613a30509738d8f2a6a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2926dfa134311d4d573729b26a3f92bfbc098f306a97fae65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h847bd4d57dafb0ceeb6db9ed52c5487296608feeb91aea215;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb91d2da5b8d7cfd47889eb2c947664959b0be5ca5fd78a312;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab1bb86fff10d9b598828c413281c34c2b5ef62c046840cec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2730909eb831602f0328f0bb56dbfc70a611d7cdead827c84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd53fa9288dde6899efea5c0f53403e99db361b8399085730;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc91e873c60080ad95fac487437996e559ee6ca0e77f2605f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4e88ef576647f342781144807f8759815c455644c1b484dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39703568139ff7cc3624f15f276a5dc501da910ce7975146;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39496e8024bcfdc09942e6b618be77bfe367a4b17ba0162d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8252a5cffb481b50dda9db7a9b4747f13dc6e4c8691b5c181;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed32e8c65d083e003d985b163374068ff69ea28fb40be25a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e8c5deed44ec24268ce2e1eb215da1ef6b9ef10fefda805a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5572e9b51d999babf0fb54ea95e349991d75b21b453c87e82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ee7739ac0763687f9dc947391dcf2af0e184e2c1a10862e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb5f6d82aab35406c4105d60d01535b2e6c4d55bb473bb116;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8bdfaf78a1ba5d17c7f87ecd253a848a73c2f3278c0288b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a5984d7b0a0ed8d110a552735be2cd4acf1cdf8b31615fe4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb04b9c4ee323b14c9572f655285b7b420a1e6eb764d1beec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5da427c418e37d84d3da9f5576c6065c5a07189c219aa978;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff04371dddf541e1de504f657c0b8a5be1698c6192d49bbf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d68a82653106ab30a415e9a83dbbc84b5c3b8f1099112bf7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h692dcc9c6bd59ab1e4f6acd5ef434e8b1f6988e8452b7c27d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95fadeb251df45eba0b0f2c7fe713b6c312710ef66c1d3926;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd88e00e686c4cfefc5600b1f829a557f861fa9e022d1ab128;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7505c31abec16e4b5587833cd79be7de3078ffc31b19632e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf89c238fcddc874ca7542848c550e1a348e521ee730c9771;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6192b6fc46c287e68ec096d5ff5f292accfee39ba5d6f2d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32515bed35a55bd3be89dbf8091c7540155179880a317d655;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b128e73a944db73bfcb5bcadbba4a9c075601185b46299f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21162bec8b6ee8a55d22b59e3f1433da7ee87740061191d54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55a0c787e86c007244d2e23d2e802bff7b61dc512a6f3c73c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7def10757dbdcff2f02ece496dcfb0e79894d60e764ead1c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2976160168cf48a3fe346baca18b5c345551925ebcd6c787f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h416fbd6d5821d40f8f5952b5b57b937e1ea8f8f13bcd5370a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b21a3c5c12c73708140d5ed03906e00be48eac756a29852e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24e081e9920a262940c7d5c41f8381997ec99adda91d7e3e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h425c9ce003991505ea951d4ceefce3c769b5a3ed1b921e6d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5164eb27db1a79d5d26e2f06f48712a37a51688d1246e24e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12be9321c67e00ab9a1d241a588f4065bacc3dcb1e6c2f2b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55b00abd8802aecc4b23cc387a7dc23fea69a5e500e66c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5df4b116451aaf9cab2ba5d435160fbbc9b58414fa4f3175;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfb6853c021a004014e7f25d3873f565271406354ed90a1bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ed67e8c7eb2278a45a1d49553deb950eece00f003518a2a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25c672b1e03c5ae9d11a85962a20862626c6ec5190758a97a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha172f1a3f71779e08f2c2cf81f3fecacf73cc0ca54100f43a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d0903db8cb58f165a823b52d5abd08148ca40c8a3b0647da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42bd11a3f4c459768c9d996ac75a7bf43861d61de6336d0b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65fafa75f03e9e534cce041d9673778fa00bcbdb2413b3b5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h853e9b4c5add988d6c4f777536024f4e3a510178e36e05a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50330a39204bda6270e6d81f5fb1248e8e58376f4c44d0ae7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78c83ade7187db4f9cd5f2ccefe64c7c9b663ad59811c0fdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h898776d1f9ad33b82cd1a4b50eb1fc7c6400aa0ac623a9400;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7621fd2f4e22d679256dc620c55c250b209dcbb364f4b98f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h931942e35b16fde14a983472d3634977b1a013f4a49fffc9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc395e902ff168e936df38f77007459ccb7fa65c2a7883d471;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed5683707852e2c60753315f756e25d6d83024bdaef347b15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79eb9997e2936db07b174f812eb4ad9a30e1adaed656068ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3997a5148b60908f738ff9d037ea4614208af54c64760aa1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c3f90d4afd9a79f736ca79f49b9240849f26a7e7c2f3b64f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbe5170253b654a1b2b41a62a441f0a8c3041b3eca9d52af0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4c814ea25d5c5040dee93f28af7289f4a30860ba5bb8e02f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7ab04f1d2afdeaa62b6042d13ec1d6e4a106471c983e0596;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca1c812d6a6cdf38a3634dfacc9bfc37b7bac2bf94001e2de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33681ce5b039f41e11a150c16ece87d24e4730f3171db766e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h148e8eb6156fb6db139b31830ff14de8f05fc67658b5bbd9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff9001380c5dbf78e861eb055b8bf3f979eba9c5d60c51f5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb84b09b614217f51e8e27e23732e1ad922a158742ff88f307;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd50e969b2ff5b954d6abc4ffeb2f4cb59014db2d635659c2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15005730889dba4c32653735467f061708dc28f020098fab8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56fb33c0d8970a5f049bda6fccbced47cd21c86c85af5bb94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac776fc8fb19f3ce80f4dec8b281abb01ec2feef9ed1a1627;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a2300cafd85a763129d705c5ed48d6ac0a9d6a9551140f06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf339d0204e0586157f09256e967bb944878a50a07a865426;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c93f91316ca55738fff44b340a7412b7c2d6dde7b5e757a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf75c21e0b51bcd2c55da87b19fd5411bb98d5898ca9cd96d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a1c40a32c022ef8af301122632428ac8597546cfb08dffe5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f0ab6b1a20eca6a2382a352eeffdbd5d9c90f57d1575759d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb508f577e3a1ceeb28c81e934dca6ac4c51672d525f44bd9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae399501add2596df4fdc6dada3b8635e654b0441f459bba8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45496bf3d601dfcb82b670ab2bf6cd8b43d7f138fc5e3a775;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h418f79c2b874a7dde0506788c545cd311122717d3f7f006ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5183dde9dc1906dcae6294a0a80436473153a0f0d2c1002ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b58261c7815d53cc648ab9e13e7911421cf19f8d5ce4473;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h684a46c627e5a53fb16c4540c349963b89b20c8ea32c85fbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d76f7e6678df34242a0a279e57ab97e74a4e8e667bf5b728;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea819c4c913ef894298f63d5c1604926cd51f88b82306b6de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63d95f17ae9b208916752be52f56193fab5ebf6fb2893b220;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dd8ba9ab69cfc6eed6fd65558be3af738762d00ad3b9e74b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd1299fa1b7da958567c786a203f94d6c56081205f21e5c25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf372b02374ed30ac916e962bd758f46a26490d0afe71cdbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c8c195cbdd9033a329e4ab8f17e7a126382085ee5457b014;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6faca3b458ba1e44a1ed6ca836c97f4012e52bbe2cf3ee7d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cb87aa29fe0c0ec7731bec9b412347479a8702c89774fc4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h429f7be12e99b75fe0ecdca9c2a950519a0e4793ef61ee5b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd47cc3b5b78b2a740cff473c300fc96b1701e079f2f02d5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha678a2bbfb1a054a053414721edf323de24b80543fb9de0cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f00f4edcc2d9035a383393c3cbb4fe4c2e71daa756e209e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h748731645061ab6d46c7bb20dbf1f1c31af5206ac699decc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde47c77f3c9b4ef4e104419fc1da5a06c2107fc7e304530c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dd5a481ce5d236a8aad6c4cbc497c75f944b6d56336d01f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ded8209cff6f3ee65c24662fd47081bb030dc322b5e400f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbadcf0a49f78aeec7b60010f3c10fa9ff664a354ecb3c7ae5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf034fa7c58f0e642f937f4c27f015b0d8ddefde55e054b86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95b32a332d77aa7321911833db008359f1b6fc903002e7910;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7415d60ecb6489dee388061ca0a512158060988f504591eb6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9771189c35e784a92260f7c102b150177e49ad7527fd8e2b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h465752dc5cc3a82debfb3cf75a3e0647e7619cb568ab46561;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3aa3bb96bc0c4b1b61640cef99d5e97fcde65b68e7476a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a40a7d7085721b423e347e7cc84a7d8f00789eb70453f990;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a33dd3bbbb373946c493baa42e1592f63f9dddee415b9c82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf842b0b74beeffb8f19f3d673236799db5cefc56d5c38abd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72d9eb77f874077591d784bd50ce8b9d09ee2f1623e7fda30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bccde254f4b7d7716143f5ea6b1aa3b9f660b1258e52b68a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45cab3c7387ca799837c8cf3f63a1ffbe5253c23eb042a7d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he025be36d2978c8ef17dbeafabca925f4a085d5d9beb96ac6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h281e5db43606a869610fce5a107a7e16b50dc952a9cd774e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb999a0edc904591965fb513ba6880417168fda8bd86c25f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9a5ff47ac785088c593074f7c3b638c8ccc89bd9cb470205;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72da934f40c0648c422e54af4d8eaf9cfa30c0259868dcf5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25ec543aff67712274a23bac4a8470869846266931b992653;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ee45a31b1d0d9fd8b1788325decb46b34c35ec4a5d79dd7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6d393b7089bb5726db07f09491dd8781b2185b962ef2fb65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbea64fa9bc733f56ec44212d7bf4a22dbd6bdf8ba5a9fcd46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6aad64047e3740dae824de69cc6eb6ab9255f3a20d6f30a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6584a997ad03a675c44b67a86986a691044fa4876cee2ff09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86a4f6016423d8812d194372c35bec74a33ba4d27b75a8e40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83f2421aa18814eb8b82f6f706d382845c1d1be655ba47577;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d047a2d1cd75dd1d4e73c15c37fd702f3fdfa3793e64be7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b36f0b5f510f8e02b6563bae4924b79f62889666eb85de43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6da9f8afc135b6aaaa03d922b22e7314794aeee520b675ede;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h589413e9715079b4894c0a37cb8335a5bf681df0cd271f383;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66a3a80716d0bc033c2083bb0744b228c04cd0c0a443fe479;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17d68a54498125b09a12e463b238d83cba8fa5e8ea4539386;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27db8ad5d437db2686a797cbe4c6972ca33ea3539716766;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd137f5bcd34178efb6fd01ac3ceef83a908766bf550722516;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6abead24da31e6b7200e912cccf3ba0210ee4f979679304e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2ba5dc172b017912a72f0043c0873214ce7a2fd39e20e000;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b23f555b8c5abd835dd03caf34af94b3db2089f7821839a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ba3977295f6fe32075c7229124d589daabe3012b7a55fae5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef0b3f0e926a66f90f06af5ffd1b61e7f87fbb17499047741;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf85058ed4587b136fdaf5beb2428cce659b886910d883a89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h579329abb612db8a1136f95cdc8cce6fdd5a6b0f809659b23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a0557b05af038ce46daec00a29679fa7b57d9c9f1769a438;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc748b60853aaa1e15cd5007c519d8489483cc5b674b16cf5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccc2020ff4a5e285257139e09af55024d53d818b6d7e30c75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2fd8755ad8c959a246194470369c30729fe0ea42fd0b7ca1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha875e58c908de06f1bb78fff9c43f38bdb0393a2f69bd022a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66d12068a5e9ffde479195205848083e9e00db3f9424b97ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7338c8a487b2075b7376955fb7ae8cd19ebc88d00f141cd7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa119fcec85dfcc99311a858c3134bd7d05cc29dc34dbc967;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a8469789e18f10cd68d6955848898ac11e7e559ff3fe8b96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5d76906f587e133a9080c5e93e87ae0f7f58e9fc632bc9d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha10cd087b05245ec35cb19bb0b8fbca9ee86bbd9401735b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf78e62aa627eb33f5c2c82fc3d8f4d1bbd4682b566c99979;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79014e66ac6678589f6265813c49f4ec630fcefb7622822f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4093d7f2a3b902fe8001ef9ba65bc187881111f61cd6d1e3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2eed0b0fc0bd4398470b671c83a46c2d66f30c204e5e9070;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc545aa7e7aea8f58f13d9f1eb5c085c74faac13978a9421fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha87316ff09e8d7af53df8fd76dd9bb7f60a0a60c4e6ed6a9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c3210cbd42b685221551a749400bfcebd1cf6be96c046ec7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea6246111d3f69c634fd14b49dba04685bb5a7fd1921d4dfe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5120b8a3f90e1f6fc349e9d8c2945bcb05ad453e758a28a86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4d16cb88343271289217d321c08dcf654fb2e5c8013339d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e9100d57f4ba019e13f1bb5be1d8d4e8cbbdcd5d5fc92a38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h669d156d5e09bbad3c18fd667fa1a4d92ae41c74c83189602;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb838e8588d0bc72a04a361fed691fea5bf049735f61f9f2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8850513fff8ba1bb700a4c384c6a2ce3c18e07790946882e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63a876480ba4381f07a098e3678ea3382c586489150561cfe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92b1c564ec7a7d8f64d3975504a98753c84aeeb052ca2de4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f41bb78eb5e5a99a0ae6ca66d29090bd9bd8ec4746aabf16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f5d0e49a23902e14997695cd00fcfa608af068d6aa910a43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h913a1d5d8d5a5c158d649df7125c29e93816f470e9c4ac635;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58cba9eb9e963a39e927e20927571b6753e0d503aea985cdc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he19406b24341b47adffc3055a6aa27855aca77dc135563426;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76bae8debbe93b52bb312c25bd9762cfacdc5bb023994cfc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2103e71fdebc70154021910a88531f8f4200b4934e0a9859;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31f5847e1baae4c5832d35774c52edf4c22b617961dbdb346;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd2477369890a81de5f3f9a2c2d42b72de409995fa86cea05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ecce0de5062de23e258fe80d8efd2fa608a9d9656c005757;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26a79cec1f69d5887d3b41cd7e4a6d05f32b87c83dbdee2a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h370b44504308deaefdd8e9b8b7f092e21a6e0748501e96a46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h495681f7f98801deae731b74a15e63066a4a34575e3ffee8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9768bdd36dd4993067b60f67e79a4a1ed93f7b23ecd208c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3774fa2bed82ecca15ca0b67cfaced13d16926b382eb24151;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9577dc441f1fa22e963342b2fda184a955932076b0f361c5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58ddee495238b409475489dcd26f68d67aa4afb987d6c0802;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87fe7aa133ae89911fdfffe36ea05e50127132ccf330eb089;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha54937f56c1cc9075c22f19c64dd97912f9fc078fd01fbc97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93de193c30d861dc436902d0eff92f1843de090cfecf1aba4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2cb371f1ead00a88f6a9108fc850a17b74de1c3fb74dc0ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74661b928011aba975971402209f3e461e423b39fa85266f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h749c9bef3d61d83004a3a7ae1c66a9ce90909977d6a897d02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59aab47298381d2f35de745bdad8fa9693cfdc029e3b51c91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4af9235c90bc93f93475ffc05bdb92c7090c8e6c60e1cf7e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a73bf7cf8ade120d49dfb02973f34eb2b9cf239747851a2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h900f83a277c583b20a7617c5789abda3981e42409f5412dcf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2231b1c73cd70f5004964ec05ddeb6d677213bf163236efad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71bb986834aeffa274a4f4461a13a003de6d4f34baadd9e18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed687fdb386b719c272b12bd0138ed0368c6e52e05767cfbc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdaf5b267096d16d0e306a2804c5807d1d0423fe141dbcf7bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5345debec15445e7e56917a1e620e91b33ee628f55dc0335c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf76b5342d23612dc9a393641b2951f96196684198a25b545d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9aadbdaef7976b36e2685e7b5dc4cebaf9394719ddf35763;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7142c067d14004c84ab4f497ba06dd7cb8c2f4aae1248b1a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf89fd18de0406d521592f0a8bcb317869ef3eb502940e39b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7802db8b5aaaf24179e49f00f01eb63c4ec33ae45d45097e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ab56e3cbea66086e018a7cbc716555af346e3679720e82e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49c2fd7ab87cf78a1d308fe63cb19223acf2b3e7862afc877;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a9cc366fa9290d47913cff068e2154157766ee26aebd95c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8587ed2df67d78b05ae4e6ebe5c47cc7c4954bc49b911e67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac43eb9758bb085adc9ea9bf42bbb7ddef0a54243bc878bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349d1297104fb8b9098b401c7cb6897e10563d4533fa33d5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8658744738cff7de651fd27f3303835cb94cabe98aac6ac1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdecef96b613a341c064fdc2f73548f3512c13549836007bd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69703ee5987cb8084727e02fb572690c155c62e4f4bfbd826;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a653ead3bc194a217064e2c5571d4fd092e2ee6f0f6d9244;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6e1e9ae581f431ce3827aeb71b54c5c646e667c7800d84c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d809a29719e5885e4d221538f5024a4445ec5422eff8d437;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf12db93ce460fd4cb3d174f3a61f0566ced27fa4a125e2c99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e9bc8e1c32da73349120a6cc1724079980249e9491fd612f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39807c5f14ddc1c42c93ddd3e3cf0c23931f88b8f51539b6d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37e374532dd0addc7f576f9ccea2953e357bc2b5d2754b72b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b9d28e6590e3d13801a8e89154767ce5504875ca2deb67fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6cbd7398a35e501d3af75817a3df0a9e446de9a753b7498b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h692613f7ff9cca013c71a4d544830b9df9015c6bd2683ee28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51d091a75764278746edada9a76991c2affd0a3cc6e11899f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d612923bc5ee9b366bc3585a19fc87e913593753ca3b68a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48be71ffae2c398f490400d7f0370cedaeabe284cec84b0ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f3e88ae8481c1202113bab9f2c34260e6ff839d795b7a657;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfdf2ad66ba02ab720992dea06c45897a12c8bb26e487f056;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe415f24f9dd06301c8897c149cde61caf743575c5ed52f19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e55ee6e54646495ee39b9a0fe9ff5d2650f6c04e5071520e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc28ad19873979f13e99022a40464af7e3f6a6489d2b8bd5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h862e84bc976257eaf1c337b3487071051a26c9a51036fb8ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hded12f796175d7a3eaa1329e885add522d9af749781b2ec3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43da98e767bbc2d02c675b67c99a76e73df6bec29f9859020;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d98bd0dd1b0f576d4d89178f06cd78d14e497a3696317dd3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58cbd436655b18cb78c9502c4fcb282e809bd8ec300790ee0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc13518ac6cf990ab7b24499ef18e2554a3ee7ed37f652e1ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47cf1866f01fc4d6f546a12278794855059b3496e89697ade;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a28630ad08f241d01568a1a6a2a2e074958ef458b321367f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bf704a67286812b3594cbb8a887fce0faa2bdde292aa5150;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h667bea1ef729b514833b39557055426e6e0a60d3559e06a12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6ab21247208860bd209584824a4dfec52b0fcca8642150c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h756f7880541ef487152243a1ab51151e95a616a75b6c3f2a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6ce677735a687d5db506843b3d43c3e0686aaad0aed9e48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a0d48a7bf3dbd1e57efcb04ad8851d409b25f81cef6b6b6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbb4d204e173657bb8226e0d7790b218f40d568637d9b69d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h730d0cc3070535b17fcd4f736e25a9d9868f57b06d6d92cc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb33806ddf7340de7c08252380d9d72e4df26d9796a7cef8e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e5764ce5893407d920139e682a318e5f57e1e14209f27084;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e4e197b60af0c0d84f977df2cf0e7af06303658c8a7ee517;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60b79d38e14591fa3f6e02667b05bc3b586a43be6e993629f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha196a5ee50d54dc74648b9cb25d595356aa5fc36f9e9032f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd437c495193c946d89d6e36f6f5518b0739bfe5951bbd86a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c5e495c7be2d02d2bd536395289ccbf291607619bfe56d5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53cf8e42539f2d175810352170d59f389f820b2d8ca769a33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc32b1e5b337a35bfe3ba45fb42ff6037fb1a8543309cbc3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1db6f827a404d58e80412ff063d2db6777cc18cc0e94968c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26bce67cf235316ad7294d05541fdc3f550bdb74860d15947;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3083e9b8fb0864b01b791d768f7e409ce14168edc1cf1fd64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc73441434863f32ab0ede61571076b1dd73ba50e9ed86e47d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a5b27d22a77699925be7e2af30904b70137d0e055e1b8bb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7515ffd08de91b8933c086e9552bfb01bfe042ae9b7c1c00d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9220303c4ae2cf5f8529efe12174ebe190958d2fa789d2130;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h589896b497756659d2fdd0cbfcee3b839a9f5d223155d30f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b0969734a326f8ddb4d8bd92f57b395160571b435b6f3577;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e19697559d9698041bed173f43bcc2408e669f0c06e21db3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb688fcd2d5544988560b00d854a3c5e34c09cbd0084d65568;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8928db37e095dc28d022f4abf25cdfe89e1d41af0f772b49c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd40d65036e95ea9d23a7e2f8a10e9e591c14511e4d7c4cf3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h332fea5977772378e48d27fd4d9c6228d120d737df1eb54eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43200742b4e545b82252b7a4f201bd9091baccced00137b29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9bb7a2ca99f9f36a90ac84568c6bca3e626b39429308f193;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c056fed5f7df2004191445f289fa0c3ee595d161ba66b931;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b659e9e2d3aee23be03e51c2a32c94dd060df8d84f9072ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1fe532f4c8a0e2819744e7bddda7f43b6f17c55ad16b4796;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf76d5274d0879689ef307eab7b0b3f6e085ef1d98fcaff157;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1a8065d3bce3d6e9c0a01e46cabea73974148faf158c1925;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf2c675503018ea8fba90df09d7b0d4ce6d9418fccfda0a9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ed4e1a69b5f378a20164a35daa0834c1c34dd44cf093b8a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha649010529fe5ba7c5e27a243591786a327510e3821f0f95c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8da945aeb5e43554218e4193c8f0d6a3186750faac8657e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45b8b95ce9c0d6477dafca9283a0177471299aa5e48bfe4b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5972077a4ebc47d2573adbb3703fde953324671f207f4e9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c5791473f3ebaa4da7a1c5e6e60f283a9d32669980ff594;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h708e9ce0c8e83f6a5c96158246a719636d6e2cd37a76d5797;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32e0b037c5c2df7b4b379fe3d77bba689ff135b9a6973fcda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha56faca62a4b84bfc7cbfe8ddb3ff1370b127f7eb46d622c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69b61cd8c6aecd9bb54d518960cadd68e686202e63e0b877a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h717def5258323ea6bb221e107884c392f3f3b4201e4c9907;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20810a50df03b0b7d2fe6c9057463758f4369cb737153eff5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h827ca09b7030d04eb2f622149c5f7c7c2b9126668e264dfd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd878b91f11d2dd31f736772f9f3681871218c3b7d5a218782;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haad78f72a72fdfb734185ba024c21cde0f358843fc7e6d527;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88a75e2338aab76174070f4eba3504aff73e358160f782ba5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5bbad9bcb72fb1a9926884ab20ba611ecb5ae66e98052826a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha03f6382f748436616152b5336727bc3261925474a57ca0dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f17e6936757ddd874f45bb3472e2691204b13b7667cce6cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f57058d890e5385d647569d82501128bf96139b9c154cf19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6591dc90206ce0220f83dfe2c2d98a288fbbd00a9f395889;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a1acb67b34c5737639a444e7ddb92ee7a657d1e44abe2ff7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8221244d4458057c1c7805a549ce64f7a0f703f4b90379f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he740ccda6f30ca4be9753e487f25388849112a5c7e11dfc56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a20857a234331b5141ec05908152d71a1f00ae346087a85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h830e84b82abf5495fbf165e2eab0ee50a9aba0e993f402a95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86813010d72c1a12c0017a9dce11da797238837a82859f3a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70c0b793f907d9ff386a0c0f2b71c350a470a722ebe7df1c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc02bc9ffebcc9923fbbf4bc59da398765c1e652e5d4af508;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6858b109311de2adbd2a8e3295da751bbcfb4a5ab3fe24d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fbf6b4337d6f0de9319f9db2a354a56e9081c687b6da525c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dc441dbb0a36ded5e6ba28c32eb0ab93b388108e45a6d5f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0db31182fad626ce9915296897504cb75dd0968c9cba89d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h282f7e943f8d9070e6ac196846ad995dd6e284705d365c02e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf055da10aaff68deb7e4ef01a9e0da72eb54567865203078a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9c20387c9edc76b0ee8d3b6f525f4a39364b1ff6c698f47f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42d1b6156c8801840505fd81759958acdd2006e7ed25b5a7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4662738fc8db358c469dd40563515b839bd98ed824bce2cea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11735bf990d2807eda62bcd7e5e705b946a933727f570dd37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19f1553d9089ad103d269641496f687280a627d32250fcd9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bdfefbcd84b863a5f904f83932ffb6f308eb2c5db1b226f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c6e5ee8a607abc00ae27aab94e9ab988e3f352732d2e0af7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h303673089d24f840c273052f8bfc5f783a9313104ccde44e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc78b0b28f5b40bc59eba99e3aec077834686b1f3f7add2902;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4611585ea1455ff5f90ebda6fedd8439246a61b354454346b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76a84cb172cd3e2669b6edfcf2f0b831ca911b8917fb68d30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h395a82185339d312ff5de87561b9cf66ca5e1b90f0157cdb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14d6ca755081d2d996789ab7292bfb62daf78ffd5b20061a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d66ae743a8be144196e806731a1c469d317f20453c2ca45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h753ea27dd7f3fe7a27399315e00bf8cf4916cf330d58f7fdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h976ea88dafa2fe5314fc3e911267ddad4d98915fa75489b50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf737929d1653a93c6cf1c3fb85f41feb7178ae830601db967;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e20192b5c7a11b6f9bfb8dcd5fafab417db4c93780242a14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f903cbad8159250dcc454b027a161256781d72b7ab52e32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha054ea87495a8a6347a7d65120c9f3b26c08958ab3e2d4644;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f2e4d8f843e6692ec9313668a9e01d9879dc43a7c3144db2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ef757a8506a2460b199ba88b2ed243cc44bad0ba3969dae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a18a05d84f7bedefbd7ce8630389707824ea470dff2eaaa8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h512d4579a3fafcdea794079880d44c6b947e560529ee924f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38d927cd02c407e5207aa0051dd6761dfcc04011a1e68d325;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb83e6a768cd5ec4672b3c0df0e7f0ceb7b2eceb1c70fc66b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60956c286657d150d20bd8705205ef14c4b8f36df30e8940e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3898d60e9860af36ccf7d78c2eb932a11003f2a041f3826c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1e1d9c25f0699d8fa996f50009b200116b9896a5a30f0d0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41d02d9a14ac3c520224bed09d84f4476c1e40306abb37072;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bd3cace1b258b933da07882d97388bd8477599600ac8c83c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e44e925b2246913fae6eb1b5fdf8cb3f79438557154ce6a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74142ce5834156b123a78f8b9849fcf3a217fa3f8fd3a7265;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he63fe926e6706a38e789462d8c30583eaf15a0a3285010fac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb564290d4e279a2eb7d91c0207302b65b47f0c1933d8a24eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43d3cd5658fa365515e1f48686d193226d0059f6a3c5c6027;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5efe8c4d6966f475bd60a1e1e693b836d6e0c90425b90768;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58f2cbe89bdeef7636342905785f6877084a820d98caf9fac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f18795506572ddaeff127be23aa32241a1216f3660d73981;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd04b7645d57efbb8bbc85d136c39a77e86074b630f3e72708;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha82785adb10792e3093da5d421dae44e03bb09311803b0bc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79fc3b3502779450e556a9284dcdcdfa52dc9e0158a9e015f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65e6922f0da41ed694290c4747a5b70dbb9af223f8ca1abff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54f743cf49653ef7e651d08a0d8fbab5fd0796678e9db3f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d191c8024684e6f5cf081dfe1822d28fd6819b2643bed4b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb85c760923e47711d09dca03b521b05a41218f942e29ec2d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bd5e1e1e9660177cf284506309791c2dfe303f0f7469cc30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2356317d79d048e617dee3011d64663c1428bd57a817be486;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7ad477b01e35520ec0c48c28a0ce012bfb5d24f9a398d070;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41486612790cd2bd0dc3fe4152e45d21f034e041d30bbb098;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6c842493e5e5c5343ad06951780d715841f015a23ffd2cc9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63b7675d34ab65ee78841571c4b00b4e0da0230ca1d9e1436;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb34f793c82001e5e760663da2accef033f2d74f6a1482fcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81f58015703450413df61de4c859361ebc51648723cc70419;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h426ebd1e8c3c97be242c318d32ae570a146b6f359ad972789;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1920b76163b8430af34edb551615454ca03183054f584b372;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h740079fc20697764e50c00c1d3b1d16ed9d82594bb51e094;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h942aceb447c80b7d6652a9c98aae28648f017e43cb3bec25b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha65f5f3bcff276e401c03daa4833b148998cc20225a728094;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4640ec724ea62176e0208a42dc6ef5600643490eac7a74b7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c1419f565db9d466628d2122b31042caa2addf41097c00e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he69feef8e3f3cef3b219131afb49529912675481b51ab4892;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha86365219c745272e868b216553dd4d3ff0734aee191fb055;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3ae062ad1bd80005ed6fa86f4a77e6921bdd111dfd756c0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h101809b0ea38d39dd96f867579887ff0432079cbf5027ff06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f576c5806b48aa64214d415b83e049f19c931b42fe6b659b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6f265dfed7fb91a46de4c050c194a0a28cdff57a0f2ee27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fd4b9d921aff499578c7d586ea7cfa88b5c7dc2cb7d88705;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c75b0cd34ca8fb514ab02eb9388b2d70e4627d50383d9b9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7314d8c3a458227a4f6996f8414115d7663da959d7a3243b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa3985ed42f95ad86ba96047e2185d5b22c913a8707ce325a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h584421cd6af878ef925320f1f2abcfeecc2f81bccfdbf1665;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83a4dda902c363c71be8ddc5802140b994cb6cdc50b45f350;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h352f115069cb3b1dd1372a793780068ad9ca796bc64f9f6bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f8b696724ca86b0fe2d55384f026c47b96a63ef8a76476e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73bf23f6a65bff3751e7b4de36c924e29973538f4256c1ee6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3022891ad67b634da93b763ef4a30da76f69debf14901f82f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h547f8cda37f750de31a7f6c110a6afd0cfc57dca273daf760;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc012693bcfca13e27809e8a0a7ae6bce5daa720a28e218ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6a11f875675a41c53ead5281a294e4a35f258af3f95b9931;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1010274fdbeaedec4d68b0a5eb123fa54070ff99bc89d909b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f6bb26bcba9ce73d2d2ef1448e8d2e81fd3f223a1bca54d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1697236baa51dfaff029d44c04281896d08eb8ed224822ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3eb4c3f5f23d402a520b58714975d5d5526867b2d6329f55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7b6b7bc66b4d12c7e5037813646e95fc63d98454fa7e06e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35841a2022d7f28e0d46205558ee5c6523f9d9102be8c626c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12f98e4c7734d4777cb1d239f9386436033f31a62e527120;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7432309c4f7b9e7f29aa679530740ecf0bb9138c9c37c1cb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d59cd0de76fe7cc4c759cfa812bce8a2e089ea4cf35c55d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he92f649b2eafca400b9a53ebed62ad5b93e352291f1ba7132;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h800af8d9a5db13e32303246b39c7ccf25fa3ad6db24b5b1b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe09921bc969f5e3f25a52f9d306a733a086b4b5649acfa27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2027a7111eaf2d812f1e36bf65fc8b62da987e998f6596554;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h847c40502441d1520adbfc4d1138c6f43ea5733e06ec5a108;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90fc79be461fe62d266dc2cfe51d8db15afd354e87f6bf91e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd02aefa1aac77e777207f3a72b28889690fb9c4a36e146890;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16367704c310abc55c42e915a9807d440a03eb2710b74f9fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69231f15088f42dc375bdbe921e10afc0a907be46c8d108ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6fad0fd793831368e3f84c4c611d677add95d3edd9cc29b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b2a7d7cdf9188d11a4c51ee2e49a729e32d13ac22637e6e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95275bbe90200075ed259b3296ac2bcddee7a4fa25d7d936c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6587283074ab957b969757f1051d53146c0ed688ce3a5271f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c5418581dd265e4e83f435df564f9863cd0d9123bbc476f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb11e503eccffdcb18d22cd6fa38f8e03e25c612ef187e8c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacee416552f2eb2760d83e303c864d8e4c376b73c52c114e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha73a3799749b7d099d7b86a1d81248d17fce0db6204c16b92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52cac6cb6ebe3c8b133847721dab4ed64517c44e2fcc79e4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8cf8ad60a77c0968bd7a24328d18cbe4dd092c2283955ef7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84fdc1a9cfb15e4c08f7b3701799aabe7b783ed4495e78af8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd69a7de72f6bb5f4e3b0c9c375cea9762b7faa41902775662;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8482c7b31dc846639a00afee7be57448947fc28ecedd38058;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf854dd9834f6431a25fafa2d8ff4979112abad9cc522a0c70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd641fdf3e5fb58976d84d0d83130347b5ab8506813a36b69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h734d09456c3e014b1afdd7051f8f55135dff0b813e6ff4f69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59ae36a958a5c78297e5e10d0de4eae85c3b6b4ea9edfcff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haaf684fd523a846aff2cf3fe018abd9bca6142e1eb754587b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89a6c85a4c0af1f023fae58182281d0a64efb5068e34c4026;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf8ca22f85b3bd9fb135532d103525c5970771ce226bbb893;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd817f9b0310d1bdfad3e742dfaa236d9551a683fb7e256b49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d6240c70c76a1f9fbd3f16b5a6b1dbd12b8d00575aa0911;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a5109362a8236fe7db3c9b2295ca68a699ed7a693356f562;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3c149aecc8bf0d8bbcb81c0b171cff2b0020854927ef6865;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fd0f06850860050982bf1dc2c0aba984f6b55d9485a03e6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafaee7d396d0f5992447e2eb783c4b0daa8841fceeaaafbe3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62ce9de4071362ca46b27c39f1167702abea99b20a608b40c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1fa436e6f50187ee996a59bb5d890ade1e897f5781471d6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4925be2a894f14dedb9f26c700ddcd098d6e7701027d9b08b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48fc3bca25702315d4fcf1382ed6103f8bdf673708c6c9505;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5163d572f6c5669addd06885da70bc3702b78c5a2f5bb67d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2eecfbc643cfb588e4135956e8f990892a314703f844c6457;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb7c3c14278b18de8b21b82c7e3863138c6a9ffd41aafee4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e5edab4e078ae78fd50aecddce6dae06b654ba7aacb543ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58deb6075d420f03f5c2a14cd7a20c1c6c15a6b0a441fe9a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11d10c93747bb6b5c669139dfb8a0568fde9005ad53d4cec1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73acef26d710ae8d26e6a530c93059023fa8f76b5aaf070bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82fb08db8a332ff6cc6f306443403acb9dfcdd8aea586b943;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35ad90c27ec66add09e5cbd88b0fc498d2c9650c5cca5d540;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h736201562ba41273c43e931b8e682b3359025706a36610807;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34d18e5e771f3d53af7e6745417c4349a7819e855ff145d59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha92f695f93863ef2264c2a2c8105e451cea06adf11de4c16a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3a020b8ccdbed00dbf397726517fe959e2dabe83a3657d64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5243ae9f32eae06b0f0883aeab40c67a6fe970cc04690c8c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21a671761845711137191951364f4c04f8c2dbf8a09e47c02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29771ad0b6194d79cf621def0a40421c3fe871414a1b18d3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4048e018a54d2455b646dcbeed3929ff365c716a2bb763416;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc99921156c9eb7f7e47b4de406eb51cff24d2859916c0042b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h646808e08746210ff5010331f21af7974b946daf577abc375;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0650e214fdcb91b17baa3d4627286df4f5df219288e0e90b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c423f3a42b3c67fbb52de130ef831df522bfa07476e7530a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde688f56804300669fa1b67100d0ee00c53d39bf2e2dbbd2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7690ee555064cee6d5a9707a321d6deaee03e6352ae657dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ba6726ab0dd5cae795251afc4b3eec7cb2e59ca0950b0f87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1eeabbf08eb4486d003d1929349f0623231e632fe63c2255;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35b9c77a3a597c29234b38cb25583f00ed6d0ec648d5058af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1443c161729dad37062401fa8479c294871c4192a00abdc0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6f4d6ce0cc4da3f2ecece6ececaadcf9f6a237cccf42b1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55fad95531dce73c96b20ad6e70f5075dc4559e03a73f7825;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdaf27d2939dc5fa3f3c883f376c03d5891005d1768a47ffba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84333390f40430320d3a6a9db77bd2482fe1daf32241e709b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e700ae66601761f82958cce730f3c07d41d589c07ac8dc69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5513434268459769f7e039af0bf4fc80d8060710a52e0c07e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9656ebd4f2178ec8159feb5ebb758d9ab8a785f460e350554;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59ddc58b9568ecfddcf714f6a2cb50a451d44fb3afe53067c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12e8c4493409f7265bb316bf85d75ca5e50e7101016d17e38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h350548344dfa4ca4428a8979096dbde86047cad7285a862df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc87ea16bf2eb6897820574934f397ba7ee3f2e970a9367b1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2166e0930040499877ee01621cdb28c07f31bc86b0f99e40a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc25e4b55c7f91812ff8f09aec1e3b3cdc9682d0fbc36b906;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb74fb257658ce72624260545d0c8264514c1408919fa58044;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf472dedde8729b9201c1079f1fb6f8e87988bc6f59b681dff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b3be7760729d4bd8a03667d78aa522a6547ac9da3d75a8b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ae187e130a4d2ce9118f048d87770f65a72bc4403150817;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a05e2bf633f143078c5c0a54107c3ed0dfa039d7aeb61e7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb912ed06ff67af9e1bdded0735f891d317febcad8475bed99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40e707aa167b7bb1a208fb73bdc5db5e1dddf0e4997e39023;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61df6b9482841381b31ecf32b6f297af93e3309dd08ef91f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2669ba20275c9794719779d47f5c3afbbcd2b5d1f5e5225bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had26c00a12e92ac6e1ec95148152bd8be1b0e5e06565a6244;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bf5b7547377f606df2d87ceafa9ce4a7abfce4be2edf2e5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b1a340d08f12ede2300e3dadca6e361a0157fef1a29fd02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h206f61606507a89019a9a60e441160fd781f0320ed93e05b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf93754e674e3fdfebe447f19afe6d5abab6074ee35799ea5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65816c39a82e6e97578f36fcb4d58f634193fb1b0997625a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h190d1c30705ccbcbaa62a30e0dfa5d5ee3cbf211dcd1c0496;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a6d3240c8a6c2328b7dea95f8e54574c2a726022d9c496dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecae8ee5e5b20a3581315579a9602f165d982ddcd4eb7cc8e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12612952b2a9dcde78027b9daf791e2679d8bc17813df1abe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebbf09cebb90fc851d2a285018b11bea7b4261ebbfb0162c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3cc21bd955c10a7ec8bcb8f79d08aac3f85beede25a85b34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92a5de1a2cd02f70a06f713cb025b977905c4ba43a0e97d01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcf0796e30c05650cee282c557bfcf3da10ac9d4553e07910;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ccaeda8b377aa4817dc505a9e457fa288b2732efbf65a48d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3940955f14714d035761423d41eb300af2d70f71aab34efd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he990a9b7296fb37b875eb675cf005c098b25f7cea97f63b28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76acc9567dc35f78b9faacf3f130696d35e3cc7838106d28f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h328258118c990c51a88b09cb5611da4c5448e94a442ad8dc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6af46d1cf5abe835e749a530597ea98a5efb7ec944cff37e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h245fae08e5378338bc4e12c3808fed57bc48851ee96283454;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27b98d8a2a482efe3935214009e3eabbd0139b262ab2f810d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1dbfa2e449a1115933a7a1edb09daea79aa0855aaf9fd070;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde087aeba2e64f6ce197122ccc949d768df9dfb0777f4a4a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba86f9799a8e1b67fa5f3d87b0b252cf375c9478040228dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcc6199d58075eee3b23776add2361d1453e6020074b56347;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ac1d98dea6e05f929536b9307af885ce214d2dc8943ba714;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd559987bf6c247ff2cce0366263403a43042e12a62ae7092;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8791959039c40a5d2e9b5e4ca916497a649a9e954df213a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb65f46ee190d0106872ec79de72e8af8a0ff350a74327aa8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he64b71d6c3b26ea7dbbf0a77e29c15d341ca30d71fb2ff4d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14918a8c801fc663c28bb228573c71170a2318525e2f87c53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he614d4040c7088412fd2df28d46597406fa580808e9016df0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc8943ed45530bb2a33f8b002dee321fd7b4962408a62b07a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cae81572a33205c5f3e656b7ab5643ede0bbbe66ac24c2bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1271d2fccc58e2bbf10e69fa6882159c6257eb8417d1da9c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc461b31bfc3ac7cfa7a5debb5334429ba5f50f30a174df97d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf758263704d8ebcb2f2debee470a0fd473e582d181ff6633d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e1c0d354f7b600cae94c3b8bd70e02c72adb52f9bbad3a39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8964e8bf62e66917f616c0e236ef372c19193715848b0e28c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h950a9525bb8258f6b47ab767a2784de87e644e1acf9c3bf30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72b674b19e765850a61f4c686a92305ed0b0849c96418f788;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b6261647e13c988bd4629de2458a395d97a04c75632e1eaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f8a12fcbc94b2c69d150a2934c67aa5d233a3d5337b467e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h951113753bd1c2a38b0d31f197a4c7b5e3a237e9cad72413d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78a7ab5ebfd788a5d69400fbd8954af246bb67910057a8c73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd79e009f104c3df965ad02586e408a3b467e699ebd805435e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf512447f449aa3e394fa738584b556955fc677f367a70d25;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc496e3d92490c61cbef7dfe681b4e41c51053c8dd5e170417;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3eb6e805c28c7babcc847d3d36550cf32fce1f61e112985c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h425b5172de1f185c38ad9921b60bc4a4043910f4e5ebad843;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11a62530a56f8186234a94dcc7b380b0f93ada2c0f7101d2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89665485a0853ce74a81c499940dbfd32d4a3a9bd1b9c4041;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf05ec77bc0ee48757bb9c4fba484ecb262337586819fa386;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb25746e3d48ef20c99edbf09a811f84631c0702526a5d77ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0e728a308f09d2eab7a96c06ba605a716acb0c561add6077;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h578cc452debfa3b393c3baea0c7ec07e943025cd5964e21dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda541a02cfed2f45f8d2ccffa59917964fe4999945c25d2eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55b98edcf46cafc9a455207974ef5f06d692bfd793f4000e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd88465ff15ea61d2b9d973312860aab37bff86c10260e7645;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35975116e4f69f9951c8d9d9dde92d0399b07d4791c7e94f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4562bb5c78b39c30a87e25587ce9e60797aa8df530d437b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1f1bb7d758b64b7eecdf6f3c576852d6e72798e46641b6c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16de3168e576362387cfb3f29b887378165dbe92880778d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee43d138ee7a0df0a51f9db6468667bc8dc4df8fe894ac05b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcba36b5facf526049696be46d4d8f4bda50ccfb84ac49c327;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ae6965255644fe1d97f986366ba0af92bee44982e719e264;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc94ffe334a581d6d5a0fc162364bc4c730767dfec61faa35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d6ac26d69600f8532576f23487a767513f39d75f2f2de130;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3dcbaedcc25067d9bbef488d2302d52fec7ad8ae24cbbc625;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58870229b367a825003f784823243965660c72413cff7bff1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4379a76f7caa0181088baca9bd5f2c6192717c2236a30e69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16a7a36c324e9302bbdcc9602e89c4317df3dc9b57dbbd220;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6031569f1c124b5c95102adb49f05e43c38efa076381ab03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5be9845977bb80a8add5ad7c5e93f2a5c8e1b5d22d157fb5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1efd9b77a6605c1ded1ed775dd193552c1dde39d4ee227962;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0e9c0c55c7da6c1ec308b3b91adb57366dd692ddbdbb3902;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c49ff72f5fbcbf3fdc50cb66de1b37d514792eff5831db4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c0ecce8bd369907601b5ec7a37695723dd66f6d93a7242b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e8ecd04b6be46b5a6abd960a629fe7a84c1e53d1bc3b8fbe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69031889375c0cec2d51dac61fb5a8ce1b8aff0ecb5fb51bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43e64ef9a923bad9eeac33ca9aa1aafb275b87c32f17234c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92920d1f954f3f36c98e37861651cfff8ca41c104790d69e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h230b00a08e71ad3dfe16315dd78d4403b723c1db05bad8c96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8bb25a60ec0f74d51088b7b5dfc665dace2bbd3fb1da4611;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he63d7aeff64131bf853b6dd5e2125b8b6ece57c18ee690b60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4925a63859885fb2635ae37fb03684f24f76e71f8e31d7ce2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63b3ac2042687f2c836e8f2890fcb2d8b255568b8d54141fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4fc86b94633de1e3d87a9c6cde7e3576dd6ca5e389934c23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe6b3e5b5bc183c7e8a3af60c36765836b82d7e24ee65a02b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31c2620daf49e143a435fbc993978986a696f3a9adda60fb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b18a30ba7b29f7a778d5cdc2fea22bf508f00e3b785e460f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3eca4922855d19d9ae5cd7bd7b525f740008869e5b10233f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5707866db454ae1f784971439cb44936008f3189473ae3a10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98878acc0e32655f7fce47066df5eac33fab9e1fdfeca69cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39d0892c0a33681f335bd0fc21ebff39137756499b5f89b0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f223d8f569200f98e4b38d12ec19d6fcde87169a78f717d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57a7a31adf37ad9118e0bd8f37fb2b5e1d967d286d4f90b64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h135f45aa52ea1f3fc716b91502d71296f6301a9128db1b509;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf328941a84557c9aa2dcc111d8eb7e4b78c9292c9037f325a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7039cb8c87dafe06459590d2d43fe4a0fa69edf1e67d35bf4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e7d7e95af8af2397d84a0f8269e979891bab94e8ba6a609b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d0fbd8ec6fa030a46791045c3d5ddce35ea311d4ea8c8a41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf04b71f4fd4636821e073ae31f5f1724211d1b134cb62f6ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea9e7fc39f2dd4da1d10adf36c74aec2a18b1c36af1a60ef8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0990155912b3a8805b45b67ee5fd98fa8fd4a52ff3a67915;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f36e5fac913d8e2751631cba39da2c718470e139423999e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f868f808c384450fd5e4cc79e49b0293441176d7f69d5c29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e49e404ab62f1ce402bfd8a13fa7363b1b2bdac66639cf09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9be080e7adb74a74fa354a4cf3e1a34c89be8ead4b3e5123b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84e83e0a8541526ab87adb49baf6c39b5149970c1044bb2d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fe24084716d11839c85e75b6a54be84e6e15d833da5001f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3dc11472def0801df7538c7396b63666b45b1342c3a66293;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb7233c8d432abc38789abebd33ce55c4db4d06bb28233672;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66a67398785e38523dbf486871c4a7d3a9b8a7ab86ad4788e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1bfddb7ef60ca57f3f3a01b8867bc3684bff3ec0f873372a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7661351d9e930771b63ed7aa61e3128d905d69d12f82cff5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bff85bab7c0172446cee3403cc1f7627609ad919eb2c7e5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5565afd7417c9bca80f78a064cb37a15dd9a065af5973a43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6c498aec09ce5538da82aa070fc89afc3508686359a8bcb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87d3891746def0eec3addb348525a91be1a28dd1137071238;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h270974660059b59fe44ba693efc91bd9410c819ebcfa46f45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68541e7a662f39b9263f1aa9f1494c9919a01e25633bb5c01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6effe07a063016c206997c1b1948bcadd54368439d769af80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c988ba18dc7b9c211b0d22ab6f62d75757b735e01a203e2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98d8769102cf320f5d7d184231b5f3bc5a1e0d6f8d6287d5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5d9fc2884d9fe2d5b11af2fb656ad41c38c5a4cb8e05173;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87ac049121c21ac5363e1a8b568d805af121b59c79d97be97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha48418e9c5fc7f5af8307c1cd95771f1ab15dc9f53f490154;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ad6a662faa11aa3230e5faf180ad44a41e2a388f14b52e74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bfe50f73ecfef4012ad77df26bafaab5b4c67d71b0530af4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5b68860848fcf6743bb0d8b18c1158dea49b47da3049f1c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dcc179b74a9c87e54d26d0a4a98408fbb75fd5004734c91c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0b5f05f824f67c9ac76f8b0f9059f947651f2e49f3bcfbfc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8a6696f7a893dfd3cc9d950cdecc32511f7d70daf15c9fb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0f6215ffd9a52837061b46950e3cbfe5374ab206d65c635e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ea59fca851a190cc9e3e812e1ca43d3a71567f083c36a33e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac602dce4c42b9f04840def26835dac7b86d601c44f60454a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80e85281689c48c7b8623f2434f2de5dcc190806ee0ee150a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h687c9558d0772e28b479e0aca5a956fc171fd77799bb89210;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h685259a7034039b631e747254f3c9bee1801f5159b33403a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbbb3ec8d24095ddaf76e1b6a7422363e29a3400e13d60da5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2fc6dfa4362195a503219a742b1d73e56334aa085e2e91cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1ca14e7116b7737beb52c5dc8ff1acba5e3d2896d099ea5d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd737c396c673edd47e82b3fd82750c97ef181ae084908e57c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb16958e03406f41d82c6cf41e848f5c0ba67640ab63ebb17b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc592c1135a85f5961ab800347695c881ec7932d384c98c98c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8550814dc14d14a92d40ed4c450c0f628d4ca5ffb4f24d54f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36da253c5d889ad7cfe73cb4b67677fea361de116f4f4d0de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49d5b30ae0215fe931bf1a73a2f2a832eef58edca223e6bcf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e1cff5e1f5bc09eecdc363b77454699460c96d4278bb6814;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3630598e0747d774d278b455a6f5bf9f495414629fd27f958;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fb36eaf4f3e23fd8309ebc158ec6c00f4ba627209cc4d93b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h526404869b0f5b8e5ea4b87eeb7a3991f5319bd43d99bd461;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hface2c8becbbab159dc0be7ce2facef4cf125f1075cedc5f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78d2d2a14482280eab19b94e2ec2c586e7ca208b9eb2c69de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb547eee61b64cacfed56bf727a8842f1ae4bbb70643719bf5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce2f138a0e73acd3a7df52b6d0a7677c2ce04cc4f19eaacae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39db149a89cb9ddc7de4661b34010c37cc120f9b11ab91043;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb4c59b948bd00a2a1aea861358ef4ef18a2ffe1338ef126;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h212bb387fa7581c9049edc0de041943e22670aa24ddc025ea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4916eed639f066cbd2036417e734c7fbd8e64a4db9486bd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4178bd50eb095740fff92e19433c1bf3cd064d20b5271cc21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4273454fb7989bb2de02c40544802ea52da6844d1d50e224e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ca6c375e2e79aaebac0f62bec3223c2c1aa7dc0fec64f0b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4680544556b705684bc935e86d25cdf7a008ea85e78e9700;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd490b6536bfcd929799d34d6245f7ee09c6a659fea559377;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b2b8fd9afdff10ced3db752ce635437fc84b106448923b78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h412b7480fb3503ed357e21c1b28b3ec97922533f0a27ed233;
        #1
        $finish();
    end
endmodule
