module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [18:0] src20;
    reg [17:0] src21;
    reg [16:0] src22;
    reg [15:0] src23;
    reg [14:0] src24;
    reg [13:0] src25;
    reg [12:0] src26;
    reg [11:0] src27;
    reg [10:0] src28;
    reg [9:0] src29;
    reg [8:0] src30;
    reg [7:0] src31;
    reg [6:0] src32;
    reg [5:0] src33;
    reg [4:0] src34;
    reg [3:0] src35;
    reg [2:0] src36;
    reg [1:0] src37;
    reg [0:0] src38;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3])<<35) + ((src36[0] + src36[1] + src36[2])<<36) + ((src37[0] + src37[1])<<37) + ((src38[0])<<38);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ffe137fcdcf465b23fcee8283425c9f492053a2da769867f4787ce071cd220be0b004b5733d9ab7364a4d51833c13a2d948;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b081fa5c869f8412676ef6b9b55e08a98968be32386b884ce956f384553a47b5b0e493335cf658ad2eb20d0a769ffcfcd17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4355e4564e506f78ec780811df76dcf5a3023e5c9f6c1c4056620756d5d7c73057ecce871082e374047dbbe89274b8d89eed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b3e44d606d6fffb58edaa578d12186f4317273a829ac0d00d147ef226e2f01e74e491e2e3fb0d7be39cbbd4385c97578212;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2770cbd039eaa1e5fae91b3267a52e13d3582f8de59b3d8d9b273318708feb48944d18c647e9db3726ed5f5f0c869267752;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9c31fda3ce3c065e77e24bc3580c7c5221e1e211914012ca105abbfb85950e1038dc40740ce9f9b4cfd929c9382bd78cf49;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha11876eecd30eef6ff3f090c0fca33c8b51a14a9324f5434ebed196e889309bae528419cb32514628c0bbaf8c267e9a44966;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45742873b24fb000c7b31db095bbb75e487f9f77da1bd1e6d5645e1a5fc411fdb5ed4e776d8a63700669906fceb049c430e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h126f01db6df393a47251519aa2b468a6cbf5b0680bfb239308edff48b96d0789ddaa06c8fc2e33d8829c86fb674903e1ff22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2500261aaa8ddaab6eb63926de1fe8c806893ba9d1d8311485c07fcf370a96e0228272cea104ea21b6c3802fd4ec1ff2c934;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb635cd1b793f4891168363a8c4c68e24040dcfe5073654a230d02b9f29c47a5ce471005d7bd0c4bbc520c9f3bf2ea233dbeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18822ed3fd41e9ce073c594d3bf837b6c8c26f1e094e6fa4558a1a2742318c64a69db2a6814b8907e231f1b519b5db82c854;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68b2675eb4f02c5eee636cc13c56a55c42f008396f3a5bdb458b42699798495ae2a5f2451687a389a3e033c24b4a5ea8b54f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8a42da70b6f04781c3af331ed51b2e41ad0a1fc33f9181917f45079425dde03edcfd184ae0e137be4548e37b65949777c54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc92dc0337093997e44a80c392bfddde56995284a8f699734eaf964d372beb8e08c3d9300d263f5aa6fe97bd2e71ff086173;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23ef54e8cdf815372e5cbd6ea18b4b6849ae68bbe3ec22bd21645d5fc48bc083bb093a1b7c8cf91393b84f3d0107ecbe8d38;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a56b8a59659940457a529a6690176df4ff2df54606f7615349e0fea4b1439005c6090082200a7594f08f893802f67d242b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea254b9320bfae6bdab1e92db2a7e13c902633d8e3ffb6999d146dc0a62b0644e2b8987bf683032f85ca3d77717d9614ca6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb24b53981fa992ca95084b3c1af8ee78cad1ca936c45e9f6a3f34c096270832e070952cb91f238eed6613af01c4ca15c0366;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a67289119c4f0752bfdc6ef006d7f5e7d5c67ee32ad5e3ae2bae44d2546eb7afe7368b8a5caa7cd795404717bb71dbd79fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h433a15d505b1e6240123b0682389073b6dc4dd436cb8798cbdd03053dd656ea4ed8ba024da47037fbe8815d7ecbc98a86d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74fff3c4a52414d5e2daeb3927901c5bc042f898fe0842d2510bfb662051f90e5a419d6ded00fc886df9f7c6d7cb4d79dfe6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha18d34d7d81db5d6f3c30e0c6f74a89e320bd5c40a1ba4d8a1d1400968eacd95622cd8fa3725d5eabc3bd56cc11a07cfa431;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h931cfcedb56f3e24774b10c52d087ab3d0f4ebbad6af92f5fbf8bab1b3b51763ba163df02948453decca35fbd80e8ac493b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7935737c8da0a37a9569959291a9ce66900b833b60ad634de746ff23223953b55dcb73fd1f28027d445849abb365b1d1467e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h825eb9706e7052168e8bb078eb9f31dd47e03b99edab7386006be94109b6a903af484cc2b201593ccbe079433dd66a57ee49;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74df582af6a6548a58167aa512aaf2f66b39481bd56ad4ccaa3d7137865847cb776f4fa735ba0277207205297e00d3d0c46d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46f1c3357d41f3c34ecd5d96d0148fc79cb7606f20eb823d54d13c51ee1959f210385ef157540b667de8d6e3314e1d0e7284;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31c645a1885a7f2de199003c7123ce45e172d9955315c6c4fbaa6c3ac22eea6b08e1fc04d4aaae9a7621e3d93da0a536b952;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2ad06736787dc411c9ac2e2244fafcae93152ebe48eb2b592f1faf55d5eb04bc99887f3ad4cc9f2e2de004733e44efd5339;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf845a2705fc1e6dcb826c0989a084447dd1de1423fe499497aa71e77efdd2ebf54041292c4525b452d6d054765321a1e6db9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h200b60c8447b8dac0a2eccb009bae387629dd3a2323388fa5846d54cf1bdb3df042d99594d105316f3e570bf9ccd00a52416;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c473c1e27f6826194a193e3bf54655de8eaebc32eac2e30af36897f1b1d7962e4c0a1695102ce0b5a2fc9514235ac9b04dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1398e8ed388977d556c19b9a300da1a16a17edf6f6752fef4b9f847454b5a0fa441502d6b7e258cea75a57dae061ad2a7be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf392a1ea120b44ac30c822fdd8e6bd600ba4da22a9db64f0b722d35aa5ef67305a34810ee1ad5f08e1bbbbcc77c30058c6de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb670ba10ad65406a80d5e77b77440fe4c67a357703ffd19ba9f0a7460d4f1560514ae1202208a489497a1673151fd5f3125;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d93ec20e0ce4bb968624fa6fe74c81492d2794f7a327e6f51857aecc33ab21318d54b7910c3f993adcb52213cc2b9001c07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha002e742303d7dea735867f66485654c6fd00cec4074df62fb3f44400905158300bcfdd66cf304e9c99346536889dca43e74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb385fc552fbe7915d276c95fdfaf92abc14d14329df95af34c68aba3fd88886581dd61373c3b1c48e3540cfe51f06cb9f6b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e18d6c625f8995fe0787d99e8d1a4659467df2d04a77b11fbeb1974f9aed1fd2b007d2d24663330d9b14ff17ca4c83c407;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecf0de96b9657e049a3b9d8b394d883d273aece4a130dae5eeeb607edb2dacbad213f5a7532e81e7c4eb42a54bb402921d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h403b5b02cc05a0d76fab1fb83df3b099cafe0bf88bffe20468241e0439968dca7bf1e66203723e457830ee11ae6acecec1ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcf7bcc2ecd83e919d4d4e6caadc62b6a2dcdb0890094b234e33e38605fefe0673d71fe8b515874aa423035a312a85b4d2a4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h171666f27f5622dff80efe2abdcaa092e6071c0c2106ac47b923b5d02cdfd9d891ef449a35dcce2dc0cd3ee5a4a50d1f90a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5bc022020ec131a841f06c056804306c0ce58360773bbfc94e71f474328e22c6d3e57938a3d1c66f0509d6f46ee0e720373;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h338bc5708e647aff14704a7715477b7c3bf2b6a18d656ca644679a6a51f780a83b24dad2a74d0d99e59bf5b1b67941efce98;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5cfd92e551d6b7d82cd8770b0cc424dbd1bf5ac60bb21aca794dce0a44067109138df110b912f07b9d95642623bb12ec385f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69dd260128d5716c6aeacb03f94204dd20bc5eef65d4afed368f22ddb0103a5ad268a35971d8f7530a846c88b9bd3a2759a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc343ea446131c3777675957198d75eb3f6a2834963b7422cbf80a25e87255a539c24caeafe30cded37ab1af71e055af869e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h573e9dd85f97ad1208e6c3e3a553b2f91fc57ebc61e581a6113529ff6cbba906254672481fb44494eaf1a83902ea325f036d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h484f3913026701c89de7863504ed9c5aad3253c396bcea1b2d36ee2137ca2228db58769e9c058ff5fcdf4eb8969a39c33947;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h879b35e10102092f489604b99b9c8f69f343bc3b14ae78f10c45865568305382827bc8ad6ae0a7cd1c61f957121b310f70db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92e472f3aaea52c1c02cc12fb472474dc0b3e4cbe61e537a5c115c62a5a835c58dd7d7270ad5e748d690a1c690dca69f726b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87b9e79ddd80ce80c1f10362d62481c3dfb4c55367661577798348fc5d11ff943c1af40046dcc34442c7f29b67b4f1c20c52;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h261a51687ef6eae703301d6493c25caae878248e7c548200b71a80a51cc8d0393c3047d6946dc889d93421406cdb3e9774bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3173941a7fde7f8151be09adad72f39eab8cb15483b89c3117574045c8457910cff973f339d8ad07942d8f27498c6f0808de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6cf1c57e5f72f6fc35474bc9a9a2d2b019b00911c650f1f8dd87b2fa9b2b1e5af391d1a9fcc3687356acf4d562f2fb8bad0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95485047ea4b813c616edded63ece2cb10e7c7b6ec5982f07282b830ad6ae40b31ae1d35dc7a0c79aee9b9a1906ffd748ac1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55826debe038a9010e4be58807193d6bb68715d5c94da35d5fb39c8e7fca27dac4ed05caf266e2581ed6f140a467bb3fefcf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8efeddd0d746015c66b56ef8cbcc345a26a8560beadc259f5fb83f0e91082180f546284f1b7646ab8093e7e88fd2ad65cc72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1caac51c981733ae0ff119ca28e1b9c4455fb2cd0a85c939cd8c6e36c4ddeb2e5dd49451b57670dc2bc877947be6e1f45360;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c01551914fbeafc52d0721bffd31a7af81bffcac5622746b5323874175a844164166b7bbd8dba5888b446683f34a89e4fdb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc01bf8aa4751f2a00fca2ab747ebd2cbaf95ae407088c044b7ccaf12136fe5fe99db6d13654dd39cdab3fb59182ddcb48fe6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b32170f6aeef0b22f2ba0f811258e789d3ba21ce8535dcce78378360c94a0e6cd37c38091dd9a2cc11133e9b2d5fd410af0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19d8c8e2423f836ea56812ccb2a060f716d0f89b5e8aee43fd11a83bac4b677970366e2c2d65e28526b3752c77269715080f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32ada52bf7b3468c70eca3b83c43eac690577b3f0ca9be9a4c88d6356f4a8205cca99812bb8bc183eeb8076bc656d89d148c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he22da9dab38348a30a90a506ec5fe77ec3384d7fb9fc8281ee5510062b7287e926eadb80b557fe743c4b715fb5b8f6760714;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3675dfce090d662f8736560409e77c3408a887d66ce34ac8ed02c454559222afeda8fa267571ebd091da18d683b3626a822c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47a84a186177496206056e2902543e5a0247d20f15a343b0e182942f78474624fd2f0f6473ad6f2ce5ab99edc271196e18dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbaf8c31ec956134b09672c237e9a84395665a565fe9f1a80dfd4b165930d6462cd1cde8cb10c78b596364c3aa7fad2ecb30d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb4edbee41fcc8441ca519e219eb2147fe1051ba836dff8e543fdb42282c2e12ffff551183d9a235dbbc82b17c46a7899eb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b5e867ca595b04dc659e15f6a7451377d6b3372773f24082e0d26431e7edc55687399507807ef7daba8dc4ba5b225f15993;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h284548d13105b914cff62542aee468a1e9f84596c83799bfccf55634c0c25f44808fb7e690c42ba3bc1bbe6da688e772618;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10b3100c69ce809273bb2524463b37969c4c25a0d98c6590cbaebedd63b83c8ec327c9b0ff01be2ef31c4c3651d4ecae0f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h195305a2ed7eed1e7febc43ddbb91d767459c6a84c9373a927e33a33b010964c1ee53deb4b94bf4f3c3ac2ffe8e38b04be6f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a1d709aba55c10e501aad400d22d32b6baaa9f436e90a835d03ad59a775dbd30de67a92924c869f6f9348b39b213cd367dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cbfbaa9d7e689a23660cadc3225649b36606e2a2e3537511ac05c6148c74b1b06a46bf1ef1916d2a9519dce5227460cb4a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf624b500c4e959eda43ec64ff61ee4f0f1f08d990f28f9fe423f73470e76f7e11fc35823a4d8f0a5b3e2c8048437f6ff9641;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9411fde85353eb1f1516db56daffb4681a791f1a0fc83848ab9d26a8ab762ef5bac89e57ba4604e90a77555e47be6f336703;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f0b6ed426da52ced2d65543e4965cd83469acd2e0551d8c615c527713e639cb859e65384814b3fbaf39d3730d3b86f913ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h717b9b03006001765620cb24477808e00a28eafc57d7af6d2d4b880c524653960c9eecad76d62e5a0aa3f8122bb38870700f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha86b4dbeef618fe0cc78083b8075263f8ac7a94e352f7dc041a2f5cfbff97e8ebf8607224bcf599c19c12ccf5ee00fdd32d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcc5f3e732f3532b1e12220a654608e6f8a2d43b1bf1d8eee1c118cd81c171b7d40986a91dcc336762450543b7f259f036a8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he93d1d2a982cc6ce051bfb36ca1c7efb546c2084c34afce9dc33ca60415fdc2d9156834e3867ddd9d4f0ef2925e004edc399;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24de49bea71e43204a10555e151d87fd50704b3334062e67748cc3a8ccb70371f1463f5b10c53eb2487ac18b73959a32f401;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d2fa492edb42192cec94cbae3d9baef828a742d5eae2ae4d889d8946018fe0e8120a46c24eb08e89e4f973006b23c8921a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a459556a9af6821261ba0df0d8f54b8fec2e79a205efa7dbc7e59acba84df92105a47736916f4bc9c8499ea4995c17933dc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aa28ecfac8f9e1aa1d6a8baf407db693a6a25e8e513f98b9ff67f6c490908ca6cf35ccb5078e0d021c6ab5608f8b26cb933;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he17b8f2528bf0caa52c15f4118338007017de41265bc61d9b9dfbc9775ef3623e548030b4d1236b739950365e6553d8902de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f7116705074c4f0b831748b163cb196e01d1c1c2ecdf475781e0222df6145c5f8c5e17d5479f293489e30598fe9e347718b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h651657a7dce6f6ed0cdab6117a5354ba4c7fa7a4410cb6c1eda44962ad4d2d8a7a793621cf460f87b63ae285f918aa9b1d74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbef2b550e0bc474fba0aa9d1da7417ad0934d688bd352c8827a735390e2e1c53846f50706c62a3c2b1a9e957fb95b49a4984;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb368ca6657e07215f4b052dc5bc8f4fee4d675a7bef5ae5080be389379a4c1b48aa2747f175a0197620691db3178622bf8ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h820ee08427d7755087094b5d3c9039322b307d54c47bfd221239ae7175f416b7e5dbd7b4b1614b7252826b040cf3470f604d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb95d3198af70d36a21bac9779d9dc6214d11a87f50a83c5dcc532430ee2e974294239f2d6f2f7bf7f2ceb8affdf664b47899;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb315532fd09c9dbbbd7b0fce87809d40cf1a2cd5d0c7f4dccf9c67c1bd8914df100464ee9f1c006042b3c97fa11ea8fdf476;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc305063bbb507a201a9baaf0f66934934ba1ffa03e6f96d3f537cde391dae5fd9999c1fcedf550ffd199b0edd6a19e013c07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h928b4f7943840c6a5c4b002272c654ae9049b6fb513bcb81667d1fa5bca2b2d5120a8adf76ab77c49bfdb60dce8027c0f0b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89a111f95deafed63da461493f9490fa368a80a31a72621606d82531cc2b4ed1134aea3ac5cfc03c5a22ba51a8ce9b5f1dfd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37e0209a36971acf2b6ee8d8abbfa5837b2686372eacd291c8d946a9aac9b8f7487ee1ad4509e13724bfbba57312d1481e19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf544d552ff69328db41d7a8d7017832fa7c601115263b25602a1790f0c03a2fe568d18ae79f270c87933a777eb2a33ce1051;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2150217b4b4daa5855f07bd32277a75ca7c92dd624584d8517d22864273a1ed56b7b8bc5119ced4dc6982fa9262d886cf20b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h702dec87687ee44e333b41910f672581e4728952496a332945f3fd95f6d7d0ac6452fe2f1d8106341d3305c3ebe9ea66ff68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4823277c2aa3fbe3cc5e8c9f905b708926b3dcd7cb961d14ea25c19071da2afc59b9cd64b433fad89368403342139ba2037;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec406bc763217d67294b4a57943ad9c87761088826740a0990f577241686e0b16e65bf2d205613e761b5f7c5b7aec574e74f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1222aa37a6821002ff7d99be470991b25e1c2bdd35e0f96623712182b215ec0b3be43f80ac8da98ab85e4c2a3a4886cc8366;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd882294d67993acf029816aa38b858e603ba79bb933213ffb6186f1b0c1efa46e458e1ee8e5c235a709355c4670bcaafaa8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70cb686ba06314e2d853d74a95d0f0cfeaddd9b9663218f759ac786ce0f7cc9a7c954547be704b1270a866aa30224790279b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h642996c19b2c6546498d801de0b18e2b4681a1dc4fc06c976f829187b488c28385bd79f0ecc546c3779bab9c1b32bb440da8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he06beb853c748e17389aa91a393b2f82b63bca64603ec256a9fc0f35a7e0f7596782d7890ecd30de9ec7f2d56841211c0466;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4af45500c8de06ce2fc39867b4344cb4ad8d1d6a1fdc22f6e4764a3ccc11c5ad810e08fda16f6e9435d5620be15ec0a8ef1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12bc6de06d14ddbf2eacc3615096bfb9e35cbc751bdf8efdc9e897f75ff61b421a422e02b7d3f670ac7fbf6f48b0fc06476e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h265f688178dcd6a93117d3f1cbeef3fa4cf408272723f8008c776efe16e7c5512fe152878c583028984ad05cc23cfd7cd7c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22a976683db1363b882ff3ee7f661eff6ba89df156d62db251c2d5ea0d0d085e94446af1a5aaa691aaa52acfc58ddddebfbd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5e208f9a911a31094209c83e5e21a60f023437a777025f13b4a48cdd7dcdeb1b1a66955e5dc974fdd2d6f882b5aaaf3ac35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h298da827be586e1b00d6eb3b28f6ba8b3610f4b942bd067bb59b174c3919d32d0c6e1740d2b3835c6819fb5a30c8bded84fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4856ae7f17013866f1bbba0d0a3e4655c43e5a3a783097d81fa25cb7aa639be67870d0a3a3b843614d3d17d95e1955db21b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11aadb7e18b8e21ff4dccf59afbc1dcf07dd6a0e10d8ae1e394da2364ffa1360e4b903d68762c4a1e59ea4c6a91269a9fcc3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3008b2edf10013415922b8232f31caac2faa356c9e8cf4f55f47df4bda92844a62bae3450c49fc6944146d7146e1601e44df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a8136b9c15ca9bdf36fe06af5c765ed10baf18717a891afd732af5748dbd109740a980bfdc8bc15dd8abeef95c4694aa3e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7bfe988825306f9d75e1f1bc2c36e887b09315bbdb06d9efb023fb7fb26e9c5f17b0445b2a05d9fa174dab3927f40bd8a9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a99f486d380d9e77f458b2841822504abfb4eb2a0239cf6d42e69c8f2ace00e5612182e3e55375941abe3ea48bb652a6a04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h342b9865366c675ce43be537881d7157ca1a799352f5ea0a3a9a9157f93f5c061736c78edfa9ad78096a9d9c7ff919527390;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2c02548987c90819d6e652b3f2a22b99b5c8fc248fea5a70bd2701250d5216f7a38d6ae1df5b55e0c6c1ab0873c83e4c4cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65079310d8b3dd0734c354061add75d4dbaf71a9615252c9092621eba928540e62615924a5ba277bfa914726f0f412c2fcfb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ab4a98221c047ed44fc215bda08dd257649c40bda31dcaa7852495d61c288d8916811ac928a3cc2803d4874b482bd8309bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he28818e5abb3ba7f42622b368407a114604d8b2c8e36429b4008840f00067adf0d2d24b227e90bd7d313e06334aeecf6942b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae6a0f89346f0aa4e6dcbb11ae198d84eddf6705aa5f0a30c30c72c46569b95197bbfd4042dc8f4999d4bdd07b56d51776e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64ce67a1b4a078432a6fe62f8e7d25f785e119b90283ec62957c75b922c2d5c538be2b9d4a98de791ae3061c1ea7752935b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3717e86a140e10d644445c7def187545673777ee12e0e641c15debee4c19ec3926f9fe036f75c3e12306d2a0f423c3d3cbd8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a669ab87babf929b153abea09325074c5538cba3ca7ff415b39180691a5ab70f7d7cc36a393c0fff2ea2cff4f16075aa8bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha000bdca2be2f2e9cdd2fff86442e4fc6bc75ab628f4d81e3b96c766cb67527cabaea03a296a24bcdb18f34ada58298df617;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f50d9b8daaa7d6474497f79857c2481f3947658b82eb4cdad965e3f276f88d96cf532d92137c173369399db461f9e219f77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e80803bbe0d9134e17866a3028590239e469aec2ab2a170bb8c03cb963cfdef8d9ad521644a62ba20dd7a7aa0529fa6ceea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfefef52726b7cc5cabc5ab7636c4d6268cccb9a493a3657d4e41614c3472c18ea0267fa445cea5b69af0af3276616654b930;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab24ffa4a7daf6abdd720539f3dc8bc723fe776aa434fbc4a743dfebe4a2c6b85272005e495ecc82f920df7b4b38709ae647;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57a1fe92b4fa58539d00f67f67530732ee6a122fc87e6030f3e7450f11c7ce34f0b251778fc13706171784639b2f519d0de6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48a6b4b7f141f7fff6d7192ba29d2ef4baff9ac31cdcd6e6d1cab626717839c33c9b6e415b008a4d8feedd54cd8c2e188e6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8e517680de636f52b53c9817efeee6093f90eafbc521a9c001bf210f8ab001a4a4eac58e7185f15910391dd9f78295bacd9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h370a4efaadc1e8d08267922e3d03c8536e0fb851ddfb575fec0769475e8903e1615ac13648c6003cd7056d8e2dd99b529f66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42c871f7c84826fb6acbce2a8146cd0b59b1d40e21d25372bdb01d647a52ffe65a86359d327725d1fcdbfc71b16bf79ee241;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8213a425cabc3bff88072897970b4b990dbff3bae033f38c0509b007d59d870c2e8745922e6d4a0be32a1e8cd67cfbba3f13;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75eda201362e4fbf2e4e15ee67e80c21768882203547f4832a253d5ebe7971519b3d5ea82d11c3a9aacd012a60d8656b5bcb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd124ba989f75db300e01a9520a097e72c06edb2d3baedf61d336014a9019c2390a2078d786cf455a828d82e1af40cacc149f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf85d3ae3dfa49d136f43d936ca5c68429a7faef0ebf37c34e1fbb55e526fcdb656eae35226c7c2409f28fd1b12c0b305b96f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6f98f26a850f7ce8e940c0b4beeb4bd61723e5f8d356be1a20ac863ce0f26af7b3da33b6d13968097e3546b3e958cf75c7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haea01258cfd5b38db4516725b0c738c9c2eb69154808f288a148884fa3d7e0a627d174d28568433896e46c0eba92275acd43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h582fe6f7d54136ccdaf90189d137eab9326abfd60cef66cfda71af17a25c79124961291c332f8223cc0520241ac00f0e3b2e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h279cc30c4f24d735caffd66a2b2bc82a38642397690dacbbfae0e5bdec3f624d7720613ed4dd2a4992080ad56f3e831680f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64e6935b0db1b5bade4102db36af2e2abaa08824d05e2fd1aae0aaa8c5fb11c139ca7639cc4d10ee1b878db472e27caee52e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ab4531761720f2bf13755826ddb22931cbd1af5e87de393c53cee06af7d39f13b5eb12e8f9cadac1d00f7e89e482e8846a8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h735f3b16a36e232d40118cf9480b917d16f745268a3c38644cb69dcf3434ff9a3a90c9bfc149d833f86ac244b7939387cbfe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ffb2856eb9825425e2efa606d21a0959218d96b5922532fabbed0aa7eaac70d06ae0221e44fc630002f586c901452c082b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h629ce5291ace010d743540474a2277907def9d4da8360ceb7a0767fb32b92dcdea2b62a3d7192416aba778bbef8d4eb8c64b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dd162dfe60d5521d63f8710928f463766b202f1a306e22212b69a0328f6d553286daa8a542e8adfd82de8ff5a45836e832a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fb41d39bf8209c34e65df2e0868ff6dcac307fd966972af4308c2e6fd47cbc14fbff0475851f9173e1fd3094628a5c4390a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88e1583d06d990a06107a8fb0f2e9ae1c2bf9ad590cf3bb880073263f1e7f44ff5a102699e5ad2992892364c3535c51d038f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc3699c25035b076e9d217e41ea0307197ea485cb38c3466693987280c7a6c5642c4d5ea648b41f8dc765834246d7e4a64cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc44e7714c8817128bf571bff734664b03b4e5105e3a95962e1720450a615e2fa782b4b2b457a1dbd39a32a60e5954d83aee2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1c8601757dad4457705991ba4e89e4ad96c1b035198c3bfe12ceb9d722676ad67cdc6f5caa35238c90fc878f6b6334f0295;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h482d6c802c67006f99a78de918a413aeef8531fb7a09d86887b019a05c5d8afe2489afa5a9c68659d1a4f964094a81f62b1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h152ec82902f56c7e6186038b0ff143f5071d72354be2708f9cd96f51d0d92062137262aa5bade2a08310d416afc15a5ac2c1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h984e0de8420abe6af7c5b10cd24592dc970280a55e007a79931c75e1d1718d0f4609ad764466349c5d20114466311c86f721;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1981987ae8009a27ca7796507b9e33e9e8e108802dfe6ee9b1c067a370049286d50422131d372e69bd9ac74e4d083541e5cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e698a71657f525f31555b4e85c325ba47555f912a8afee7b280feb73d298e4bde904794a77563377178b9e8d96c84e67141;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21d4858509b2795a6152dde01418ae345b7da83c4d2d96f3620ad86c42c67736336db253b8d0cad8e4d90f03dddd935151d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71a7fc413094dd668c96ecaeea722d033c3da52f3d1c3ccab2406f5d9570fef325f96b8c62162c8c0047ed66294fcf2b81c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef2d9ffe4535ed2dc44db2087eaa6c6437d14e932e4d80330072c611aca169d3745fb4c53e9227dc09de5319901530fb573b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b7fac288dfcff1ab1c34742e04edaefd3e8df8ec4a9898fb90596e2ea2a00970e85cf1142dc5ec6295c078f52719bade9c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h944d0fd66ff0011963a68e4489651f2e288ceefb13549d92832a0d5fa7391187e53f5a04a00d6f1e22fb5685fa2394169230;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h574b472976e9a3bb3028879e115e07e0c5f4e4e37a8376d16e9fad738eeb214f33f55582e9e138afced51e84a284430eac34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb40f0f240310dcc6a18804e328bf5e18926111b4f2e407c5cc97f72cc26df5f0c9ebe597827ceafcc0e2f1496d15ed11de83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12f5c3ceeb0835d71bef29f05b2650297d2977fed3f7b8b9c28e7915e43597e20ea2ce7b60dbba005816c8ef0639293fa89b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ceb7dd6b9b284046c4c8e75bef10d4de6081fff2f6664a4388b50388c9d7ae7bff9d48c2e1aaef895d51ee7ff0b9f787f32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9bf808678bac821c730165bcd437ed29a4405f3d6d2c279debac8e6e49fea3e443464fa0997bb0080d78b0573898b98f6ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ec55b0c113e5828f62fea3cac28d40bc25a5b8603057ad978bfa195ae50b83aaa1229d1064ecfb1037dca05021f8d4a01c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d8e7bc139da6a78e6c3f14d69032c91f9a9cce7708ed9f75ab36e0eb52ab827c56f60deba62a8d0dba2ac99f6b0dd99c295;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcacf787d6b9d1baa5f0ffcd16a5e0ac9202ed4b07c1eb358b200005f040383828a1c034ac4a1499e4f1c94a604372501127e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1850185fc3990fc919a9ec6c70c4b6cc83f6eb07dcd7c10dab058686a04ea74ce8b4f6b19c5bc11f92ebcdbe7e7dfa27d92;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb70a23ef8a5c69dc59577d3578aa8cba7fcf0da4076be6a18237d2854e05c4d83699b50d709767c511cef4162a93f1ef56f6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5b440aeb97098e4a6bf79008072bcc1a4de8dddc0098f61b8e7e64e2230bb6c8ff8fb4a50e00126f0e2b2e7239e5ae4d981;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b6f72146b36e1a97179a3529b04503b72ff3e783246e64dedb31ab2adf2199d13a43ee1b33322c9720878bde2bc46e1ac65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58d5e746b2e7d15226ff39dde3d5b7e9ce54ce7fdea071108ae499ab57ae87c6b4f6df538adab1d3a38952a85f97187bed08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h102139fc9f61f4ffcd7c97b1bfb1f1b4a9887cf834bb45cfe63f6573e351d8eae053a49b1c8f5f97a1aa51b96a2ac6af4b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80e74ed6b9703c4d22bdc1ca166dd53ef4223fd03e715f51514f4b4598ed4a2efac60038709cf515a05500b2afb9fac62bbd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5b4fea3f3c637d77f634e1c350a8c093c0de30bce02734775a4ef4444a6705bd2bbabf5a1177b2f1a8f3a0b8c2d859b85f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5c5dd0deb430adf08b7b108898be4b56b9791a4793fb06d6dc96770e37effdfbc19108fc7818e03da5dd2df38462a98b345;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h452dc1483908bad297c95fa85e4432b2215832b77f9f9597b23b3c115639374d2bc689594eb984dfc70a4d43ff80d7836a4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3918c26e4ec130a3333507759d51aeff15c972c1e05e6cce649527950c1ecf307a8820ee4af2d42ccbe6206d2f3d3eb20cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ca55d156b1b36315a800560a0ef487120d23bec23a59163b6f2b297f0e15ec57efc9b97cad9aed6376a30a4ee0f7d70b5c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h476c5988081a6b2639321a28d0c621e99a386294107e6bd43cdf0a7bc7a546f68bd999c306fe9125a46470d45647903fe7c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9edbe9e769779798d9879648c755de8f7fb097f7915b3c0c610be918feefc24aebd0837d7119520e84ead3d5e48c572a6e11;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8646824c5b07cd0453a5af79af490359608e614dd1b009d86f5ece58989c36a0ddc01fd47c0ea9cd69de2b5ea242059dd82a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97f075eb0ef7d759cc2c5db63b44fcf3180d1c50301505130ec5ba2e01db60c3cc476cdb524d13cb6a22715789ae08cff52e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd2e654eb092914c8701b0796ab606a42b5c3907fe7ed489f59bf233030efdf412565aec95d5c2d1236b2ceb7c94b4380f07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2696d520e33cdf1b84e1aee6ad43fefe536fa65128c156fdb5d3d12b7467048595bb089eeeb350f83c4ccd23ac00d99540c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec549f321b2933ada695808c8038a3970d1ef9f3bc9c95cef68a66d43f8d8b8699d8c78dd7f3e066443a1690139ff0a61488;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h955b03be144850bee9066808698c66d3fa2ca12636a18f4a2a7a4c50593f233fac4deba979b409cf1cfad93197f32b452173;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d54acff9a026cac79431af6f4a128bc3e2d20d72473c89d4ba64fb1adf0911a153cd8895a85faf2fc68349bc213d5f0c38;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d2d746d77a121e79cf004b35b8c3c6ce2eee359e4088e400b5e1563ccf944485a61a13560e80d9d0cf32a521faa4bb490b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed62e2b19a6fb079ed1c55af55c5e6639e6ecb74df3b9e629c2845782baa4c6f301d35d24866b2dfa542f5c199a59a8bca9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h608002b36718222e81d798f7dd91b3018ccff92ee9cd8c2c8759b1c06b9f04b87d369aea4523821da07899de2f57c5b5fb18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6eef7c3ed2fe2b8521ad7eb2340fd8f9e2090bd1794f68d58ed0fbc9ccc9ff7f0292958bc33132512cbb1535a53ea55b227e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h181a2f13e9ed11e981868dd7fea8f459efecce644c4cbdc7f21194e9c629eb7229c563f0213d489330dae84ef83ab624956c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f90ea2c770b8ac8abbf9b0f2829961637d15eea7ce7abbea9a6b1cc1f375f1bd9249291ba17fdaca4651f992d708dee9fd9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44af2db71c584fa8f8f8f133b3ec3ea2c92ff47529dd97080ce6e7b99985a02f6810cbdcf8d1e68cc8b28821a1c5a2be1164;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fec661bd6bc78551353d7cfd75e87a0a4e766470701ea3c61f0069705619a5010b79e309ac4f19c8a973e1925bc9644b55d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h667e09ad003e52f3f73f4d043f9c25c50ceba78a19921a00cf87b01e4c3f306770be20ea7149e14ba07f7131722d3598d299;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dc0c4c1a6648d2677f5e64d5b096b5ea02492e4775cf441b56ce4ccba4b68f2caec0c68678b9534b59852411c60d01fa45a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf67b39451ebdfd21f6f30629f5ad4083c226e7970abd46cf6eb14cee1c95525c1654f6792bc21aedeeb7bef9c705371bedf0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb639e0d5a24cdf8561075ce4e86b3f3a9d37bb81c987ce27e7d5550a47c68dcb16835cc7382551903cf6907510c903b0259d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h714b4f47fc836a98c88287a84f29586cefc75f1e4d27751066016775a0a4e9bf0532a88781795b9a0a96bed6d0b6a8a0a5f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92d8db00b426ffb2d15b97b2dbb7098ea533a5ad3ac8bd317dc5469ae301ba49e38a1dfe36058c1771f7cb175c76bd2bde2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a7b16414c6daf41fe90729615cfc76b7a40de2ae9ab953fd9c9a2935174da53ecff4448df1f68e5d931079955be54b7ea7e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5cc356d926c3cec26637c3a20909060d7f8e6c7c56d5fa6523611ec72201629acbb93b0c3d22413362ab4b9617b1c5f581d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fcfac2697fdb900932d93ea05e6c611c5eae4e015e553d4f491d2e0490bcdceb3a90af187ade08ddc9597c2f9002717b1f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd57d9d57c53d31bbc9505862515a9dbe42666c569bceac69f5187385218a65badad1e8dc7c1c20be08e946905d3d1551a928;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8dfcad28ccc8281949947006322ebceeb5ce9d964ff51b31ec8fa56cf27b4c2050ea605daada3e72a733f4111e520a140cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfadade15849cc69547df6cb9a27384990e18b5381b8f37707aa758c029bee1671ce0f712dad4d543b65bce6138bc0019b7d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88ef6de06b00091de22234957300a44289e6827c99404df4677268d3cfffc5feb3f78a98378dac93693e0b80ecc47b4416b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed588e3f68d70ba67fc4d2bc16a144c547de4d6834ce35c16b8a10ffc86776451e2a1b42e7dec828147e439b86cc4f3f9c8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a8e598ffaf86314165b987331ebae9455783b75ae5d2f795167a069cb99777272902d4e880487d0810db9cd7c50209a8ed5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h793b49cd11a55f8ac73538836a6ead5647f3cdfaa2150d1389e17a935e5c4fd6aa2141a4a70231bf6daebc6d4f2ebb83f320;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf558779ca85e66c936c0ab83c2214c3bbbbbee4f4b5c6e4e91e27da800112335391b0987a4ae72da7b722b9efbe2f7acaed4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bd70f263e606b27179c125d5b7058f46d9b8cd18452e9a93cbc706d3bb8d4a28394d0764a419d16e35171f15e8037b6019b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d379fca9578296b58fbeed7a352122841b836ed1f76d176751d228d672a8320d9e8e4bf5d74b958e0bf806b9d8f9aff99e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79be806740296b057e6b4ae1fed9241c8edd1360315735dd4b32d77a5d7b207446e5c646789f705c230eeb47bd12f4252f84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec32c062dea765795c25968a34231c559e94851dab473a5a14722776c0e12ebb0cb4cf757642972eeae2b832f9624d31d9fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50e23b5f7ab56b1006de8c80f850a0b18c3ffce7e369c43260b012904e71b4c27e9705bc3e74abc614dbffca93aef13882c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4bc840bfcf35def343bbcd0ffc960726d9effd624e8ea21f2c094070b0d9ae240c6d91bd515381806dd03b0150cb9bac26f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdefb7ceeb350c2fb61d4d290207ee6000df7520ebf431d311913ea54691c9d9277a9c802f4f8714fe24fbc09e8850eed76c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b5b63ceaa52ebc6f219941f8c78d0f7dd766dc7af837ab46cda32f54449d7f9e66c33b1104f38263d251b761c59c19a0c7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc98c1d4b41feb0e7d3b7661f2ddd53b62d6eddff583fe762e6f90c6376b474130c56ce7570cae4ec5ae43933f715704f1bb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d85ff5298d6d6d80de4b87cf09a28eb388bd9cb91cf5c633273f62b6da5226c60c598a1d0c1e32d7819725cf3cbd08a3e17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cf8fb74c9eb1c3d01839edb9d6e2a1a94ebc39df561162890952258fdefffe7d71d81dd438281cda55a3d28cbbeeaf03a1e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94aab6f869df5d1e24f0f4b1dc227ba860314e7037ac3eb279fa6eb1cbb393758a3faa34d42752dde154ff28fb498d15a6c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc86702b6e5f9543b8dc6ef661b5c7bb80b574c54b9fec634360daa1e9ef45167b39e0d450144640fa1f81602ec86d3de8f74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88a7412d8272ff31020400c715e8a70f457c0ab5ce99213ba1bcf6e333993f565b01fecedb442431aba625ce0492f6267e3e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6b0d20244bbd420798119ea70e5fba4bcd15b536b672a37154b954e7d0f234ef42a94610d39a989070eb48188b526cfb279;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3d14a0bdf1d302ea29631859a38a0009e2bfa5458f20851ffcc9c92f84beac7b06b35ce845eb14deea144db99d05bdd6da4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b8632e637038bb6787fdf4eba070cd751ebd02477b14791de6930306349653a5cc9cb62f3beb38d40187561e82a585bf64c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63659e846fe4e065525efd7ba5021bbe25bd5dfa04d50bf2d659476446dd598cc67bb4b479079a6f54399ca076d2cc58e728;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22906427b82ad2233201ce2bef0a3eaeb16a0df6b885b9cd59852bfb5936a75b3875d2965607acd81d9c5b5b58654ce1b18c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ec347c1a9cb0fca11ff64f4a4ff39cf919ddcf3da7c070ef5bf801cf5bba491e05f4e9adf037d624dbea52e766b03cf7c0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a16daab322185994c3f0245825084aafe6339247fb90b221a15918c0e14faed831055c4951bd3a44c245f26ac3cf314b464;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69cb1b0d192c76d10a598c27ffc96d2758259dc4ffec8dc9aec5218a4a965b53942092bcda508f4ca762c0bc88e9f5411552;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfc01fba3292691880180ff6c119c553a17d6c50624b86adac20064ad874124afdc7ebf643a650055b6f6af39887d2e6d49d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdfaa177b75b70c0f466b937fac35782e31ce3ef242fab7b49d2fe2925320c71d21e40f496215a3c0cad6eb06cc458ca1395;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he747eeba25ff27a39c120268eb058520be9d2c5d148839d64a3857933127074454a995c2022f464395d788460b91bcfe0ab9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23e32d03efb369f90e944e7a0b70c9ef1f97d7f68762a7f91367c44c56f27ce0fc6503d8cbe5c790d4cead4965387cf24d58;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h417f9ad9a5f2802748d1b9a0cb915ac82fb5b90bf514bb4fbded1d8ddb97d471f53910165af8902590287d73f30e7280c6fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9a9417fbb4c54a0f2d0ecae242e3c92f53b73a39ef7dbf932ca65e31da4a2e0b01ccdac3b6235058dc955b242f696597e2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72bcf2711b6c1601162f606ecefe1397180873d4f15e1c9343427ff5db90aaa328dfd27641ff4b01a9f274746880932adf09;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed94258f526348aed271600c1ad401780988a64568d7449a846566089bfe210f35c8b14d116640fd0524da5aa21ac814817;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h725d3faf3b7c3582038f88b78842e2e41a270e567002e387c261dc9de3e6d5bf0c90c9a7494bc36271788f1b3ee0a3416d7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5fb640b4ddafa6d5fafd4a72376b15c8ebbd0bae2257170069f790e86a3eb8c64a7961ad92fbd04d657e36f7bef4121845a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a5feee421ff7b4b9197df5bbe1fd015f57aa5d1f72db209b127e1911c92c33d6d1edc04da6e5c7488603bf37fcf7bb18fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2eb721e61457b380dd479a3c91e310a490445f004faefdf612853d1e5f76e0f0a1da2844573785ef7dee054ed7d9d512b3a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb413cc24a499345aeab1c8a8acff67cf0d55b44a7557eb6553812e06bbd428739f2f440d5d7f6c6b067c5922f2b66822e9e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8192d0ed6860aacc8f34336b67040cdda922c85e78c794db2393996297f7ded877afafb31ffc2f264b66a5578af6ffd89e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c92c433d1a51da59a82cc9a41cd3ac5a9b2d195b5ac51e0c940a147c04daad03ae94112a4018ff33a814da8cd72439df828;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha69f54e79c75f86496836b48aec2df4dfceb0629f1576580d2d662f5c788a57f8ae1361d65655d8c7aa95ed130499479bed4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b222396a294ad041cc16e1ae77eec6e3ba9654c3876b648354b8d75e62566498f320193424a99ac143c3f32dc305af712d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72abda3704ee635cfe44283e6fc8a07b9b5592dd3108ea520f05ead3049d5df51cb6a0ba1612c4e33998eabf83766c62b952;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fbdc1b921aa837ba65afe5d25d96f1660297af05e1b5ee9c30d38e3fce395e64216abefa7aa80c78fa111739bee983e932c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16e25976e102e08b8d69816f7459a37027b52c08127b8e3abc4a163569b3cdcc506a55b6797049b213250aa9b4c3d5867840;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ef99e5c35b85cfa9d30c5dffd0254ea3946f0cf8c445c3f1153baa0ba768db449595663e84be3606ae99faa989404725b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4223ced6806f6626f9a8d35d608402529ddadaec112743aed9c98ec392c2d0a13dce70bf14299e91dcebedcacca60245bb86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8d504e6eb7fa0e5756938ccb6cd1e6f35e1648bd5353533deda4e15533a3cd39c0913ad4c40ef5608c9bcb9b37e837116e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h746f5f9ec9a89a828b68170924d8a0c72a69be3a33916fbed58d8725e4b7efc6301c6b4511be9274f6e2a09510fe102f555f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7294f3d7a704091131d869866bc116a29c348417e2339c07f9e9e42924ff0062a0a6889f0fdc2c8654fa703ae68aabd4829;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea50002319c38d5524551baf5041cdad27d2afa20b314e44f2c08a36d56a80b2032451dcb91df17ea5d2dc9eb4bf8bd8908c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ed77cc7b8e0f6d918d55e7cfbb5b68e094ffa4f4bda058af670faf727186fe73dcd044db333e7306613cbba46476dc2ddc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h254468451847a145e4232d4e5d472ef5836769c9ada1deceb255d30612b4621094ea8a79f453f4e29f1a07628d0720d76bfd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68297a3dbb3ec82c0487c91c4c957559bb569ddda306b17370cdfbdedc3d3cf9a829443f147358c440fdab370b962cd5e7a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59605758fcc10a90add85de12ab7bd29e6c81d5bdfd4cf6df3761251a57f7c3c7da9535191e2b9910682b6515f31979a9e8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15516d44f3305667ac5326d7a75907b6372dffee0ed62542a57a29973f0234e2c3b65c3db19066ea1f4cac3308151773512f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb158bb49d63d207f75fe17f0e6a54ede2bdfd27303b40db1755d8bd1ca2924daa5a70fb1887939b38c4e6833c260c5f89818;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecc81f9653431cc1bf494b2b44dd69dc1bb67fc59142bdc896ad3f84536c597e99c301d6fd208f200e6d8459a3c347a8ea9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h114394cad537ad2bf2c349bf505f34b21bc2ec801b6b26e973eba93076b92714d859225cadf741163928989cdc8d5f8ae167;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h375a81b636a3eb1ddd384e6939d07962d64206e15160f55ef2e33b74ec1bdbe6628d10d8b3592dcf390cbc245d6a521ca08f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6566184c37fede1ab64a1e771d3c2673f0051c16abd10dd8143fc46792fac31017d7c49a89cd6009330e2125f5c776f64af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h241c9260b5779b927f4868f451cc21d4aca8e8c209c5daba5a4ef13007153789aa875bf996cae1ffada8765c6d6b3c0a4843;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8b5a9e5b8cf8a5af8b9fbbad7413702459e8518d2521563d5bdf469c93904cc426b824dc29cf11f1d1d5fb04122ccc7b3ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habffc17da7818b99569cc376a56c515f97c027703642301dff6bce30aa8228d89d454718befe494076b95899c4dff1d94967;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h345b18a30f031de9e1b3ca414d57f7243ef08bc79ddb77dc45accc0af1c883f6614b33b085792411a3e8b2f95c99cab6f850;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9da01355495168b3cc6e89e3452b65dfb0e84e1922eb3abcf5762b99a08e08b139571a5c482cdcfa43b913389867e1bf4f69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac2aeec531c2ea682c84853406bb0e774858139cdf27800e893e57065b472951cdf88bbcc146ef5182512e0dd49a2193d1f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8b22c54593d58648cd08634e76deb058d9ac260c3ef21c731a13ef9fda3c659581cb0e7239accf2bfd2c076847f99223fb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bc09f8de404ec8499dfa493dd9dc24bcd78bd065d90ffeae660e6920e49b35ebc65c0e5773c86c06d7df892290350927e19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6022322450dad82af799251ad7781da7072f68bc397e4199988de4ef0876403c298af644df8b0e02df873af6b634127ebcad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e22b01779c1703e9607c9d53f58871d2af9099e6dbcbd491eddcc91f25cae9ea1c97ac273df21e40119fb4cbd2d95a9554d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h978e24b4c03800393d3c8b36d03e3a6a69597306d07350e0f29ac04da56eefa55ff4922096c35eb2fa6b5a2eb1556df5d0b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ef4e6726dfa2e58f846fb746b4d6eeecbe4bdf5ad70527ba244fc99d1bbca9a0d8fe38646108d81b31342bbd137aef5d7c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7592c86ad4d9221b644ddf4fdd48cbf963cea387c68416c428cdf9abfd205819fb23b157f7c041e67c160fcdb55758c356e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h127cab8614fa03da3360e5f8f011bbb852bfd892c151e93479ce6d1036d3398c453b1626076f2b6eec79fe6ddab168f5a77e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h965be258bec204334c3a51aec6fa097e4049e5e9dd46b1e20afe1f62e258a8bad895f4fbb7ca798d500e6688e4c2b5a241e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ecbff83b83e5143960ebe18e216a5df139f61bc63b02edf1f5962fcf14da19cc72b26acb8c942e8ae3122f2b4702c70120d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4822b08fe5abb73ab410c9d863baf768278b4a6083a350e77a2806003d3fc8050c07b30726da3be2654ca77d2de94c3195c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12b465531d1ae0c3353afe85dd44c57691a820167424ddafe56eccdf0c87221eb48a0b2eae9a4ff912219274a66dda43e907;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8a1d189230d7bcc0ab30f66b06a91e0f48e6b1bb0a023546e6399d51e89afdd3877530ecd15a72b4cadf89af7809c17f375;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ee5c3f55915541ac45550c7ec652a43b7029f05f8594d29c955db874445271bdecf5ad1c156acdab41527f6afe0c228b89d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7689616530eec8889393613e89b16b6181421ca8c0fa7b271cc402c8cd034f9b9b16263882f743a43da40c297eaffad6c323;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa3c881c07f1a44d0034aaaf2ec94d7db017321b3e637d33461cde426ebbf28d35b927b037a6dc2638cba55d54fb0473e64a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64315fb0b1a1f39bee87a05853dcc501ecdd94913e27e99bf6f3368245f183e7f000163efacae91c0653f2715357e49df7c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b9a1d5a03a11c3d187a7f302ba75c34340e0ef2d060e3c2c27ab2458022a42ace079b806e6768a4d4bce14746cfc6b268ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa4ea39c3b83cd8e89570a9e047d6cf990586c662fb26c55c0141d2eb9cbec7c5def4ea8c3fc345095473beefd82b7817640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he382cdfc7d1bcec154f4bb975d338ca1e5849e42c41881b6530beb33a02d2a71b210899887c8d6322337210c6f4c346d31b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ac636fbce87b3c0bd0e351423d0341d60f2f7d07c5ebad62b15f57e743f4353ec279be5cefc549b96a997f375b304094dce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf573fa9e631a1489ad5310187b4f0fbf7d91e938ed1fafb8ebdc072b08daff57b429488e77b71dc75c0b164128e36ace2bc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha62c2979fe2ae2a24a5ab71d9684c1f36945b3edcc7f56d94f90a1ed5df7d507e3de302ea1e4b5ca1f50593d72973a38bd01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea1f77586d7ca53684a2439e6f8c9f8391560f679b3d99475d276c5da51787322ab4661e0600a71d19cf1dfe7d7d92307e2f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cc3cdfd27b01876cba60b95d76b2335f873fe3ae473294944cc15d52bbe56d05096f80d67edbb82b903d6ea5cbf0ceab0b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc969486595a8a72e4c617b5efb5b1556b1a55ad59fbbe1b7c2db10f4ae4c4a053cf5ef2910adccf09b5637c20be87888523e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3779f0e6f9951a47cc87b9c45c2f6da190523e8c9900bc690bcd7fc17861f41f06edf237f4dafc81fc4e4922d0fea1d77898;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b76375658cc08871171b8b83b8d9a2966260e26073381ef7d027cd2e8d50fe979f9d44ae67f9ac1926b973452ee1bdd8a0c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5adedaadf2877646a216632953ea837c2de9f9f7e83c1968131c37e9d5126d6a10e27325f2fd4dac1781e1fc1a610c87bce6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2f561dfd3de45552918605ba7403c794c72465cf5cb9379b93b44da9d33ebfe7b7c3bdfb09092996ac15bdff571e2f38ad2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd01746c61ba32b1f257af63992b597a8d9a3a2088dc24dbd7d8cb030b5517f5e1b51f93a0f965b448b422f0f65a0a0007317;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h441683b17cc245af9501499f4ebfd8d2c5f65ee438c9bf632072725ec7d1375bb79eef4c4340b60aee0d762dfc5d3e1ada73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84fc1b183fe5d66863cc65f31c6ba4ee5619d8b81fbc3d4db7ff73e3bb97a1e2c97970b23da3b12dc93c25472b9ffacbd59c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa26c22d6fd2357ada0b27e3a347b78d7a780867d0a9c375c98b3daf875b72b34224ebb0009892b37187f7a0b7e59951c5e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5515ffea3b09064dec11c73623a2ab835420e4641ef41cfbbddbbdfffd1de5b5ea5e6d7d1e79baff638d73d8647fb72c69c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56cff3ae2644aa13783a6ba0359a95fbcaa2e8406f03b46fb168b62a2a7b475ec92f4110f396faacc0bc2245c81c7985b50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h766bce7182fd7491577c9d0c6b266e9f00502c8252105a7f89e9d1c5756c8600f2a216df9a0e57d719c0b2fe066eef364a19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc125575845afb48e607122fa223fb2fa861c5c00612555bee41513f73ccdb45ae4e9c5140f11fba3eb570e03acbb134f6501;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9bb1dbb5a2247d04b140cc83866536eab9eb3b4257c9b3f7a9eda4312d1ba790637b6f8539317718e86409435f0dbcb1bc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5723ea685626c9a5cad55eccff1cddf93b23272f4405944f45f135494135583566f4a06e4edf4f5bb0645a0cc24dde3e4231;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h789ce6b3c88e8ee009e4cb0a5b1577c9e4d5950a53868f52fdf9f89595376db66a2d2c12d4cd8e13e627484f30721f0fb8b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d413a8b099e59685cf2373514730822af0c18a902a7afebad537a8e27b9b05759d40d212c659ec1b4f337443dacdbd7c69e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e59de19eb04dfc27bf67ccacfa036bd882b0537927f39bfd731fc3aef1c414b9a94f8509c50c23542d9663a3d714de1552a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29a28e4b00b4451c7a23c6284283c65ebc1d99939c7ab5abba1d7f18a36f7a3921c41bb0573beda98aa3ffb465d8b3a2fe08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7d373034ac42da54baac65bf28c9087a1d8ae79e8580831177dc57a194d854874ea058f01add2cfc673518fbe9f94fe06bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd889d626f91c2b799a19b5f66de9d9a5701f482ca29f0f97c7efb8b70f934bfaa867cd5b90ad929dd1b0bc3cbc392844764b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5427f48ebd9e26ef3d1d3255ba1c6c5e47663155a03791c7765d21963a4f79d67c63cb42355f6eebc5807398ead709d9789c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4e21743dd243997b2d1e10f6790632a7d04154334cf6cc6cead5de5b84ae713799912d681832b8ff3dbf02689f02184ed4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a5e30f5a1046457223a74cc1803c7ddfcba920c1468b6ca382ec2125056293b7cc939479b551c67bbb992c0cea6ab63dc97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22fc80c0e0532b23de65af33964795e93ea04eb292491732c23e2d30f1eb628dda58834be5f66406543003da04a8c5fc991e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67414b602e5e520d3b0ca32ca206ca10aafcfca926814d5a6bb23fe029a71f36a2ba8711443bd826ec1902237e24bcf42ae9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf00f84b87a133e57b48519ecaa57c3f77eb7e3cae5a05b6868207bd2d04387244e2351fb777ef7ed4744996ba9aa293c4678;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc7df9d3b4c6cef550d1dfe4d06ee3b412dce8d2eee29ae6dd8eb39161aaf9eabbe8c12b6503c50f25a91fa8fe523868ee45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c5666914ac84430280930efbe3635ecf847641f4773773c7da2cd19cf2d96263374b6d6b3bb16044249ea09c5a3840983bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cfc978cda0e2d853345e029bcedf51a12de4d7f78d34f8def34f0e6cf29ea7601dc40a7fe087974c917d069dc77c952c6ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93e9dfc6c7273413eda9c817d3563d02e90a811190cf7acc4e498a39323cd13828e9c77ac7cf54d76d8addb0dbcae0891544;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccfdfade8cea3af8a1cfdaf484067b25fe0496086cabe2c52962e7046d12278034c144a51339ecd6e166ddd95d2439f385ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbd4d927bc3dcbad836134669e5befd6d3a20f59c8226a2160925158902b641d306c1929d983cdc6093e21da39ef7f44e19b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49e835bb6e85f5a7eb84e0fae2da24d2107cec7873297521885a60a5be699f82e66dc277ca0acd95e194d323e6dd0bc26e6d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbc919cbbe39cf389da9013170054a4d94af41305159219f7734f9d466420ae074739aa15edb04b5dd738a26c42e8d5ef85e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3496a63fd022b91b61b2dfb7edd9c838e61f275c74b7e9d3094b8279aac7894f314c6e588c6fc5198ae2e14f63a74045a35e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b905c2b4ab3f3466f0d5f892b0ccee93a11419a706306d7135e67bd75228c75ef1b656221a0cfc9fb0ee5da45f62a86f5ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28dc354dc7eaa9c3d41ff7a35751efd8c7c21581f87030735643a2565f8d2a1fa300e9b24fa11c34d12b49866d670fb37640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he33e7865a74fac66609c6efe9fa8f33a55b397d4ba6a0414363d487aa5361b4438a3424b378e10ffa9ea3fa4dc993c464f5d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb46fde2450019987808da7a1b7c828e1f9920011bf3fb0b251b8dba359895568dba84bb6192159e01b02426d90bb1d657aff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6ca087a014490b6d1f2c2ae06971191327183440a77d22f43262ac95858ce8fed8bd53c33a31c6c4bc0c4f47d6069a06162;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf834b7a0023fa58bb4fd5fb85c0932bdcd1c8911741a312c814b7158aacdf2da5ca71dd78691e46ea2356d8bcdf37155967d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h702d677bf6af94607da48e2b5e09e3c453f25c282d5f7370da85e455278d31c6ea8c1e4c97b362f81e979fd163896fa1dfa3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1b89024713c3578b0cf18089d8499799ef3f976e762e8b6279ea00d59ecd3cb7c46f61a1a8883afb17c7816557db1f35870;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7db297c45f2712446104be1df52ab635e2793ad06d9739624811a01293a9469e9d5c34ddfd7789fdf4dd8a250b42ea71c982;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe24e607a35e12b23cd5693bd5f0ca5b157e4110c7a6677c1bc3c6ef0062cf3f8d825416921af263e2592399e3ef22a82205;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e87f37103008b20ad52b01767a543662de472a8a95927044e50cd7420cf14051d3f351f2b8739031bc752bf9eaf9325281c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0431e15a4e083965f2a2ef207203706b545cf97f1c616ad4240c730566dfc77ca57f8048aaf1955d869e84739e916284cc2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3115c828345ed15485e8645b3ee46f99ccecb6a6235bb6ce560c66efd6ed475ea7ff41eb0c15b634ed66d0d7e4860606ce31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c747f27e5ef8d206d44dd77187f7aaed88f39ec652ac85b8bbc48dd225f982f9bc31439983b6b186f8eb0a6faa3ae691e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5597fda86de82592051336be9ec1d2f2b3face60f2909d08f255f38bf4237b0d17fb75727af1fd459b89748760d3c4abf122;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff66d37bed6e961a67185367c4c6b1088b991b4a5ee5fb8cbbf5ac73c14d6933a0caeedb72b889660a80e2542ca12f4e2710;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h499c79e05b1f86801e3b98036c24a173207fbc42b9e4f305c374744dc88edc29e01732163bb6cae6a6496f33c89d2020a5c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2ee0bb27800d9f1ee13721e34a6cfb65c7df3455594c59bb1c71eb0138468638546be7ced8e1fb4098ffa2cbc72766c720c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf51e7e781bac86ed1c84aebf05bcf0d0e4f75e134a46c4641fb3e1baa2fb6d61548eb86fd8c4105b2bb2b8b51489d1c881c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbb3fd8ea7613d4907589e85660b1a5809869d968078ec44b60faff8171dd2c4def3b38ccc193fe131501b557912f63d36f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fa56f4c2125b71714948193fd11afa41e50eeb06a18e1cb2fb7c641f58576160b33782c2e5cc328bf36c90747d6ee573407;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bbec9fcafd54fb390c64c3c34f260696deeebc835914344ac91ce72452805e9e5036b8d6e1ef98933f2448929f026b1ed86;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2751156b21e1f9e14eeac19ec07d8514ea729813c26e92d04f96708fa5eef0eec1aea46087c9f7d82f1c6897092cedd566f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f09f921aee6113c1669040cff2c2b64c5440e10483c97df2d6539f2e1e60cef2610f9ca19f7afbf4f02d48ab8060dca6546;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he66fb3a8887cbed74a7ddcf8b4bfc46f221944612d906cbfbd0856048bee3d832186f0810808e3b7ec04322dfec74c215e41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h154e4811e8c3db4f61aa9e983fbae73cbb21d1718c0e9566610fe3442a0add05cbf4143edfda702ca836ee8de4cf4d09bdb2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h808d271ae306f4d29b73ead9f08985ee75c4d9d2a81099f8d89fbafba4b46e0903c2c0c050c0d107697b5c8bd1ed017a072e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h879d687f66ad8bfffdc8eaf15066944dacee4df2ab0eb98596afa029640ccb70d33dc65b36abea11f316b1456ff08f1081cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70d7090b0e5cc0e44d19ed1985fa83d9b724a55ffa89ebe08f202783713caa901823f98fc9f82b9151f7cad90b2d45b8d7ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he229dca09fbf39eb8c2cd9619ba7e7fbc200bb0a26d0b9cd9634eac5f8cd26b54fae2d6d2732aef305f54d8b136aa910ab2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77d358ae96a40ecc4b84b96f0b6f0d2a58339409ac0e0e8d6bcc6716cb7716ad4c59ca3316c8763e9bbc2f7c0beb0971f67f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3571997365115229112cdd1eac3c2fd1eb93f74b5efe730b1f834aa672eb481c61eb7604092dac06e0160f935bdd68783e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57b520abf571cb4b5f383586cb11359436e5753e1e6d9440b1ac82d8f4ae8be146c3e7183af3cf5309b69068536f5a6de605;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49cb34769f208c2437254240c7f7254fb0aa2676448e4baf14002939f94f804f2d663f03413ec9059b9709435a858b0184ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb40a4fef7b9bcc1c8b98becb29109c9ef1cdaffc62d54e7f7018df47d82bf548f1e3a22c341b600b39b856a5c9b787e7eb3f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc865d5fa2c2742e278490beaca90daac7ae913bc76067ecd455fe156f3585cb0c05e4f359c9d28625c27b6f6f65bdfa3ed9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca914b1a70d7bc134394529c323276530d3dfaff6f12bd0a5d01187c68fccf3a0979e96c649e05646612fa5533b46368b5ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd0c72c68f6592a05eb3a2808de9a6f117c7e1809ef493f77175538c65f16a64e08bab9b7c00287ea2516a74fbbd3444d40e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc87dcd00df38756cd6cdac1f53ea88404806d21fb2252c66145616ebe360ee0ac1caad6a38eaf12fbb6fa7cd04f261abd9c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42a9d12ad8e02d52199fa34bcbf9a9dcf7189c501f6be67f246c797f7bb09bd59df7679666248e6da7dbdf15a5562570f321;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he90309f4009da0bf3b6eae7153522ae8e1bec9629095b34d2d92c44e662fe59122466dd0f0d599fbf3c3eabc595fdf1e86fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1caea91d9dea7a7c4be5a8396744f79c3f0de6fce426695b4367efbbe4ae915ba78a3b1081114b40ccf2bc3dbaebecde18e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7c02e376a32b79c2611a7dd9b724b2d5214003ae009a6940388463edfac9573702b1e4de02d07942e20fec4bcb6ef0089d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36e0a3b183eb68579c9b8c61ee754791baf82c9217ca3351f652be987065963829731375e895e73a164e13530b8c06144b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59f90554476c8ff9ea4ad8edc7c84c139262fd7b5b37e529e1a0a951b951e582e8b36c25e0e9151e29f75d6c7183d7f6bf0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c7d9b45fdaa4d4c82a6fc71af9fc1f5a3749f66c3332f72818566e79f6c7588ef7df8b09423a749022730b80893e7fe88ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcccbbe4812bc557a4dce40508416da954a22031cfdaf26d1bba688f4ba82f75d8dde8f2cf669e21513f30dea958cca2e8e78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2c7ff98ed4b7ceee516841de5c02f35bdf329d8c181c750e19557fb834319f575748a24e601c9f0f0d6845867d936ae1b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfed822ee359db408cb8ab55277b095e689935bdfdbb3787af4aa40828f23987f7c157ebd1cca429c5e7e798c85ca5074f85d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc617c97c531c73d74047b6579126c07ab1070b95f8ab6e09ea07aac5713268f2845c046dee29f3fb310b7f9242c2495d16f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b30627dacfaa0757d5f66a882110a305e7e6fa265cc000dc325b898e366418bb6cc14abff53158473664fb4422a32553b4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h183ff45399ff913c663c98ac7f8ec82fc82895a9ef3b32d0eeac05283d631984eac830959c0b05b410136222b99dd4b44bbd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heef8d5d5b5c9a429cc398d6c79950bd27972fae7715ed1c428375ef8ece4f3c39c3d5d815c0be7585941ac2acb926d879852;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h898c2d9f639fb7b92f01cbd76c1aa940bfac094465a9bff84afe549379c190d46ca1654685bb811bc1d67fd94d64fe44eae8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6d17d44815b173773f2030073b8d1e8e28a90f688430f48da0cee0fecb75222847cf9d85f3dc50c87e475043f18be5d464;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e6d56926179e3c8dd34b9cf1143c8f42af78c901e00ca5f5e47aafbca1767393fec5e01f77db1347b844aeced562f0538be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17f731810c6ffc897cee1850251e3278649ec0a70d6e1cea089fff0211f715ff44acbac2823601572d898aebcbe37a12aaec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9612299cdca88783c355f71dcafa57f9af10cb7a8df90de46561bf7f47757cb21f93a4efb2e4fb9c177c110c9c97022b9b39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab8d4d6038c879b504407cb960f5d842c22e2c16492ba71dd4cd365150199e21a1ebf8bc467a1a54e5e2a78500ba73ee9745;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h975dd245a6226140aee5071e9033ad5ac7396f65b816d218df74d2fbb09883a7888e9fadd7650701573858a74363c2e14e16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c3b1fd5bbc0f9f719c3ac48ac1627f765ef307ea8eef0c42ae40552a67ce98e05149a6d1031b17fbaa4f11494480f27c741;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26b2dd4255973e36e3e089c011c74f080006397fd9b347319e04ba56962ade0f6107c5b91555765ac6644f50e57b81968841;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h474e51f47acf1317cbe86e527474080262704bc9f5efc5018f14be7926836a4ab43b104efb9153ea597785a52ca70043f137;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'head6b13bf3838452527836db1b81fb433578954deae1d41ce86b4b638f07c24f10986c90fe4d354c1aa44ccdef73223eaaaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95b99a42e37ff6b4c8a39e3203d06c33f26cc74e36abbebceded7014f8d6f5db7a3ff754fae8e75259190bbad477bceb735b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12bfcda3797f76aeb6b1d6dce56351dcbcd183703eea2d16614bf8655280840829d65a8c8aec1c747f97cf206ea5ac0dfbfe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbeb21928eba41ddef9d1caac4b2fea7c673c019cd9b53c5285e4ba7c1d6679f847f38dbbf7e8caca980b403a7519eee7f30a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h274ef6d2355ab5c3f968767fb901153332443e5a6232e3954abf841371be152fdc5aef4a7e76e1353e3bb6a72094dfc1b0f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f9f228cdea5c145d71073998e8483b84c7afec21c563b8e2a6f27a6bb6e73e4644e1ce36672422374b412805d7279e351f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha082533b26870ef39a38177730aa24b21c2340beb0b7fc689e701095bfa09c3c1a16d7476347aa250a6bdd0e2c3df18abb91;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h611d70d6aff1158af211d014caf85987ee0e04d171c8c27ab0fb1f71e991f76dfbab8d0ad0463c4ae5021c335d24f553dd25;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10ef9f8ee9ea5e036c3bdbf6566df8b7ef8ea2e33971e65413d6a127cc159063858a129511df0a1ce1e07b5317d76741bcf2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c9351ed9963786b3a3b9629412698a878dd064ec71e3cb32865ccc8e341631c5a3d4d4f445e44696f645962af5eb60467bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1b90bb95dd9b70826a904f5ae2b40956d7d8095518d4fd028688674a7381a9bc409943b762d26745da2389bb5e0f4cf343c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82d0e5e00cc2e333ec5a41598de32cfdd62c024fe136e411b298e0c42a2c139b5982d0c4e45f27215b1fdffbcfdaec29de9f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcb34cd980ce55850a53145a5743cb0f19955a8e14f41468fd6c4269c2747a5005d2109523e3d783fda450f6bfb7e9a2726a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe5a975d46700d8b3aac658461374b05fab4b3497a93d89caef459b5d2cb4ea5803cc8e22fb0ae8ae9b5982ab15798edaa0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1645dd903ad1fb0e1249d48b1099c5481ff5451ffe0a20a1f3619b7bf16c595947d900a6524f30382270d7f38dd5caa2653c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6078d9b435ce3dc61e2b2e40f8db8bf1378d456a93437ecf0e3ce72eaac761399f113ab64fbaee9e6e27323fb7fe504275f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58905cfed6a0d567b7b8fb7a7718d9af5ee2e9953ed2d0d6046854a983e3e7bac497212c3fc1ff9cd49aeae808802717a90f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12759f0087a9670a2c5b3fc247dde061b45b64a976be134d19f9426e1a06787292287bb5e9227fb3020fa4d8dd3aef2a4023;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29eddcc012f9b8b78eed55275b359938a269c3cb88acf812d432f5db8d9a0a9e065e55682317d5985837c314dd3802a1f83e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd75008305d7d98af467108f6d1ae00a4f39e25ec28f04a970f0bcac34b293a88dcbd0c7565145c5f0dd7c6d6a91e3e6a3cd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6df783baa9f020cb88b1f6fa8e21b48117aefa3b1901416ef10e62b371fa1df16e62047095fde2472717773144e00871c64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7d9778da08c6f7a6242235dfb6095b345f96dc39981c84467a28e1b8f155494104c621fb2db692c113f4745471869b1bf24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16cf1173be8891650f8e68a4290b9f5cee1ff93313dce323fc1ad01bb2208bdaafd496a5d768e95a648d7d34762e0c0dfb71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8c676c025c565efacfd5cecf4ec341818da010f259739c919335cd50aa3c150e8e6fcbffd00221a5fb9531b00b5530ae77d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c17d51653ab57528acb7a86c2110a24b64e436684c84263d1c20bc31767d9bc3a1ccf2009c4bc1ae85c5a8f5794d9bd5bbe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9fd276021d9a81065629ec465a6d023dbfe37d15ae6104ea20fa74f7acfd1dfa7f9ebff43a25441ad557eae10433bc391d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h510db59cded16bef44d6766617f837f62ff4b659bba10abb64cfc559f36fde8d493d22625f2e00bdc424b0cb6958cf92e4d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h416fefa5a1c7f021cbea8c804719c0cc0418a8540cd93595cac64c5b26f0110e379529c1db71f04fcbb5746081db9df59f38;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d3d841cc8b0459bfd21b4a22020a272b202a2051ef8deb045a10e87cc410f436ecb0245d7c7ef768c212acaa6566536ea80;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1c875b2d7c4d61c028ace16dccdc7284043968440632a97c4ef72566a5f2795e85821aeaa3bd887df84703cc5c714e9ff66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f90609e76ec1c7fc311e55a1dae42c375097c4192ebea0368bc881bb7ada769819e9f552649b50df68c1c45e03f91813df0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9bb8f78cfc5dc51369668d6b3f0c597d71797e875b89506f8c00c3f74028bc7a8852aa0d11b6221dec3d16b7ab682867661;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7717f5e0a2874d48263849e5528e82dc386efb1b649443fdf5b5f515be02bceb504ec74b4a4477bdc9660e826aa64102c1b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf289ced8d6fa59dd8eade179bf1c85a57bb5fabb4cc4b08af1a587e80138831c1e713d1b594031ebee61536a69050a19754;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc491c4d322c95baade5ced29bc4104b166569e6b09c179e81fefc1d5a9f4fe6106d807f8b19a730626e3aa9f9052993bf03b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b607ce3458b8dbcf6383eda8034145c2fb27a9183c6280647cfd8da86862be8cd1c7c8c106ef037af61ab44b8c865b0814;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h997ed01395a6a547d3b7b17840e6d566c25c345d4e50143b13ecca217f3706774ae6b13fa0498e32ab626e74707c5dec6388;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64c976e423ca985d455fd12957e4c320ca1b81d8ee90b97b3fe2f7d5e1d5401549a4145849ff95b6952f061cfdc0eec1692f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89e5462136a49c9e9ae9bcb8fb494febacd790fb8cdb0424e220a644ef3e0e1d97a32cea7464c30c23e953dfc6ca5d34c2e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd934a4e4408dc64fd462882cff82488c80f070c1f60c574744127089396c42a43da59a2807bf1bfe28ce5ba0f29b3c96ff8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79a69855d62a91e0ca30d7d8dfb55c3fb214121fcb619ae3e7e9dd5c987ed9f7ab22b6254bae259b48a5a17a6c3621e99ea8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5231b6fbd2938d34cbd4b41f63b83e2eb475b8f8f9a2b60035dd4bb1cec9de79504372f9482c2c846e8d97c6538d8c317a15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65550872cee1ece0db03a0482f8c1e5f68f592bf7c1ed7c7f7b52b331bc1ac374c7ebdfe8393c3dfe3449ede5747ddb229ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bc7a41a807caa2ca539af322489f89222bc4ed06d30485bf562382f5a6683fc361aba5ec4e216b66716ee2476fd6bb5784;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc256f9edfab0d9fb152ef7de9781e6703f1a6e8fe345edccbe3f1a69e88c2e48a0b8cde5590024f16c88625fc2939b178e87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h787cc389208b789331f3fb06f706a903d7b929d62c4d745b570232a9da2efe4f66ca087cbc0627581724adb034ce679a194;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebcecd7876fa434cad13c1dfcd073b0cad04105f2603493f53f36baee3df3e1bf6926ab243f6d9b82b999d655e08df14189b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4317a1493ca28361977f70e3b8928881c02d6afaa410fa55192b2231d5657407a0656796860613545b6d3492d2d76cdc65ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7f7997caac08f9ddbc413d0e35864d0cfa996bca2fa75f8f04f8fbe3c2108318a107bfcfdb0692260255c8d00863ce2f606;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h791cb5e9732184cf25a4aa0d5cb5eb29a22647c8f6a54305ad2092ca5b73b2f1eefa321c5eb432baa1174fe638580540c84b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea22036badd837c0b2a4cbf9e2f0d8f9b41a3b77ed6689d220921df7976b28d53432ad62b965554495ab1477250276069a5c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfdb5fa81322a6c216bd7b3e4b6d0b23ae863c1e3346fa3168b23c73e2af86847021c783b75c6ae9bd21fda7a856e5389f0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5cce3376ed826fab1f501f5d4b761d0b2009d0d2f34b346ed39be746b346df4a23c5f3433069e10a56f36556b030a9068f25;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf05f837ab357707d9898918a3f16eb9f10b9007fc10e77f5175cc4c90e6cda6e78da25be5aa702de607de6d927b6de1a4c32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ae683f7e959cce99828dcbd19a8ce537825a18035e3d1a80efd24066a69bc9512c951d2d7a1adf85a6a047e1bbb089c06a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he39eb746119e6cdec3e9f8915f8f5e5910deaf2e196446b2f043ce7e8404fe36e0bc948a8664bc5f3244332dac8ac8ea67ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb91295b70ea2b79a9fcd2e648ecfa5dc8ae3a97c4e1356aaa40698a11d951eede03e64bfa21041a56f8e752bf371ed18b8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8e440dbffd94e1484d84563d7e6d6cb6f295e798a59594f26848f0400ab2bfa4da15f50b9bd86863b3172bace8f7bbe71d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14f6b91c41b3f97431c535a40e6739ca71bd2fb2f3f005d915a0f3055253a148332d1e2d6816387a5ee41e66e3382473fc8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67aef04cf3a0933f2d1c607646f913487e0ece4af230b31b9ae38279339f0c60cc464fd74d5c6c45621652a10a73bf26b6f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0035c45c9ac598cc907b19a2c3305b85286fb7081a0d8e4389ac5972321d8850d507b2df8e68cd0580090e756d107c546ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h915fd4aa59faef1eea72726e321bc6a8f190c70534144716c2f102eb211c43378ccdcb246a2028753829f13b9cffa1b1f832;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h962e498a893b9ad8dff917b030834b50801f15a1d077795deb782112bef1711987c15c0b0dfa4bba2c3d661be2f3e1c6aa8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b112083762975df4d006999d501419ac1f10aa37aaac444e1f5aed57ef0ed7fce2e4085570e2c950c2f631e2e7e87e8ff73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c91bdb0b256c5c50a11c4d4d5b570d0e4f6c495667d6f139c10509474ff79adb28f295076fcaff409f03b55e9be7cd46916;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b7fcc98a3958c5a69a2643c3b64efc9c4562a237d07903a077f3a69bd59a5d48094066e0cf5638ea36445ecb8fefc711fe6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87c01169a847fcf1a1c4ff2efa557cf57cb5dd9da6591bf6828b1091759a6ed0c19a2da67556896c99075390d8ce7e69613d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18d98eb4bde85e1ca459b2f5948ec313fccbe62994f8cd1743d188147fd4a3d69f5db55bd1fbab544128090fa4e9ded064e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1fe6112f01cc2550c5d36eafae47f70453cbd031543b9e129fd48c7c4d4889ef878d279dd992a87553e976a6a333843735c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52950c1a24fff25aa0c94b262ba4821f1ba69104bdfe5fefc55acdf54350c31060ed3fe19ffec705753b31bc1a7601e3076c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4ed2043c5a937d6c51cec25be105a17736d2d966e02978b57fa4caaffff6bfdb24c071831e916681a231ea8c9ae41376d81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59e742049124b27da983d040cc43cf8b3209cbace63311d5f1207e45ff99bae2d4f3bcb00828fdc518e73f680b236402b31f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb9ee6e76b2bf0c5ce6a686d7882a925e91f11c57f5b1a98d76f9c181ef339fb61cf6a833cd559bfaeda1e8520b93509b618;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25824c632fe86da9a3883b1244dd89ec59fb87c1ce5a16e86bf8ae8fcac9758017c0add48cbdab19fcb872efbed248da700e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8abc8b758baeebd3914b10d3d7a5ee199ef1e2fe72847ea433a984f359f046ee921e66fa1f171a4b812f343778a06e34f75b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4243473e162b2eeaf158c2b8d51db0eda06e6e50fa56a28c7a8f4c9e42ab94b54c40439de1301ed152c6c3f5172720aac51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2841e8eb0e6a5f48c75b4f13b73871f66e9b57100af64f57268ded4b31900bfae17cc253d3b716686e0f39a8b836dbc8578;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdae17c47171afedcd185aceccc9d044a3832fb32b66752149d52c7d2649e76cc968f11bd67381adce7440cbef960a09ebb94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc152d629a0113e1b5a2d49337d0a95b0b547facaecb21e72f299089c9248eee37601895ceb3e3eb368afae27f95094cfcaf6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69bd6eb9ff05b0e423ee096a08bf8facd5ca7fd6ed087cd0d769d52343f356275e03ab5f6de2d4a841d49c0c260dadca70aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66c06ab40e9a836fd0d57eeb34d4f82910619c5c8393c5ac43c4a547619ed583adb67d70eedf04c963883743e1a671f4527e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfda2fe95ebf59e0bab2acfa574499c8e97821597c2bb94ae35d99b9593342bb67ee428d46e950ed8e0d91ccadf985a6bb4f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3146b49108a86dfdcfde319938dcf291e72c15ace69bb47502ed2e98b4b6fd276da4d49d8864914570f3f2c0324261ca557f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5281b9b72c59ef9add583c4308e3d128ba797063e8328a0d3ae0032a41161f9c2093e510364643c40e069e6c1e13c749fdff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h471bf76e635db8a67043f917d8fce844082bccfc5bcebaebfa5e4393fef30b12cfbddc433457496861a3f9b762cbe704ad22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ff2772f5be745906218a1418260192e7a2d06a21966dab5984313c461b79f93cf6da9fcec2bb42f2c94bbd408ee8b7a5886;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98093bd20156f84c66dd7a1b6e1a4952f4584b00796db88a666b6323434984b0e97bd84a8dfa90365069813f869fc8df9218;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h936931cea711a8cab0df9bbc2a3681d915353f9a44970e9113cd7f9ec5b9c2a3bf95b26cc6f661bcb5a9bf6232ec6f3ba1ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf62d6e69370196c06c6f8f7ca308d0e6b2fdc30c715fa8ba6ce589c7234976893b0bd74c50c995310823a63228dc879f65c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0af077485f62c771edc166fbf68066bc8b5c49e09a85164c8cab52e6a546dd12838d8cf9ed2c6235aec720a0daf6f53c0e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf8ae35a71aa888e3f7249d0019115453405d95dcd752490907ff82114b11466401f901c7db23ca3544209f7f96835c230ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e795d75240d3a6f9d9077a5568c71b6dc45ed1c6d1676ef0ae10c29f4318a1fcdd8df7db26ff5de47632773005cec5934a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f851fb89c9277aef57925732697c557853ab699c0e53c0ac192a53e4b9e08e0e6e8dcc42022335faf3d4f5a60baefd1ccad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cc0529f8f4d818e252116a793873867857b68496d9ca7f8086d6e3ee1243ea26cc9e49cd2f7d710cd760cb18901a8a5f992;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9df2799174e5e8d5409dbad5cff8f7f89e059d17b8bff91b90cede8f046747a228fcb89539714f772d70f1e32d71edc9b4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4ffa4936f691288affe50d20351d7f537161781cda5e36a5591d2e40b85ae5cb6ce0393fcc560280e6dbbc64c6585fa0d9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ff38c6d3f0f7c5086991ed1f4ebc61c517c13db804b32dd99025158a9d12752e2a31c4ed5db4800567b8c46f08418deb734;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4490cd007b31ac47e6076aea57f7d3dafa7477b9aed592772bf9005e12cd5da27969bf072b74c2850be77edf13f5b99b05fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76999b61de0a8c639ef44e03a4b22513804e3a7d1d97df76f01ee6f22a15d69862cfd27040f4c19b7458e2b6272b85cb030e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6efddf88d2943f4aeb0e9b61d524b47f19c665bc2d53c0a06bf39ce206ddecb37c94bd868936007e2f6bfaf5604e6257ff98;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0732a3ed63b8fcebaa00f3a013460d0133c0df8b91b77ad7d0e62a166e6c6a271c5f1e842ea1570dec084b20e0b2e77e19d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf044369d96b33a6557d72305053fd64d4afc8cde82e3774746dfa2e611f029d39e58362e961e70a1466f711b251ebaa8341c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf63480d9d7a508e69a1c474024b9e63811cd01ca2d2207d80b161ceb82ce0101335501b256d945d6e011a5ffaf15c47a4192;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f8d3e242bc53b1778d1a72b5441a3097b58de3d682192c9f9bda91a699b625038f4f9c7c9ed9fcff9ce1d1c654e57101b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21533a5a45b4455aeb744f4c415f75195762c49605096235866d04b8996877f2318bcf77f3da648d41d7e9c963a6c40e078a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h694397790788a2c4477a3042dcffef9ee1b74780dc8180cd7f93b448926e2cc9a03d6d9ba12725d28e28d277037f078f87a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd84826900e07e5eef259296e4e2a50feb4c9809aedf5330018906ac53635f4a3af940d9455e59593cc6ba011408871e30959;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72ef4e263e69cbcee98054e7eac70dc94d3c495c66080e950605ad14be8fdba7fe3f4484928d47b7cee83c5fd32e2b2a107c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3e0c2db40dd607e2f670a61eb4674aef6ba2fcae2774df2f2090b39e2032098b45e9725245e47324485b76c14fec5a456b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68d8e93be9c931ced4188c85fc577dcbf713160841a703a0b0fec0eb717cc05924a9eabfdd99383cf65bb4fb0f9dfd7cb7ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dab1b1749d12e079282906f16104c503b68c52c45db5dd85a1d8223abe060b1355283a158ebc0599e8bf8b7844d8f60b5c1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h718ad1f71a31d5447555bb2b6971f449d6c26fb43644e0fd73b1ecc4bd37153f2d2a3b1624882e4dc4cef28cfa4877b22ba1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e3a26f781773a48bed42b6c7ceba322113e8d7264cad9c3ad760b2688bde47faff73784a909b24211b6fcc9039e186da0fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2026cd8438e1e2024bf557a2e11779b136051650018853a4053fe019f7dabfbf652722c26c9d59c7aa8263757208858c1d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b565eee82a4e280265db4daa48b0e340db4126c27dfc6ec06caf24e68099025fb2e34523184be2b13eef833d6881a77ea8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h725127869cb22962d8d8a676747a431ed374bc925cb5b538fc1ecc45d0fac7b480bdddba454a98af3af4c18bd3c92783701e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a0e15fbc422873ad982e895e89151e854893b4be46dd4643a4d00cab5ee1a71285030f71996da317770d748f2a62241117f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff2a866f22f534796917a3e558a681268d205209aa29eb0d45f612120eaabc3164fab09b514e3fc8ff500cea83b0165185c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99f6402ce3705d09a303c9edb6d9d570dac4741ee930524e0ead1dc5c0fd4d68e7057ea2a6cc653610cd545e210cf202fcfb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d600eb70418f9fc47f0a43c785171698e364536cb9fad82cad9841e1767c750c52ac51decc8d1c8c7571c188af36ae040b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79401dbf0b5f1201f963ba88876f7b19a6744126c6fe86044ecc3a3d574c1a88fc1ec2b724f9067572f1e232c941e857b08e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57adce3faafece514e0b53a1bde8282eb4efe92cbda63ff039ffc5747c87b6ed8b74d60d425e317f2a8f764110187facb734;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b643ef6209aa6527b8ccb05093c16815872ed55665e9817f42ba4121ec54eeb4bea58e339930835c2b40cb234cd175d054;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfef9f1fbf7d1d1d34c0745eb31f6317d55789aece3a946e81695ef4e6880fc1b4f200fb37b53bc2c0cf70d00ceb3396e4692;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26880c631880915f545e8dea9909b3cb2b7e6bcba7415fb38cb39a00f084855d378fb6934d032468eb4bea3ab3c0eee412f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78d7ae95690ae9a132c4331d9c8f99363e5b4c80d62e39013f2b73e8ebb54867a8ab857d152cf5d821c311c89906d2c1a05c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02962a93e54233313045226eb1208d25637b4e26410cc4e37178e0c4cbdb3921c88ba2dd317d58fd8f73a20683b5abe5569;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde55dc61a896e283fb24fddcbdc2bac27d8b7280eb078eb00cf211f3ed7b099e38554151d63c3a4cf9b9a175b749b2a88562;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4a0f99ccf764dc78d6ed4fd3c40338e6797e01028fec369b2099f810582496dd626519ca63d96dadb885d613fc7cc7630f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he32fa4de62149ae161683ac777ab68e1eb6596889908ec95d451a8fc0ab2be4f7f4e99d54f5567b8327f87d3572022cbe305;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88b189b89f47372d253153b5adcf6913d82b96194d97b19bb53a6be05906449fe21ede2ece95264c0a38b6927af176457159;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d1dac014a63fab94a13612ced8bfc16b60a15edb9aeb5bf3fde70924c108e234b24c025a035622bf7d92828594399185481;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b2c9cb24e449c5a4d63e85f8ef4d0e7b5f1b10ae7af28cecfc2d5333b39966428a83d6aa7c99614f3363406a3059fb5d4af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed1403e15d41e93207dc18e9023890c69c02ac72585ed3e049ad04e235b50d741992db65c0451d3b1a1312d0d461146061f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98fbf08877e5d13f84d640097f6b5c67aeab127686efb6c05bf47e3fba05ec18988f8354bf0c4bea47b9bbb0b957d7ba507b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7c368ffa1ccceec085246d1700023d4774eb4e1b72df53ff38171b23f44d45c4220c0bdef0234e16a7d2e1b58d30eeebe5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15538efc9209048f0273ffe14c6ea3b848b0c65f57163ed73db113d23bfc24006fdb03c3339d0ce52e2037102117d5065e0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e62bdc38cf31d15db33cfde0d9e5aa61c9cb096502cb2edd59894d5effe60bdc0b71b6bd92d1a4a82f7bbd377b357683c85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbfee06e69122a7de45af7200f0efd53c6dc6377e6d7e7fdd57cc94a0370abaf32c7245f6290467e37571c028a0697e21239;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb23ed5354ca2057b11286c273c4f0c5d7f6842d302ef9ab2d3df457ca2607cea2ba06c81232b68327f9bc4ecc11fc9fe43cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73cd5178b9120dd86ebb916cc167bb320a5e001721d3945e14fd4e3b5d22dbbdb52ed64c1c1f4aaa629f8b2c54dc20199ac7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8eab283f96040bbb6f3850db04cadfc4f051bc1168f01ccf0ceee1ef8db48f9ce2cb0adfd812f07631e95c768f484062b8bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cbe749a0973e493fe54d9957148b12d7e52a449bd36d594d560d8b4b15e3ac22b8e83c060cf0562a11efc3b4440c9238f8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h825bff11aaa3daee5ba802d9e268e3a11084e6baab6a3de73305fc35a05f05b90785ae7e4bb97cc4c53f4bc949a3e153d993;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86691795e50b645c44d26e2821ec895cb3389cbe3f967fae7c80be74d466ff7b5d71d074d4da6cdfeb7485d3ad3984fe8aeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b79c60f7e0a46ec7630d7541328592b49f75465f25e3879f376dd944cb69949aca97a7a9b41e1f89104e5ed0e4b4520a4e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69688bcb50786d71a2d85d23fbe46a6d47fdb686225e78d9795d9737aeb414a2b7eaa9d98b65fbb5ceab30ca8af80925c3b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h641a033592749d11317bf45f7fd1dde5b19633dab41937a9c90e660d52c4b8a2ae55a1cc40b18d7aa923fa8b7e451cc36295;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee7bb47191f32c937fab0adb88f1370e38e0fbb977b381f5fa625f31a131e0075c2d315454f491ac57861c0de5ab56cad882;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9955d96206ee2ed09936e0bbb720a9388d7927490467707dc9503c6c3845c367411e90b93e519106d06025add65fa9a40af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89624d29c275c7a58ead166bb4522736cd48b570b98db8322ed4de3190374e0c006ecde19c62fd9fa1b25e452e8663bacadb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3067238b72249549761ee1689da0b6780f7c251c5d980df4ea70e7a05a79197a66739fc164862b2808e037f593a61bf65b7b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7446282c352229b46ea4778f879c09c0f4643202877c74abe475dfbf9068cdd3b0ce9ab7ee08ad57c8a07b0181ec7e5d7a16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf223f554ae8cc3e6d3fa89f3f9306163890c2960eb6183289dcc2df7eee0669f33d5b92f7c6577d0ad2b8e802be906faead;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he845935017d0f741c767a3281fe518620e561486048295e8f87bfdcff7499fd176dca5e32c0c6421074697c4895cb5fe31d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf8462f57c8abe44ab87653110a2849a9038a13da33b9f2f7679c1419cf18e9a305026982eb8fd2bf5f114f2c6ddcd365fa9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f235dda3b2a0008b4e5dcf8af7faf326079bf729a2ca1155e8e1ea9683a884f66995384ab7e45fc7570f8e8196e7efd56c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed23103cc89ddb90b892b64aa1955944a7a363c8fd38d740f2e029b5157f8b87b06f3ad2afba2d7aa5ae83430a05967011a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c5f6dcfb6c6a50abdffbd8b99b3f1110de2452ef8ee3b1f6e866c7a07625bf6a115fd4eeef18b3ea57d0fd97f10e8aa7903;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7382455c725bf29905b7f937bd2dc0759804c60b7d52e7358ba0966cdafeeb9a032ebbb70f0334a3194ca5498222fc26914;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41fde4ffe8f4a859ea57e324b6232456ff30386c7ae9e03eb6db821947ce6a12c98cc0bd3ced2f05dfabdccc054f9f58a90d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf97f00a095d41eced68f6adbdb3a0b7543bffb0c068ef345e268ad8d04fa164efc00d79689778198e4fa62c2a5291f7013c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a33dec22d81a46d18036917c84ab92b042563431ca8bb6d75c3f94acd40e97a0026a795351c7dd5537daf2bdab45faf9391;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf00c8cb7f729fd4cea270a51f2a5c52c0efdbaa511859ddadac8f4b354e4e98548bf875505c93de3adb4b6f9aa21ead143d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha46fd110e455b0c7e27cd795eba5cf5a5abdcb243afb83fbd16a26bb3269831938c57581974aa4ea0dbe31d630cba8a23b83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h871daddc40659110b16c4a0dd42bb566697ebab1e7f91f1903d91976c28fd5fed35bec0ed3b77fbf50dff9ea522d23b90483;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha15a4010b94e5f31f26f4c19a69faddae8320629098b162be599ee77c37f04e7c949e6cf0cac21968c8efa9865a3042eb632;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbaf33bbd2519eabe99d9f02ef3a474aae3b7b7944ba8b40e492b2de755e80366f30292fd99942a7f585c9f02b8d58d3566cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b09f9176d1c3e083b68ba12c493cdb4cbbf011cc04a12d31a159ed2528ef6d9f6676544366b07c9ade16c82e19529b8ebb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c831e13bc4f7a030eff06c587d686b8a9e6f20da6d5213204a4c40c925daf04ba7f4f77de33dfb524d676d7be558f13ff9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70e30e0e1dd7db85723c2903c8600e92d96c84b9ef21f99f0745d6dc12737146d3d2b345ac18c28bdbc8d3dc2b396e23e06f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3db39ec8489a8f7320e192a7dbeebd428a5384e5f5c7284552475b8be48f4f0d5518dc36e58a80ce94ef2ff373bd6772d791;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90c40952d2965bba1302cef6bd18b143ec4ba9c07754dc4790fcad8a57f98c14bcae37e5560d835d42e7dd4fadf148196a55;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7100576e9b3c6e386a7306c2ebd82466a39344e243d26d6029c1236713429045cc2cb8a861242f50ab97cad6d65565bec17c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he88ff9833a06c436d964e261579dd644692b398b129ad48824884a8e3da849bac4defffa92820da84576bf2bee1097cd82c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3519daddb2e81d01cfb20dcc733a0567c6abce69d5ec05661bae638c2bd5a097706111c31ceb663e672f96564820849b322;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h676cbaa95289a3714239f6c059bb8ec6185ba0b7bbacd4c06420dcaf25ba47ad8899ac8dbad43b982c7e509ccfd76eecf8d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcadeb3da5b397f7eec471db3a036da336510649e0085d0e192527e1b8d812657d59a0eff89b16187ee7e17c44f289bd22e91;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf03ba755f2faaf2827f950a849950a3aa03e7af9486a811e9b4a11ebe65e59016b026934ec73f916a9ae19f5b77e0e0d4e9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h941733e169000bb87cd8a8fad4a99eeebc9c3eb4eb61690767717bb9dc2a12f9041d589b650996db3f5863b36764de849d24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he97056d989966a7f9923ea50aca90ba105b2394edd6d54e5645e80d1a61727489047049bf8c2400a90052c56442b3330c0b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55e0a046e7451ecb996beaa48a0716a68d2269850c180f72daffd0d2d101fac0d3f65f6a3c50bdabf9333c54aa8b41fa28aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89897e8a5636f829cabc7a88ed26b2d5b5fc3222543afee658a2db63c0d5d1c094a738cfb70ff63cef141c3bec0916ee4d31;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9baf2177b65dc5585f3b786e704ec8ad167fab1f3b5318d65ec7d46ccc27bdd946f956fbdba803ac63ff318fe1cea690b02c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5af9021eaff05150b04033eddcc1681fe8d109a30629bf689d85d56b6087d66f190c38de10f61bfdfcce17825776140498dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc8a68592b7c62340d47c778bd2f9ba5b729070715a8c69062182ae2c906c93ef13b829cc14c68e1c20c1de6757812ec37ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4e047a59587de92b5a101422170985d636eba12ad40b29657850925fae572e1005170e2649ce0559155b88fe7b7c718ca2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha53081136a3b7eb4af3e2bbc36302f3fdb970d3ce167082a61c63672be0cb45c8a11b8f742230e649028a4a8e1ef161e6a42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa91515a53c5118378e643450f540464b49be992e1d95e89654fe78a9a0c342fa4c8e8d49a3eb12679e6b2d77b80d7b2c9c1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8849994889220d74a1e1522ea1395140dc3b15dbd94053808d66c42e5d79259aa8d93e460f6a9169d70a8de3421f20c26d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h972bcddf335ff903bccda52d115272c66122e7ee421dbfc0201984daaf4df568cc1bfb8863b2263654d548b7eb0ada304906;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa4c4837e1e67191c68c1e98c7405cf112ac27f2af7111b42b39d16882350c2282a541a50e380610855667ce28635b839ec8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd085efc8ef18e52054ccd63ec5aedcffaab63010efcd258a8e6f46737edc4c16fb06fd405b9a6e2ce36bd4fa946738445a69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c7bf42eab79d1b1b425baf9f4f333ac4c175a941e413e2313dd4a639d109bd3ed73ee3fdeadec65e343aa6119591b247363;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4e1e232ba3c2e3dcf003a13523d85c2f56ad200016344ce3368224d931c3ab5051d10fbc341899cd08e4dc67b9c29234f77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc653ff11bf9d53f32d2a1390bef73d5bf7a4e5c34b4b0da59633250e0aac6c862c28391138d938f5c4a56a8da25031ae8cde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7e5f55d98642f80bceca56270acaa061eb5675fd69ec7427bb5a4b1be0db81981be0b9d94b231d49d6f82ae5e4aa3587580;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2beccc6682b7279b56447222715ca812dfbeb834ea538627d8d526626dbcb08e8fc10fca562d002317bdd38928dc5af27bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92ce8a97c06c4a006c52fbc3f6081c04ed240cfc125a9f97fa1d8dcdd40db5c4539204be9eb7f19369b9629efd3263baaf9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h265de6ee47774babf39f4de3a0392a08cd0a67ccbff3e8c834a890eff9de6b8cedaae80a8519c8980431c2870eb2b15a324d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3a2c4750371cdd13cefb33535de3586ddc2b554d63c077b12087fb9bbc6590e936f7899d61f8d22538cd97086b3e3f86a3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4c3b7687256459820671d810025ec19101f39c48dc45f338cf6541c3bb01cc3ae5b74e72838d2ecae5425d3f835311d5fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76441de92fac7dc222f6b12ff513a8ffa88abd1f19700935908be48a177368540532907390a64b95b5a5268eafeffce93d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12fb60bbcb90ca8ccaffe9b311090cb916821e30133e1db65c3a3a90d2bc75884298c4827e4a9c49cc6efb2a87e83387e8ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fdf92636501a70ea8ac2875cde86cbc5329e6a55a5e54a9d34adbf27210e3ae0f410041a7ef0749162a61b735a8db3a9e0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ad88726bb13a9308c0c316c33ecf982230130529b7dd9e3c2119a5cb537ddc15fdaa107b85ebc7392336c1b9c93c0bb57c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ea591ca44fe29569e522c932e4c4805c2a5e0f07891a37c645fe35ca9fd02c843a784e0c736918a22ec6f5b678987d92e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h666362ef4361cd1c1610e1f0ba403de4f0273a7537beaad7f9bb7dbfda9e9a20750073481d5ddf31703813ef1f411550d340;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h894a7a891c11e389ce245ce75570ec0249657d315beda791422b1befffb43bc663d623f8f6049f33678b2c968734245594b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb3a0eda47d3ef41eac207f6464b7855e6a39ab04aa1287ff3f227895c83579abf1b269b91ef39d8154cf0755ba56c78f2ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d86021d30447041b4bac5b144f4ad70d2719689da00fe33edb0d8d00e4fa88712ae5e3af9be9e037ee6a54eaefb3d028a66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1da301fa0bc48ed794fab6f0f483add50683094051d2f4b14530836b455d961ea8665a9e89ab3d2794ba6c15a5d10b7c990e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8dc099e9f5845a68a3c5c8f03ad08d6a81419b417b62369bbf339bc6018aa299955d976d0cb92ede7c157cc242b557e7a23;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84c3ddad85f28f7e7b51dcfaab590c0b1b4e1a3d95428e4ae888bfdc99badbc2b3573f73a876d0c61070e98e5dc836e760c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdf6aa0537711fc442b264ae4fcef5107440010d5a7e254e07cb6511dbb6fba5590dfb72c9f41976492f01e87e0c4ab4431e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5c99ec262a7354ad304d83f7d8994ff6f47c2ee1aa3973157f972a50298406b9d9919e459e99b9fa2850de1f63b2348db59;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7657ac62443396d82b635a40d719c6b9ce16d272552f2edb4c98a26f4689b06451d5eb2d4fcce8da7a1a877aac20c5728cac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h232d808a3c70ea0b85a3ec9a6d137360e69b63b7f42de2d9fe02e37b2af35d222e65b88402e00d3c3a1bda2f6a7566265c62;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71f941da7a06576a2a083c4ba62a111bc118236b0a4f194dba51d8f1831ec0c0deb8079be6b414be7435c898634dd7a1021a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43b9f797a29dfa5c0e2817d61082f15fed6e50a034a4e661e4df5223df8d45b561535bbb442b9208dcdad74ebf1b34be5567;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce5bfee0499a888830cef3d4473b58f87a514df7cf017518b6c4051468f8f4f3e05d545ddf1466cadae7c0c1970778f49768;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3993f767d0d4a6a4300368abc8385abd3600d0baa636c42721f2932bb69320bc147d0d0d7cdc4253c92c8db6cfdec52f48b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae0821ea48ae79076feb5793ec80d37a3d330e8ff69a5d116c2be67e98116807e2d2e53fb6524b7e13f1da23af4a170f98e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44dbf28dd9136e7d95057b2dc90bf1c5b3bcd29209eb93b336f8ea8d97fb93e3d211f0bebda97638e563134ce990aeddbdd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ac87b922b86dafc56de04b98d87da97946e1e3e966542a73c78a755825a2789d3abc546f552b12fecc023a16423ed74314e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29c4b478fef2469308bb8cf8a6e72b823f4150f8f2c50c7ce530fc061ed2e5727f9e9e531fb1dd1d8493135ab1de07587b3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha18a75ca5ed1aff4b7218efc9efbaf7cc2098d7a748bd00463cb7ca856510393d43b91deccdf9f5b83b8c85c0887845d06a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a4cd025c83dbe82cb92ae14b1e369c183064fb65f72e7748388cde2cccf606fc70ce08517455879151481cd6bc51f423574;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h555214954a1cc11b3fea27fde5448b4e5efc1cb90a176ac65cb1b5d3288f5c867805609b80b6995b5bafa6142c687b65c593;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had0a352269a288392ecb76bcb817a4c9949d263204764f584f3dee5c0379869b6a97cd1a756d0fbf849bd220174c50b57c7f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cba871ee9122818432b8d8b9ff0bf971e1456ad99894438b84e8a6d6a07c81c9e3140ae09519db694ffe65f89d31e994f24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ca5eabe9a62dd1d1f2d0e5dedee1b4a7e5f619627899cb32c549d494a3ef3cd22150a2ba9591b57c39d3b3bbb19a080bb2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7231db0137ee14eaec31f4c1ee6810c193a383c1df87bf73e852eeae45bca6aadb0fc166509c04732eea06bdb651de7b5f08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a0c314cc5216377b025051c8b98512eef11e3bed2df7b8bd566e340462dd807c52ea775006e42081c8b1bd8e5f79748ba5c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h933062fbb9343405dfcd4931ec2147e5c87602fd53671719bfa5813ab3517af7366a52fa7a618de81293a85fff03e8ca157a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ef178a3db626775b9c916f94fc8edad2e43fd37b86c8d725d8c2cca9fbdb8313e98c3db68ce6c8e07ec8c91aaf9d6cf25be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h316bf77c57059bee2a2c6eb0c22f2a4295ebc3e5f3dc371fb522fb5f7dfa322d3510dd9bf17a92338f70ea9cd5f584b0a32f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70716fd44b756d2c94220ec22220999feb7bc61129d96a270e2648c6e50cd261a9b2f801975a9626e8df720c28f1f7f6d9b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1760826f23d88bb3a24876a10799294ced988d9a7daf3da1c93395717d3945953f6233e1a9a817ecccf9d1435f5a2700cca9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4938a755704941d52b3abafa5c5471239d26ef01b22b7e893142645005261095025c15c37612ab8f6c2aa49953e44bc67de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h835e55e6012a0588a398fdf01259d35ebf26f73dfbeb6b82cf1014564fa17ab55030f43c355425805e2c384f70bc94c0ae00;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf95a149f4e2efccd4b5b2ed36a8d6f3fc376976f75aa72b7173b51ad40a2ab5b20766dac9242f75c77fa3089b10507753477;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha703c859651ccac12fe59cbdbb5545f5ee51d7cb372766e479c4efc08cfd81121445f6bdd0321baafc2bc7c64004f3acdf8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h339e874c03ca38b3f62e960406b68b608dbbb234e94f857f4abe2e51d23a873b426377eda64ddebef939427576aa0e74ad32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48499fa90435f06139e6e92f676f4c6b7f2e098fd608d3b367745b632a48ac9b04991cb7f95d92d7e9cc553505e284ef7e01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h283d168348b39db1154e3c49bcd201dc09cee9de5fcc0d22242c0a30b74bd765af07852f63c480b7e6d1f3d2bad6e979680e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb97eb34c5df1b956ca95723400a062f42802b6a4d3eff1de5f325278532972c50f2323b4283d8f6820067e0945096d72448d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fc9c001db4d4249cb895397fb4b4f4ff08020a93149fb8cfa4c8d8dd5425fa65ef18337c17a17ae0d5cbd1693ff8541a0cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6b2b2ae2b85989c4a11db979bc53b2ddc94e8c8909dec501b419684d5df5c871d440cf11db201a331f4ce09b4f5201f8653;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2247582af58d692cfc538ea12c0942c802f1f7c343d01938f0d1856c0f4909eb2f8df8d16e9f8429bb60fc7b11cf6fac779c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe7f571224b5b3ad676bb188716f1ffdda331788333d1debb75f5430f81abda0ef6cdf68c06abfcbbd317f42548a322fe241;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f2246dc45654f785565b59c83d5c47595a8202a177261062dba7c794d649b24c224714377727422eeb1fb242b82508367af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3bb5d3f59fa5c0a460ac254b3478f387d3a924084a6a5219096270540c695eeb96f2ad1153a9d59af9fe89132622cdacb63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb43953b71dc7b6b3b60fe4a0146b97e06e8b59e75b95bbdca18de0af96abd42800214747498f64e5481a1d7b9060f661cfef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hace24003af630b3d7d414741e6e7a28c64362c4a3956c092fa4386cdcd7b11ee02eb963481c2363019c53ef1f2266df42f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdf5b06ef8bf7c0cc5863dbceeb326a362912cb20be7716214bb7a663bb43b1b591e007d422ff3d47b5e5c8521aae4422f9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16c5ad328c0bdc8ea17fd07ccc587d1ad7a01edfb0cda9ca9d336979f1673c67ead1b008a8f1d2e832d81aeeb32e4d346da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48fcd04b1d087f3b0a0032636106a17737d19d8df5d6fa52feb2b117b55f5139315e76e13490204b7d2b183bf2154f0ca8ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdeb2f53c8759b58dde38c11207760ac841b91b63266dcfea36809ddce95e8924d4d1a7acd36cdecbc8b8bb1a29695ebb43cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75daac80dc331db998bef1384173312dcce5a9756024208c2e5466c84a9d2c93a94d6c285959157e6c0f1787e1ff7d7ca116;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbac03c706a869bc46f2c5b4b9857f1b1e716d98af223515d452923cf2f72511709a8fc54f2912002745ad00883336c8b0089;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b2c37853a9a94470b20fcd120f99972162e7847d4c38f6e9d17fe1196006be7d0e579ca20cad0e73a97d14e5a0826fa5221;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1f967aef26ec6153ac885938d17866e4c5d4f8a7209a4cd8ee3cb3855e5350c42eda6af515ecf71e4df007e1432c58c3ce5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0f8f5efd4b8f72df828683c6d364dc311c4c91fbb51d8b73d955904f4f7474db890a32dbe1454907ea95ae0d28b502278d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6d3026a10919e4a4e622f4c40fd82d10b2354ef36b80e6b725c7e250e89be7056b606aa35a37463bfb206746f041eb9bf81;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he702aece9a911d18813c7f35b9db62df43ca350eb4a63df34db25f3fe1f89b2917bef6885c987b42dfa5ef4ba63d27b2399b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h168d159d6316b3538e9a66e7313230571201188ce5f45d72f1f164a038ce6e1c62e1a539f756b685adf6fc99c6f4da12ebc6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1962ad78dccc3c73886f54718977f882b4cccf9fd221e73e7efaf6dadb1a18c1de775e0ac33f275d70a9a21bf3931f556e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96b33b25e411555e1b646c8fdae4ac74176878e4cb78c24a6cb128128e3c3df982ffe002b58e2943d2cbd474730a32bfc24b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde7174a99c20389e4a0d067dcc424310dcf8117ebac9996bdb58f9867985c0d40c6d0c3d0098f8bf8165af33108929d95e7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb35377021bdb4cf35c11cd1542b3c572b5e128a8a3ecc83515fca82e33f5f54c46c90baa84c780ec7598aed8a5951a21cea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he721c82695d1fed91227acb48efa0b2bf429282ceb7e23717ee3a8d4553beb4b10ca31b1e4645a939e12cfe3f61a82c54ab0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h444c42e797854630f1cc52db068355b7909c4a8159445f63663b6cad2c16730e3a7196759cb59750601f941a7db994a342ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7ffc3b255be5419961829b1204c46dd76944825974d267b08ab62a9c8a5553c62ca575fb013381bd8958d2059d8f1334784;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haaaeb64388ab392a614be90e52a44671d2368cd514bed27381bc8b62813b7b7797a7b5d7f65c8b58a3a57d9253204a042e6c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87758351f3a05616720a2f6e2f177215e70b6931e9cd18165db2c305608cb60520fb3580ae27dfd088d6b03a4c03116eb560;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc65c8b04d4924d8e30ab3e6079fda3af7505e131db5bdd313d51e13e90dd910bb377e906f926426a7bbe74207ee8536d02a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d4ca9b3929300586675b1b0532bfe41f9ccd39fcee2160bc3aecfd7c72eb1fc194e79864bcc412b281743b5ca126dc7e87c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cca5af9d1a2c4e2b366d5775516fb1b958cb5ad05b883e215febda5a774e692446b70a694324eb49aafd94aa28d59da2ad7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde208afeedb99a18887dd143c4d1f9573d7146fe146fa86518c8b39512271516220771c0fc608f746d5734be9f84367e74f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94f149b72b9b3d68a42a0048e11edd1d259536361477ef20140955360b08fd7d029a88d885a249ae1e7688bc6bc94040bb72;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec42b71ad6e9f555ac53c721b69d3f28c2e9101b1fc6476ab647fb013628854247e6e052bf95a1a2eab1670a99d2fac71b94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7dcfe512bdd7f6d04b4aa31f1f4641559188bf63de1215587b1b39a704df3fbafc446c4404bdf476c781dbc10795b4be4f73;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had855b9a713aa42730d90449c5c8b1d78e2c75000099c4e4b8d0bba74ad48c3519f23099e9ea2f35c3fbd631ae3fec7ee753;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb69de8a17163bca7dfef719c6db94325a90526dc9a8d6de33adde5142df544d8dbdea00b2e2e74532291696178690ed39e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb762e9d95060e39b03e57f20500cbc0de2e38336708176c3a3ccac6e5b82b804f431de824edfe1d820f094d22e39bd2552b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5f04410df44546982921454e432b7105ab25d8cff7a2760c09817546884ef1e431b26fbf96ed63ef962925d520e6c57e66c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h608b25c20e879ce78583872722265eca65df8c70554b9f9ad0b8c564f7b40c909c2eee1f8a16d4d0558ed6e0c17b111b4c4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd883b323137f1bdea12d62bc61bef83c4df599b8504d6d9524a0a1ecc85b39d3533be04362aa4a4ab6b73a7596c7aea8213d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6cfc4fa391e44f75d3344a52760f9e0bdbdc7aa799ae2f0e7705766b5c29aef522f04319a2634524e4a9c0ab04de419ce24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb4ffd54ed5b283daba8582a141425083e9d84585d19520ad52aa72f814d3e473aa23ce4795245b156278214c176247c3576;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1720fde3b0c3196241ecc7248bae4cf361e8503ad01f76cc6d6029cc5519bae4507006bad6db756f6cdbce7940f3b5a7037f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57ea9ab508d18ca8964fe2048920702e4607965a6717a09419244dd086ee21f0474325cc6f6273435b020c31ac27e65cf689;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4e2fc34ebf340d6da61031d723c954e48f4885ee761e751ef46b0afb1d95e161a3e5ce394e1483962ebe95ca8af6dd6fffe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf898aa6ee19c249faf214b2548c13bca87a356de2f22424dbefc27d29999a06be64bae9b943c04a28016f00e7e7a0320b0ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8fc7ca80f907ef434c86810e0a2961973a3f6ce658b5ea9a52499271f90ef8c2387c3534af3f5fed24f8453856c4b0467b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f92f48950e54da906620e02e2fc828d5c85997e8970b876b9c40a1ee6151c378da9c621f449287648080f104f35b0015cc6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd91494db4984a203ccbf855048592f73f7f365f4b74a75b4357e572f6430548c8538882392b78c51a9d2772a5e5642d873d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4f0d4d414d5a6e92c1080ff25030be16030e8d4198165791055f6779d3ae859849f02c6e4aaa1a104757bbe150bff234b68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fd510f3741def1d5438d4e665e4bc86906fb990808ad47a26135699a2322e15e177fbfd5d507a5f320db9edaa6279f80f96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e1d0e4583ecb8ca58ad3e575fc374d32f9f7a6ad8e857e0a3cec7b238b86d9004410519070a0448e1e0bcaafbcf89447559;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c80c0e3acf4608d56e212cebb2112be7321631b08eaa42e2c574975690a554389acbbf1aa9ce659fc112d1db3440db0ea2c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab165c368708a76b90d650a3dbc4d40e96d5a9fb2e31e8468c3f7ba0a843ec7af9b363725f572b79626fcec57bfb245e1c5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5caf2665caa1f370e08dc7bfb59390a9c59dbe18c7f7c7736a9ce3fc031640e77f6b647d04b7889c488355caecb09cd4c84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2f0d59adf8c5be23d3389fff2e9a4fb737353a1e17bd0bf20b8b06e8636644d428aa2536dc94d426891609c4e12197f96cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3876ba72ce51799a35deb936336044974c8918e98919a71dbba484745ba7950da4dee7ebcfbe6e4f0b739c69af9a1ac505a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31e6e0305b228838a05a2aa5e1df04946ef2bd6b3d64b0ea967cfddcee0b576551a8e9725e1b022d06b7d971fb033353a940;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he68d8d46f23ffb63d3aa8d18a42d61758baaa8d644025ab0e6e3f153f6e56f8b3a33c4e9ae585f4fb44127287ceb034c2291;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4465175d8c470cb89d5381a07461612df5f9bf07376dbcf4d58dc2d851b3769dd1c7c4fe5f76f66a41db436a40e56d5ff8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c0d84f79edceb0b9ec95eba939df2517f347755e28df34d68eb680fe2e80e1c234997c96452bddcfb63d65424c534cb80ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e7d459a6b89e3bc37b4115478dd7d390c24a74a74bd31816ac5627eadaeb584e70b972806a3ff8d391a89a92c1318a3940a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2750667c5299e4c9f650a246f4c728f215adc8bd5effc582fc45af63c59df14d4e6768acd73aa1ff0957730e3767e48c3f65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadaafc9b2e1be69ed0319537e7db0ab76f1b61552c03ad42f2cd4640736760d78e67356f37d2738ed4dc3f76bdd22792d323;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h322578abb33d5fc292dfef032ff86550891d649ebe8e93397f5c85f067cc88b245d3ea4619fc57ec99e1d6c5d1ef0a8f963b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaa33ce51fca511a279c9a98a56fd6c7e68ea21a4c467e134757e005fdbd1415c12c40faba4828d737304b404e4c9bc5fba7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd738a2ea5085657ba576697ac4e782c252edbca31593054b998673554b0f7d864cceb2ae858740c15767ee2924896b80517c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ff1179e2755e8be6c07a8ed2eede6610adad0496febe846bf4e78b3917c342e39671c5b0a601512f785b2b53d450ed8cd71;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74e34658d8014d210e8560dee0b6617630d769a4bb0827ea5b60e27145f6330bf84d3c18843c2f5c2cc99c8fe28b14e67d42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf7759b4a95ceb88ed76d574e8d4e436de0116db1c813ede2310c930fa666e1f67b0f3dedbab9548f6ad1ce1ef9d2c8abdb8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e43227dd3d1ba41274ead95a3819e390174a5ae8b1f341d1dfac2fb42468226742b2d9c9b2a8abe496fbe7ceb9c0b20e0f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47f9e1603a8f7b8dee610270bda760059c94815a74e1b5c9c146efcc87d97c71fd519be9b857f85e044227d651819d0e9640;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4565381a69c50888fae61972cf4268029ca85ec28a7aedda57e8385d0de9420cadce08a95e44704ad21f60569142adc7965f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24975c51c290ab3076edd2ff51691b32359d07c41e994c14ff7edc65579666f8b1fe5de36326e96ee2c7001287fd15eae4cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc36b2e40bf29a8318837475c0548f9822de4cdb37b7411796fdef9c3ef7c7b4713c79240d731886de048868ec9040f007c75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2f50bca692254ba50560ee46ed061273db75a661b46c3db41ad89ff9142dfca2b07724d81e9724851c9d49649affd6dd16c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54889afb264787da3fc688f6a7e00c436a711058c6f7f3f88fe45fc1bcf47686f765f35273d54bce69646d42196ec727af53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5fad247941f3fb079b2a237274b8fb2ab7f3d75e15e2d8dc38d84089e600835c740f107fe88ef59959a3bb9952ae8c8e7a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5e7b69e7e7deee6d7de9db8ff445d112cdc5fde243c2619d1ebbdb06227a29b0568b8544d4fbd5e60b6a87b363f430683da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22fe5ba00710fb0fda1a0cc891bc56314d75e84ceaa6b5ed06696d9e0e66cb9f8cdec0eb689c65049a1e05874484475e0366;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52cead43f534848e2f312be9e1dc0d38b688785498d1289f29b65929b00d7cfc02b5a9a34f189c997cc7f05fcf8ac34b967;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72dd445726bfa0cdf4bee7d6938747f0f9f86115523ddc7766ab09467945d94d80b611890ee6c036054769969f0130c87170;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6b3a4e597f84e4645b31d92e015055e5cd4e436a6af9a9fedbc154888cfc1be2fb540c29c60204ebf9ce6aeaf21521787f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf65080af899c8aaba8770ad7bc98e69c983aaafee699f025347e14c55cc4b112316226ee1127721fcf10794ba9da968fa231;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9caddbc315dd8b06b8dfe741580e2971ea4df58056552ad6af384666c598fedf0e562d50f72c5cbba7d7d2195739caee6e69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3d1cd48ee68e706d83451a07fe80ab96490d3ef91b1fbc5a623567e6f3e48026b3d9ec846d948e8fe0e6152234557e57712;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee94cbd78cf399219430ba1a96b6e0b9bb21f127ab9d893d6855b71b3a00d5daac94a407902e5adde1b4ffe7f8f12d77944;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ef8f6af3b5255365a8a98630dd348135a56505380c484afb1a4b240ea3990d7439d800acdd44f054e17ed74959f5ea593b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f0d23f6eba8873d24447cffe1d4647dbdf95e03599a58100ed8a30c4ebc05dfe893fcf678f0e823f720bee8f4f6405c01ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h915f2d5d42d5a32fc8a86faef441cd7f4a4eeaf897b03b27d60088f4bfa9e12359e4107c322a17f92a500f7b8836f2704c7f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5024d7847ce2cbcad4f4ce3441a47235469804e71fce189fc115f5ee681dcac9750b36272c22b062f938f296cd116266016f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3656fc37db7954e9573282455f6377ad61474d2c7487a0aa15bbd8b92458e746905b199a82a332932b62d74cb83d3aec5b39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4126995e6f3fa55ba39bfc7e881c1754f371fd561144f16f1665808b8e802569fbfe94358caa5caab2d2ab82f92b9590ea6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h298d11cf5e06e8e3787959b0a9f5b9ca5c470af2318600e308a086f6441c39badfea52538f14816fe11b6d1cacf257856a00;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3887b6c8e1ce088562b422f6dfdd31c517eddc1dea1c7d31010408e11f907815c8a8693e7842b49357aba81076e368e6a33a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83f197a7fe443d925aa7713e7fa464f22966581fb7ff512e49998957966a827ea31a2f52938bbc03a8e42fe6064b4805c410;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a488d2e77344213c7ab4d758f67571f6aa9b1345dc62c7eed737a5d01174f72a61c382ccbe6b300143df05265d1837f5fff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8967c858f420ef19d76e9d0386812cd9c8c55074717fa9f48fdcbadd73847a43c09240a716beff84cb7c9444bcbdbd17c96e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h521b68328be2263559f00a0e02990b8f585b5e7123bd6bed1e641c5daaf22d9ca16a16dbec39789e02652d6363ab7887c979;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf250fcd86fc53a45295b577fea6906124b25024b7028a31e8ecef4683e57867f27d1c34023800148e5b8e579d818f039005;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbba60e6684cea713523343fce7a865d2e7df507ce694b7d797416a33a835afc6d62cad80de5c8e7cc38b9dc0fa41614e1861;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h693c88e0ebe01009014cfe52c0fbbae9a1cc98293197a50193b8274aa61b18e6c31d37b5b14c84574e37935ed28ccca1b16e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h325d0ab71427687a3bb0d29d2ad890a2b232c1fa445ccf74fa33ed336f7a76a07a2bf3abe1634b5ae058700e727227fc87d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h581efbf39295aa10a195f0115d30b4f8186e53c3bfce5cbf9be12d53e49f87c0351541adc68c0889fa3202819a48ce5f4385;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h359ee1934e81e6065ba07d85cbb28ac58e614702a5cff52e154fa6c9aa68bf2371d64d1128366f288216f8b4d03b44edd585;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h920d72a758548e0feaef9831d1d77748a6eafefc626d9d1dcc80dba8fc6a535538eae4610b20e978803c9cb4ab055402c139;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb95a78eb5b8a3cce8dc5f8a13a5893894e5fe08421fb9f20e57daaeb35beef5f6aa41437e5ed762a0b39e031d17160d0b17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h311f7b1303309a34c1b4a1abb971c1a50a8b4d575b91ad21fe62bb00feac645334a304652fa7981de3ece7aefbc96e3f92d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61429b979cea19cd8edd8379b5e840732030231220cd7446f0c7b92fb02f5a0288dcf6e7accebc66ad0eac7ad72a0dea398f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15267d67ebf174921c5d7935d77f34136ed4380b50a14e863f29bbff7f3c6cb55750391c4befb64cb7ec55482cf0609b463c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda0b97fea0db9a49e903a5885fef784dd004f0431ab8fb75acd68de790cda2083f8cf0cab95f65d1baccbbe7bb7efa07faaa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc39725501dabe3854b2c7947c769f2d9a56d9b16c1778dd56f68964b5d2a99d01d5c6ffa37a05ffe470cb6d99e2305df1ded;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8869ee820ab49cf58f8fbd612f6d3c730ec534ced4beba0c8c96b0fee8374be7dd6b5f8353941f55a2413a1ac6d0ecea7a10;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha466ae0f8b4b429adba557d07e36769ce8596c16ed800f227995308a3f8c2c9b9014de6b7f99522846aa7c20277d01482ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46eccedb4f41d2702240fa78bbc6dfaac8701febda58f0484cffda8a3a2763fe5e5b590f963427640a14ace99241d1ec2944;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb89d8704d4a8fcc646055100743dbbf49c9956326bc927d216bc9b10122fca139a95ed435417b6ceca22a95cb0c34cae1460;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75215b17c49f205751ba6e4e45e1b7d1999f6871179d0b0464ef5993560db927ea7d52e9b4091634a79c2a6d011a45ef6eea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha80202c0fefebcae31570c79d5f200c23d6ac7a67b7a9484226acc8721c756413209398707895b1a6efa841a1c72efc77f4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha781d3bffb1d79eb1f4d7f40ad56a9c6e24c68a4d973bca9b3349f68edadd6a726a88ee3ff865431df4776a23bd6cf7cea0c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a8c4576f7de19986715c04b0789cef79937101c1ed5fb7917531c0c5e75bed100bab1f6a3ac5d1d04cc3180fc49b74408a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a036ce3edc5f438058ade792cdd46954693da845d4795ba8caf44df02a40af1f6217a106900a16907b1cbbee500e32d2022;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc33b20f2fd134a3e20641e12dd0cfa103d8230ce8602c4978b0876b3cd9d393da6d81da0dc9e560df1ff701cf305d4378a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h961f02d160ba572b97d803e38804bcbed17e5042d251bb4a49fcedc3a2fbe04d606e5617c7162edd1c5e0c15cfea79d1c8b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68366d8f3997ae15a065a6ff0fff18dde4998e59fdd8d87cc645835e214b7be26ade7f3112e27ed81a3726cd89402a94b3a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dd9f6de480e3e9a352667ad74fec83b8f13a5ffd19ba38bb5bf7ca912c2d4425c415cd78b6a90c74e8e19894ac8a380a195;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8b2e0956bda1c21c4b13c1d3b1711506e4b707486b301b4a3c45892f995938ec70518a3a9d3b910e9c50b879b6b3c50fd15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2978cf6134abf02e77cb55f12396c254c3db9421ddee0b47c0a42dd9fc60034cc52d4d70081351cc3ed12a2b718569b7721;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed626d69350b7e461f734b1951074a5e32a8e23f34717d53c8289053313e5c5f3382fc6d42187fccd029703aa4e1cce6144a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a4caf134059167df420bbd1320e9c9922350ad330633bca5e614268b38eecbc9cae02046c01b548a7aa5b64533f6ef2b884;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h301bc7906dad5083a3aa24ed36eccf3263759f577cfdd419072762476c3c6e9f44ca291fac57546c83b8d4d4b71e5facf4e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81011f4023f79e484692da389670d079196730d6e64005751bb5b19eaa631fc2375c4e787c8a44977f9f04a75dc46e01aaa7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h275c9eb4948f8071e785dcc25b1b830cf30f85503b7274ae5e9d08cc403d8ac795d06843da7fb92095d61377d4dd1a3ee129;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd36e371b47445005f2deb376528e8bab898793c7d446a34c1943b5c6c4b42349ee908fbb62e16ca1eca41e83910e0f1f0652;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha650ac4f8c60201a965125f32fdd77cde9620c7f2e3cc423ede0c13a5a0bbc7d7e55769e2e5651e8334049349a93185a21bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc018b23b7c91b4be1ad9093245772b8a17e42abd5946926eeba3d01d0c56932d8728c8120e6f0a9fa2f97c2cead1d8ab346b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a7694953828b95e1bfa587bf2584007739600b204faeab9ab0de646768cf1507bf5ec39701c709fd9ad54c8169c404babfb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7c5929183147916585e1ffa25ff48b130dc607b5a36df6e14afd2fdc6e88d2437177ba396ced13ad376ed509f4d82f0532c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd161f73b52d53a0c43d6885014661eabf718e2dceb5e977bc3aca77db854d85f7560e7f07cfcfb278a0522794422ab717774;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a74f9329edef3c7a807e52b6888ddb195bccf7b902325dbe63dd2ccd0deb47ec5cdfb869f74ee8b065d342318bf42c9d0c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ef559a0e6d4f26e6f580f56b64f27db1e221c53df2b7bffa331744219ea1457787cfc6133602915eb0335eb7ed06459dee6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa5812c1823f0639cea2cff9bce15d3f0d5b2da425b14bae2e3345303012671c6660b9c93508b36bfa9bc3e2282e40ea0241;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h694922c7a3319dc587b79ab49fcb493788214192b17c92c7abbaf5d47fc62bcde561f78a99656fa43e8f37dab7f9cb69cf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ba61951ce70adb37321deff1032611028941cdd3c57cd36bf97d4fb5882e52a6b6e6a23dc296795982c04e328a7d5ab76f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h895db5c09798b4699e2ff2d938ffa51208ab653c5a262a97eb5da61fd71af4205dabc001761dae59d8a159692e17b2266598;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae99ff60be952f99c1879a71916b3d2090d62cfd04e60d5e7b14fd96a5a88b8888c2add1945df18dae4ea50814002906b00c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f7129dcb69fcf3d576aab253c387f57f4b9057835b08bac329e5f54a60e4569fadce0662bff7144a6f0e7fca164d52b3c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77ab45d84c310677a478919381f1b8986d073838b528b5bccec093eb4c029421e4d94afbea3aa9564bc75fa3c168ea14037f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5fffc87878329d5506d3c88d5b57375d035c78cac382650b0dffb5ac270bbec554cf4a34ce113c88b2a6da60f53fe9e6cf5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5131db7f718ca633b0d11d3361f341bb9e3ce5817021c312baf0c573437c92641b6013858ba466dc2ffa029e2d36f1b79586;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ef8465e88ad0e5271b03531790030822a9dc045171ae3ea6faef552f9428b22d8118e0a4a22ce420a9c65d0101396bea8b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h255e26c058de1060b084df7677a1cd03fe1f6bec447c442a8e266e566c41a2eb3b6417c672363504f031de26faa0d5846629;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7be3ac022bd52b51610825d092dbba1491839613b2e979ffab192bf8e0ffcd06e3c74fab441e847f99ccbb0c2809649cadb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51c4f043180a6668516c902c21d32f03db075a9c5a0d9694564502a62c4f4aa985e5865bee49d712950ef4cae17a407b3fed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb9f5128b735364c74ba122d6129e1b8c9e487270fc148a52a37d06a7c8ee1c41bd6c9e70f711ee5264cfa502a537602d30;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb2e7d5090baa2b7a6ffbe13f9dde9bffed5e2089f545ff09da7b061686087c055739b4a4f43e5b9576edde790a8d8610488;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3816f61f03cff8311d75a0519f8590f68d37ab194fb961f3983f3272254495255209851fa75bda21f7516735585bab9e4251;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6440d65bc0ff91588c78ec3ecda8bfa405bcf58ca63a312220320f3c3163de9094bad999a69d02df650e85a2cc851c0b2e8f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee1ce6f8cd0cd58cb2085c30d904ef3512903132748f7349704b1d85e8f1cc17543a87351fee23045ce43e54836ee28dfae1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h380ee15fab89c18dd75dd6ef7b65c284d6c5f30193a61241204989bff22d57f983b27b03ba4c32801171f50ab194692c72d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1560a28e0fd8fe9cb45dacf94bd6c80d57e2af4f33c977ed16316d5122920d78a577665e398829c31071a9abc4120bcdfdd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h819d1329e6c0b9cc0e06fcfcd6a5632e581698d47346174c47f83fb6d1140d57f7f5194b5e3c9a8a6eaec29b9618fe868d08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30e1cfa0c6d6eee736e9fc326152e2a550aaf7fac24848155de56f15f0217d206f857e3fb9b907429598ea5150bbaa763aa6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa70948fe75bc89f3ba961c7023c678d407a05296b6c292f14b6b82634cb4cd0ea32ecbe0682bbad48620ca90bda092187eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f805b632c6c27f871778ec26ab0c349a6f2bf34078e2440c44190c3920790fb9fb462baa4ca3f8812181fb93712f27c61be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d81752dd0719542328cf0364550c380a5ae7417b34da810234e4a47b3f7de58df676cb74c74948938203822e153f7080724;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a5eeba5f20cb023ea26ae38d76881bfc081b188c0119bbfb4acb945f072277ebdfb5ac293df9b3918a37c1d265d6b93abc6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6eb63c923d2a934348869ade0e1c0caf809040846d27c0882374e6e9cb56449291a177905480ccc1f84f24512a22523c300;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c00ad07ea19e393586acca7ceeab33d9a10f1b220b92e724046c3fe056bb88de4e2c5dd1c7f9ab921ca3ca210f2b4996652;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h955c2b2ed19aa4a672c8fe638b455938875e55e8b8376817dba86ad1aff6957b1a4ee84eb15637bf71f2a0289bfe95de7dee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h119b280455b1e892184d82d2fc1fe8eb051655a8da17d59e2c3776ece9606d59ed1cfba8ebe0e7cae2d4313a975cad61372f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83d1510c40b2039045a958064b3768f2db17385528ced3f414190b4850875a3e44fc6d46e27e2e765ff643a74d83a91d5564;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf2b6af26c88d49a1cbe02cf81a6813a00b3be05af4ff9f54dfb038c407cd195c4d2591c5d7bafe3c187bd6141926fbd4c3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h481c94b6ba609945e6a1983634e1653e3f63cf3110d45a7f8a1961c43e440fd9b0e806edd45812bfc0f079111a6cb0ee5ab8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h676339f1911304082cf1df442254d9074527f05b061a0999ab81b6b89466d448e2bc9f5a356961f18bd95c0ffdf8addda594;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h407930c50f233657086f7112e634caebf8c10ca48dac2da2fc6e2b2ef5605841e1ade1d0ff90860b75c9388318ef1677bf4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3efb378e83527b15bfe9a3c8d0beade0058e2a4830b90a53bfe23e1470f52dbd75a43e1f76c890627af90722fa7cbd0aca4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf3ad569d84cd5798f7ccd5c6d3afa80b59d249ebb8d68c311220b613f0d5cf8b5ddaa593eb9645d30bca4df1371b4672ccd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a57c9a019680b178c76c9468283882b20fcc6c3f26d7d431c6a05d178f8f82d0b99501dbba8db092a8a795de1ce5f683f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b33586fd1cf36feb35990554b1dfdec159a98ba211b541525cf1020fee0b5b8db3036ca3772cc1db328dcdf2fad59d8c62d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h974ed75feee1b14be0c92d1505b9d79ced4cfa22523944335f07bc90668178a1ff9fd188664da83d4fc3ed1396ee4ec1134;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b6b8259e00ab3ffe61c47fd78df519c28a39d5788cec74add8b043c59f433b43c939371a8956823c6f60dada16a7b82e262;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66b3cce9c55316aa51857926d4e478f3f493a1b77a67a4e69a9f1944ccdd626f0eb950cfdd1449a5460453356964f188cfc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f3a6d80e3a0aa526e00d5c19cc494e07c5b574ef692477849fcb2c1aa27a1b5ce7c8cfb74baf61b6884e6730a526f3e6419;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf31870c5652635d53667b5300ef93acfc9d974f5529b20900feb2c936e48a02e12e6acacac2b1a2ced62c64c2a1ba0d343a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6511905e59f8ff017d9784adc05789c73da6ce1125d7c6cfadeb255bed12b397755cdd274ea6804464969da8eceed3c72f93;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd276645c880cf271ecd34e566b382da2d0c93c186eb1841e90d490e94f3d7d75ec1b15e571f2893c8cb4161607803bf0a05;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34f927166535fd1102db6a506e2badadd9ebfe9563bc4aab4222731d26592b94f2b7d607b04be1bace5e8e9f792992c88a01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb9766e072e09f78dd24734d44c55d4d0183cdc3c024de95a53cab058c30e006ea0545765de51165560eda1bac347e80ad5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he48361516ee8e002f324a4f1340f068f331bbdf4128fedeab12646aa9c3fa0e9b1e4e830159984f11153862ed86b2bd876b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ce4052e579b1c3c3beeba8ef9f1d8d124ca1affcaa5f8df1e2ab049b9d19da0e493156c4934cb5bf9a69b408f0410c43154;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha877d5b7872c0a53528c5c76e1f4053b16d7235bff5317474cfdbb69088b659e3a1c3bbc885a9fe95a02c9951ade737e2442;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6f4302a25e2c52ad4fc5860f894f5e1f596b682bed5624d25b46ae2180e0aa4fa09e6f98eda996740e8b90b6d7beb868dd6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h414f8789fa1f2bb8ff782c945dfa91e97096bbf5ef10ded47fe8295e5c2f6629fd2020168c21701e75ad4f1b585071d0dc49;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3aed80349b31edf89411fcb160ab353527acdf73b5ef96fd80ff70535b5f513a891cada674f5a7079ed8e22a61c451193be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77a007e4aae1b588b60ed9f22cc697a64d1293cd9e4eb26e1e2e2983c8eb8d03deb592420bc34432ab50ecbc634e8087bece;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf3ff5bf32398c18c2d8479e952ef9aadf424992abc672b28babf25cd0ab23cc865f54b34b6420b166618df79e513935c8f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e089d69da9037e59968f58f4ab7de0b194e5e5d8bced93622f97baba037b1240effc57b422fc0ac57a7fc532a8072546198;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54b14a6b76a0933f2340fb9388e7912679002f3e0d9d1e319b506f0d1156f163e1f1f64bbd84dd89a2134cc632d161ddfbf9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7776166ee127a096698e164e760608fa73014e6073058841ea1af50ea99b48ad3222ca402e1ce09ccee78f8b20c0cf315d22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bbc6efb1a86e64f20b6ff91c09513f4aee51b19f417166844dced3cfcee85b306e8082f7b1f035401b705df95eaa16911d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5881efbe656c82e2a82c1e946073c4d2d5ea06ffc604af08f349194f2994731e43b5de094ca1392395c22344b5e2e667fc6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ec94b91d508cf81eef334f50807ce0a5d4fef917d2fdbf36c8bdc05584a7b2c674891491622506d0489d5ce9eefd97bfadb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36eb75475bd34986560a3cd6e71f22b8e301057ed534114d293a991516d97970899d5abc2a7de3aa46dac87080d4cc8f8329;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc82e91a2e5f9970acdcbac474538528c9dfbfa171abf65e7418759bb6b449611ccf2182051cf786fb28d26a6cd47ccad4c36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47b6d7d89253acb242176d74c6f71f91dcb2600e0406d33fd1264f32eaf7271bdfa1c5b1784cf6cd683b9150548ceecd6ead;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac6f16aa0160d45fdab1c735f328c3ff86d004c33bb219b69df370196ac7ec07b3eb40500aeab177e701785b014c70bf07f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5982eb1c95770a6b2639a784ff8bfdc7389c34a8a2ec5d1bea03186d76d3c7dc30a3951ee95dc85e6e8a56011fc08ca90a38;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86af9eab347bf14c1969520167be3e011546825729a4608bb78b3bc3fe6493c1ec0e47b15167725a71c3240cb5968c26322e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h409e6b930ba1026e07e80bd20b89cf5b17671c8b6c4e27dac99411cdfb61a3ba7bf20f7c950593d86eba0d0aa7a12ac2806e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75a41271d988d9205ad9595a5804c267add1a1e23d39dc82210dff9417cbe86c8c63aa86f6e6de0e000abefb87d5b86ea1f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42b818cf9610d014cb8aa198a5924358cfb8837d6f05402aee19487bf18e1994ec46d909f364caa7518bd86c64568cb7be67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71e28fec686a5ebed1d843f774a1ab2a3dc538fa2de7c9fcde0f69f2191734dd49bc0a6325f0d0c28c9c877342bf14778864;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36669bc52eda81edc6a7fd9b790d85be1ad29ea07da304cc5fa18db3525a09184418a32cc75b1b005d9480ff47c26c4da7b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7bbcfae82a244b57be9c14cd315c745068a4b08e62f26fe935aa312faaccdd0aa7030d322b018d764cb4f191763c64ebc9a1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3138194729a244254a66c6bbb8cc979093c8f1679ab478ba3d2f626bd1ae85e2e6df7625525f6bbe72b95397a0d87569043d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8586b3f1abc6d4b7296be71aa39f54767fbc724dd8b42244bf0200e5dd9ddb59b82fb086f915112da0dc589726c56a3fca16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a4a470d2971b8cef80d095613d0597a51fc9a6a377aa9422247dda55ba43807ffa5758f37c581a31844ebe47c6a4035d977;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92110e73442e19a43a7b808196220b1e1472a7a80c01c0f30e52d9291defb9b05ac5c462f877583f6d779397fe466303983;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20c53ab150ae8916094e9dd7320619d540da74cdadb5e087f5daf82f094ab43c154327c989f9a54386ca2640d6dab1929e94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5d041b17bc9058bcef849606e621bbc9fb3e2feee9b3fbd5de3d84a9e1646ca6a0df86fea54d49dd327f89f47b938ba322;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7966da5f2b3b1e12cca7cf1762891da79281146f55550fc8536e1d61fda1d45f1db025946d4648efb780e68bc45657b44f00;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e9f7e8f376c09247ab4db0a12dc4d6346b1277c968da5f1067d28accb3647ab14b55435a8eccdbb0b523d7c16f523879bea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1966c0bb46bd1a69d4a4a8b0b05c949ae5b0cbf519b872480caedfd67f33d267abcaf2d13c6f1c423f4e47158b5f60aa649;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d417dd03310f171f670b2e53072d4ed5c3305729e8710c7e917e76d8b024bb1c161b07ea2e7654ba08527f9d8cc24b0d687;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17e220069dfcfe0494bdacb81e5ba9209731bcb17c25b690c42d9dd29b2378bd3cc7632774c286e9ead2415208bc802b0c42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c50528ef92d4a293b61aa45f527694133d3030c128a6bd6c0857809a0e948f8cd8b23163147b5a43e317f0605d7a7da60eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60a269ff5bdca3c3a0e8f97b01b02d5149045d3f2c656125cd71349a75c10913221e139ddaca2f717274b09b23c17e5dc1b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48d4d1f36259e8b249e1c768b2c32602d7a9305d7bccdc287c4411e27d9ba1cf9717c34728cc015705a5f87157d7e741f0b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h700e3fa09242deb8cdc38c4e38f0460551179f3261119f3d2a17c7e74018af3e493e7c00c3253e3b9b6bdb8244d7ebda4e68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccfd3f2b79eb3c12ad02c974c330c2e610b903044aa169dff5d6497fcf44255dd9e3f70f6c8d7655a3f9e9f6d37eeb3d6a4e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b29b4552191dbc7258e56d63e4e4355c6dbc85ec01c7ebb63209e004ca7180598df3424151321789859922bce1122baa9a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27e7dca2967d04bfb3a56ecadc56fa3a421a081ce33ac202202ce2b047370e10dbb1db0a9f0a8f88ff2817949a769d5f3b91;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19d976a8f6873df27fc884af9d532ce83a665663eb5f3bf058f8e2b3da1ecab5b632e75bbcc473ebf07067a51d73666867e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5b1e3c67ee61ce95e6455c65205b2259fbbf3e716017243bea48acd6464dc17a4c3af643faad6e06e4b4e9c72687139c9ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h867379c8aa76a3be50e8ad4f42ea00308a72bd6860cc0ad9a7fd4184eff3a6154e32cb23099e052b470e1ee6c034bda74461;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h436df61d9c13743d1bc56c57bb4f8b75a2fd553cd3eb665cc7b4441932b793982a2812f78c5131ecab59f312db3a71e8fe3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h486464dc0855332965454c0b39da188c0108876e885fd5b6786051a665e724fc315fe74a9c113437d4eb3928b9922cfec301;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9248409f970422253a4dd900449dcc78c137ec67e9b3d83554762f14220fe43f29c85d5ad1cf955544963629a8da4b791b21;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4317959a0cc35e038871ae723b9702265b5dde37f46b16996a925ffd3b3a5c107e9d29e910f8d9d95ff33d47764d99ab1b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02217d8da48c0a782f55652745d5ab7a55fada43eb7cf9a335b8fd9a2902ff65280a7cb73566461dd0f30546e85d98d6275;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6d2463984d933c4e9c1dd4865a5386c72874cf047e75f0e157977ad4fb19441736171b9d58259db7020ae503fa9a99cc936;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c8dc43da5d7cf6470488ae662e0f6868d64a41749e34c0a6a93e83203c046c32b8da160d71b11b38b2e74691ad50049fc8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had08f2d161785d60b6bd268676bf9c253685438a66d5672e4b5fe40e317b4f986e6a7e43736f6729b9bd77e5d610d43f5d04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf436705f66e26102298de18943208feec1056b6041af23309e37ebd5c33ab5fc45cb00656f15fd752005fbfdf88916b07254;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bdbe139bd45205487a20653c36e0a42df9317f23286056b51a9ed0aea0dab2fd7bcde20a4e2489fd995a46264292639a615;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb999020fe9aeb27335e045abf406485f56ac9a69f167514ac9d2985e869f4c93750d557b8b54330e3d3f6a16d983f391a8a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c6b1a153f517cb7ea0b1182669186e88c1086f6e1e11a3441229d05981cb56169b3eeb7de1bd77b3b4c096f5df7aac10eb4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafc94ed7f1f1c6981a4fe3e1326053ca93c4401cd71db362d0ff2c5f7ea5441c0994ae900d463708c829dbb4b060b4ae01d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb63823c820ca6e5efd7dde27889115b29c099cdb1d12647b87e7439ab041cb41bf3ed98f03315920c9df01abdedb9ca15fe3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf67cec8becc5d27c531b86a7eb40b18b2eb79ecee9f6952234c7a3b3880197fc888724238bbd46bc805ec47c556538859d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd1120bfb189aa2cc1bcbc6fda65f86843ee8b7c56d87b3a0a405f38a7e02bd77a233f7c057e71ddee9e25312fbff3d994b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd9a795cb18dbfd550ae953d160e132f36dbefe5852853856b27371ebf61b86673de3b9a87d2a877baca40e00afa9fbf0004;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5e0c930ae59332fc6934e33c847d901a7bada9431c01d1fc03868de9d3482110b98f1b940a064689e6070d6854bb7eb29e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he07815ce82935919d0ffbd5fa24741f33b228ecc3b4bfa0c20e3a20b63126212b74df764de8e3e5f858f6c6edfdae4efa9d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbad4d96edc91e28f32fa422d4530be79129d950e1ad3635b38c4c95651ab2c9209f289cd2397aa13b0b87745f45cf653217;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ea09dd234f63f9e516df870487db393e8f91dd844b2d5a9f1e8f0d65fff43f9cca5ac7dbdf38965465cfbc42bfa1932e425;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a4dbaaa84adebf87677315dd7672fcaec9eb7dfea9f53a1db09605266113e9cb1b097c5f4f70622d6d4d307da34bb48cd0c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26a3b65ae428593a0c843748cf203caa0e323ace4506819d478942f56e8125b381f3e4d5eff5406bf4a6e7c0266f29223bfb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb27dc3e9e5eb5207348fa7dcc0ef3613aee7466782daae1885c53e6aa974e4c219989d490637a7f1c5a40c1299ed47e25858;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he908ba701a082f51c3c89661f89ce9826c8c5a397dd0d55a0458ea41823eca6521a9ffb53814d4bc08e2a1fdc18bd4c87427;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45d22148928927a6c20bd6b5210d22a9211dbfa73ab89bd1b6911daf05c6464487a6a35004b7c6ab7c66931c26c8f899390d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf29ff1b9271bf53afb35f94d10843357bd306d35cbe1fc7c0ef2323ec3f2808278c2706e3afa2b12c5b715a25fd9d20a1274;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d74872851e5a9cba64645dd7758fbb7ef9750fd27a420c716b40a3edace0ac669109d6cc206449bd61fb07f18e5f786f927;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58286ebe9974fc9c675967777ffb3c5081ab2bdd24fc79a37f2b4d311142c892b4d5b3a228a16c73104df164d75fa02a96d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a70378215088ad9625555a489b055127221539045dc074ffc8c91f83ffd354000c201cf41ccf8c3938e6d539bd595c5b29a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8ee438fe31311e4c192392506cf3611666e91e82ebce17c4353dd1485b068b23b94b70b70e2daec7086cfaed1f31ea12793;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d220c99c8a95b5f25ddd9ec8a5b1fbd535cb6d6859078a33a89ca9a1a31a10d2af2b719d304a772babff819621fe89d8607;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd86cd06392fa1c678529d6f33f87d4607ee2e17c1b4feabdc88eef3f6f3b782ec87adcd94f5ce5e11954739cba8f6fdb5b0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f73efabf7a81e32cf6b379daa1d2da5e8736d4750d0638f2cb4a7215cd7eea7e2b2c7cd59ac0507272a29e93c65c68b1a4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a69cd66e7c96edc2dbaa4704cd93daa7ace42265e7918f184257a5850feb8c9b7811517014afb4015526a3697cd16254525;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd372c057e4b40412bab6fab5a3cf63c4345fdc0fb1df01b0b7c3dbeb5aa72e9903684ccd94c7758b41f60eefb3b29ebd5843;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd142766ab50c23b51440ed09d4045a760c59a82bc5f8f5246bfb5d91c5b54442c64b904a61123f35302ff5d605c9a4156638;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he31fdb4305b97257ce6adc6e98d12842acd1867ba23daddae28617ed6f87b8a9d372fd8adf27ea3c2ee233a53d6f22d0aae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81a90d67d7fef1af53703000bb5aa00e0e6a60dd182dd37b2a6a57833a564ca4d94f7cfe0fa247cb3ae92411ad9f68d86ba4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb010c09d20114c4515f476cf4b64f543c13abc4fabba7e54b327afd7b6343af95e9a90ff32bd869157637ee01b0e2848368f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ec1fdbda74cb810650c93972cd261b251ee861459a715b58cbbcbc04d8cbc53155cbe2c2d56a243610598d504d5f2204596;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habb8df565204c0c7e5afe92aa95286c52ecb652b3af953167eb1865c00d25602c7814958c52f82a547db054be261afb55797;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a4ae9a43d76dbae597c95243f626e510cbf282d1a4361d993f28c104edcd1625d80f8f289f8776866f3cac4d949f8d29d1d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc83f6e28571c3216c4c152a6182fd42fa4ef61bae71d5ea6a6b5a7659ae568636d98515030c621981284e8a0547054f91c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf7937fd6bfa93b67ca8be968f3c9aab45d04ac65e4f497392909a5cad96f4dd623e84899023d95092b998a10ac781b3b996;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d6839b321c4e75341a0b025c6c057e04ce1613d4faa1d19dcec174793bdff22462bb2ac3ef5492226d0ed6838c872a2506d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc747d9319fa5a2dfe14d566b7388dff9655ce7909b2cee1aa2688d81b284f0382cab52e80f23151bd0a33364f1901788232;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6056c74fe3bb72be21ae896da16171e3a076302979a3aec8c11dfe6f8371e79bfed40da22e567c8b0ff7e4927947e411ef3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9681aa894452a6e867b0de5c534613072b311734eab0e6d2cf5a102e467887769cb11609fd3c0f8ee2b112aa04bb3cf829fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb400a9d4d330becd3aa3cd0e7e8ef08a564434f66c2e078dc0a6c3149658c6e30809bf1687cb87b1b51a6dbb4e813de08a36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h984576d0dd08e78d72b728ce5c6878f76d2997594f7a30bb48e80782c53274e03a446909d197ca68819447d5d1636afd1ad9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd14d0aa9f24016bd63da91cfc1ca5c78de747080c7081c6b07ccb4758aef78cd6525fd25a477f270a390d7ee9241ae70ab4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha28d1a7e87aadb463c759d0f72b45faddcdcc6c657c17190e71250c7c37d55332d02bbec2d473bfc8d1aca72d32322daaf42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf610513566abf8517383d12f4bed0069bbe7cbf7aed4e8761244856bb3ae5e633c9cd0ffdb7a3613954bf08a314e4670482b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1d91140b44373c382bfe0045cbf39f86d2ae16f1a4ef647c768ff9f2b8a801c62a329574b5f83ee91432284b3d5b51a6266;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2b9f68ffafe6e827bcd108632c6ee15d47ac0448ada60fddabbe148206893d2ce42b6659b83fb6ad6734611f8c935f30926;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85a56fa8262e880cbc7a1d587fc3aeccd593476555577d8b2180c35bb4d8c00649157b3da13fae73ed819aeb402ce98648e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9194b389542a3e77df3525905951572227017c752fe6900006d2fa11ba3d320635f3cab01deb27bab687e2baba23a3435bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb556603b3f428e1916daaecd998036cad64ecf65d5d5863d7091359b2683101b2f8b66146c756a6e80dda398adf2c45a690;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h437a0ffc95a11ea0a02ffa0daf50080dc206e9284acc9b4bca53b8ebf4e3015f807a21c741659c4850e23ec3af9a4726af2c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf4350a3d729ce96ae96c578cb0f7cd9f8aa30acb0ef0a330cbb9ce21976639f755a8c041e974694fba1958c27cb883571d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf856988c53e5aa49b142c426662a8131805ebe2c968490f31933e8da66232e5250d4a84952bef0f36decb59d7b54274a0967;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24d6ee1a64609cc7c375c7fc6f96fc1efc75a7305509b9a57c2226031e17d2bc9a8026c5564f1b9cd7f782c239ce4ecdc5da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f11882543463cce01a7baf5fe4cc290bc6c607a079cb86fd82bbe33996e589f1c96500bdb8d5382291ebddcc219bdcc22d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1c7161d24ba82e5e2285f298dcb0ada39415b41d48b739b2763eab193c0e67d4a3e476fb754d3c66d069d73c098168ee322;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb7c6e73f1132517ce7abacb20c31debdd2018d75bf4152255353b91517e1979df8f6b1c19551ada2b026e37af8d5976b390;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a03599f6918d88aa0d2dd7d18d00e3c5422830a9f60287127c0be50844e9a56641df8c11b89ab21bcc773973dc2c338ae4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbce0663b4596ad47187a9a78c8c8978077c538b34d531f38210f14ca8e5d8225c81148611ce8340cd4c268453733c6058b54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf49eaf73c5b7c51feceebc1b543eae9f83c704425f3273f25e83c1936fbf62a73460ae28385f5fa88f1c926bdceeb68d150f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dc15421e7c37935246cbd53a623da894aef5479f35ba5531dbec9788af6a74585a89e380031aa422b074ff96f8a3eb79be0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a4bde0b45796b80b954164226800603f9ba5ca2aa6f64479eb4983ce5c6d4181405caf3fde6ddef26eaa3007d3ab0ceee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ebf02caf1bee976666f1ab60b59d527ebb327b026dc435dc970ea809920cb89d07758e915f171df0e5372af197b39bb79ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd96ff3756874d30ecb799efe43bfe31d5219c48f1ab6a61924f47b5a2d00258a65588dfe03a7b8621d1007e60cfdad072a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf20b2bbfaef684cb0d3f8f0f56f5332247f8bc1006b257b421a753c46a332c052780155f7eb010378772b7e53ba7d933f128;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd686485795e5e3287caf3329564e6ca3deae6f73f920684fe820c74bf5b64b52c165cf297a2167403018b7ddb896e9d57856;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4aa98f21316ec489ed4f92f15582aafcc87873c252e2f15f80ff7998389017ac73817ba476d5b796b0f1d230ea06db66db9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34d3d0b328a98c771812d12fc200e17ae31fb82974fcfbc48ba98ee423832440b2d65e0c9c75d46e7fb8659e9dd76e560b9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f47ba6beed8ee5aaa52213dc70f501724a81b588af12cbae1bed97c2f26f152a48921da230b6b1f69983c0eb9e5c554543f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h535c9f19fecbe46332b852c2beb8a6a8f3a8bf51a4d2de36ead94fda01f34aa1475cc0aebec2e8e27ad3b968f87902e0c52e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29f9a05619f942472d6efeb6ae0fdd30b1066b8df28d495aaa5e573930d724af730b37e8841eed2e490120b979b4f9095c4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h318d31d2c5b7c3c9f945c92e10ced9295f4f0edba19f7fb3625dda50526add2033aec4d5a0c51c057f3b8dd177a228fd0e92;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ca6b82154c996ca7cfe571f3be5f23dd74653dfc9965bdb5d65f3ff0edce066e8d065dfab76d397663f95dfc99171646407;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1d9077a1f73c1b3957e4e3beec56f7162e1d96857c0d7a4b3a0ba503112bf1ed4e6086dd90aabbd06cad455dfb13c925afa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdeca2ac8195c1e5b6b0f2baca39aca1adf1ba7caaed461e64ef6152fd41578f8d5e9ccb922fb2dce439c7037056e568379f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf038465528ccb504e07e2566331ca9312e143ff75eeff694aab09f93aef766324c2219e16b7bb1133fc7772d5c3332afc66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2700d26397e3a3e13c78538bc7532202cc8ed99d9822a186eb27bdaf116573d5dc435dff04720b695a123c3a5302a00dcefb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea46d720e73a203d2bef2defc6f190a920c6cfb8f649e439f9ff6aa916fb896d66c7f3b4ea2ede40170737e083bf465db02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha08b1ebfa02ef99a9e2bcc74cd56184ff234259e040c9479f37914e4d26b959214204734aa362cfea7769ce4bbbe05d37a78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18c7f7b5d1a9b6480fe27aae2aa57530eb5b687cc3cc9d050a1dc78795f0a693fa2aaa28cb3415167d3022a2736f9374f78d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5d0f17730847aa9634f53f6b111567564fe3070c9940d477cb1f2781186dd6783ca09fbcd3499d6de7c22d371ae4b55b5ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf4d80b8037c09185d6a8341b0d255f01ba41acb428359ceb33f7cfa6ab6ac0446add1af489721b2ed77630b4b69fc228302;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9443f5df924cb26c66460dea36ffaa43a5fd2e487a799982020a4373037c1a1643e7d52cc333238bb37dcd07aab1c53e4b20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h229f7d2ebc327acf6fabac4b2b5f6f15bf797a4cd0638975eefabf3c14aae91e7f64f0a0299d2daa67b329e5f6abf78574e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c923f77624af1c2541788d186d53727e64582f385bcb4336bb3ed1d7c92450e0387c830cb95b20b8bb5625b7c7fd89b461f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4dec7d3f48e48d34980f1c78cd2740c6cabf0c43d67db0d6d2968ef0736e6491226421830c543f5e697147e1f1b5d9e2f15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10c6f614af448dbddf2cd31fc401553c5f6787c04b561ee732898058373c46a23f616c8a9cbe97f77da1259a898347c70186;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5b215cc46b98043c6dd39a550ddaf3f46a327d60ce0a47794322ac82354ec65f49ed2bc8dd88a82064bc77bcca655d3cac8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7334b13917c9c2da9b7103e71cf30412c1bf4e3f7b5a7e79e8b3592f30a01ef91dede25cedd17dabda6c68d1861007ccf08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59e85d49ab5bd1b45801b78310d3eda75be4ec44f897d398c6ed2cd09e357785e3b4b9c68df147ab08741c8039fedf509ddf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdcb1adc41b7d1e256a923cef840dff863efdc1d9dcc92700bd22e2d9f45a163fa79717b7601367d7c8a9c45d83dd4551549e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c91b45c1228fdb83d5b5ff300266d883f32fc8b5e2be0d0b037ba14d13bea200f93907775b7dbc00d87e749fd6a7f75657a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18484ee7c09e85a7ff0d233e6d2576eff95b6dce871f0b832b63f6d09aa4745d69128600aa8c22ca844548706959bde00817;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6c4c024f7c2ede499e8a97cf37f4899c26dfe9265889a2ba89251df19a547bf5af15a1d39e98ecaa7ab2f4ebdaded950951;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16bac217d504e799230e7e31310bacc1636eb60d78a45d12fe67acf4bc982327b16c097d1d3f6ed04a359d723e29ed23d1f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b6135fe4e08c496cffa2b4d0294c0408ed9d10609ae934b8d8e444c3f29776796311520c6e7aac55773a2ce84e05ae67d34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h226428330d2057dc13f4d495b1cb9e33d11cbee53679d6945dcd4cb5928b6ecb24ac68756a43bfa3e73114178f3779f12d0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35f039644fe9a1db24ce82827fa0162d8be557f7078aed7fccd374012456b54dbbacb4b3c7b291a01d386815ae606eeba758;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2a8314862ad13a78f322361478f1cc847f59b12e025cd22a04ac59c41318ddc07a40ff143bfadeb550f24af76ea20da418d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40c579e2630d29712e35cedced02650263c3af3247b8e6d48d81372ff13d9df4286d117fbab0595fe794e897edfc89aa960;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h780af13f04fa04002c45f2f1115425421166540c8c8dd45a92f6822c0b343113eaceb540fe366720297e10bf1e112cece468;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74374020e63407662b2763a9cae8ef50f62f1583be0b5729551e73b6a8ef30ce03add11b39a96250e975ddbb11ae152db441;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h730acfb6f29c7bbd139a1bcaaeddce35e0d3cc7d32af779916beb6aa8cd7671e79b1ce819071ab8beab39c4498a2dd3bb3cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e26cbf20000f682c60fb5e2f8cd5916df5aae5114eb204ab9543092d877186c8b46cae2e183ca9043c85cafa1027df9710f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda1f90024ef021fbbb53e97589bcaf1aa5662b39a4165fd542a595c172e6bcf169d08040a2620d5951e3c5c1ebcd23b5825c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d1fc911858f89547b4deced4eedf277772b903b1965f1e560f7f114c364f9a6a8941e942b2431131174b02986b658c40e4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8698a475ac5b33c78258596ffc532690a8687b8b39037f95a6df0f0040e4713c1f0c0f5e9d8e0ac4f0690883d1406c8cc17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4b71559bba39b11c8d16fcd8d3938752ab4a67c27bb981e26616921ab684b60983a57768084c716931be9c9a5ef03bf4636;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h264ade628e3d44404febfa3c040f7cad6c9001281c75315bda96695a07fe3bbf8e6042619bdeffd03367b7eb3f79d7070ef3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4c496ecca5be98d3d9bd95f343104df302b7fe723b27ba15ec5a5471efd72942964d951b1387c04fab0ee10d730299a716f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdb947abf6d554920c34cda8db1b742ffc3d8b4814fffb0a73a602097d8fa0fda113c86d5748febf573dd57f981da301d9c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb402faff4379610866ef0b6af5664e85d233dd87f9fa4439f08073bea2fe6beef14a9050e30baeb1b2431f173dd4964a0ecd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf02e6946ede48a30a3f091286dff32dda50f08c429f8cd518f97e836d72a25396138c9d01f00819f18f2aa2d4ed916f2aeed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ad7653de05157366c4ab6c24bfc5f2e2cbafd80183a094f1d2fae9a70aeaae73e02f957373021e852bab39986ade0bc4959;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4808752f33f8e8da900f0146c3a65c9c3dc58878912190e776d429b5daf7fb199d8ec497a0d5652ae6765e4dfedde025073;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98cbbefca48235bb50f36d3137d15c681ab9202ce2c7dbe298b65e14a310105635d2d1795027c881e0b897433f3953b3c3d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h812668ac2cb5244838f958cac3a0b316ce9846e1bd2c239e15116888ef8d724aa30d8b5649781a4d8b45f27d2fb3395be31a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55e0c128eec5f207b714f3942f0c626e5b93b8f6507624407a2a52c4a64cb39326f98a7ad6cf575451fa91852289bf2f8d98;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4403abf9776e872a980d9017311db192aa2a6e7a89af56f2a23a2b18fc1074c94246dfa35644b74ce80da4b8497e3e6d0e13;
        #1
        $finish();
    end
endmodule
