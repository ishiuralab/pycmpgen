module testbench();
    reg [19:0] src0;
    reg [19:0] src1;
    reg [19:0] src2;
    reg [19:0] src3;
    reg [19:0] src4;
    reg [19:0] src5;
    reg [19:0] src6;
    reg [19:0] src7;
    reg [19:0] src8;
    reg [19:0] src9;
    reg [19:0] src10;
    reg [19:0] src11;
    reg [19:0] src12;
    reg [19:0] src13;
    reg [19:0] src14;
    reg [19:0] src15;
    reg [19:0] src16;
    reg [19:0] src17;
    reg [19:0] src18;
    reg [19:0] src19;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11cef45626b89ca53e35094bc995e84b861a71399cc8a5b96a7379e95750b740cb9a6663d6fc7d1b422c5cf26f39a8378e24;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd8172bf71be1b9f54ea39f7b21b8f12008ea8aad0d82066adec738b0944422557330c31de0fdd8250e159f9cd6f741d4668;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ec52e5eedf92b4467b5328fdc22b01fd673a10943be9afb77b4d334930229d71fc83cd8f35d7062b29b5debfdb2a6caf5b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90297dcb90887215411046f715ed9b96a7935f64f1368e193afede2e696b970fbbfb75bc2d22d9a5d2eecc31f796efe376bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b4c3f9b93c5a695c957a082986c5fc814c8453ecc0a65f16d964c497602a6f875ae1de2d862fdf8813f9b179f17660e2146;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h347577416639907a9e464b83c2e0e7e4166941e3b620793fe7bff79a616806a46aa02e51761307187e59187b8caa26d0ed91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26b351945f00c97575c28526afd94f09ef480a7a0cc3c3d0faa47938c47ead24039e922e541f572955e1887efff2c7e1071c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17d197beabda792c53eea8a5359ffcc5d69a2a34c6ff03bf900957522b4085c04c55401715b3fddc705d31c03e9ac7512e64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71cb2232977c13675e4b25275b927bf1308f4ff1cef85ab3b0df25a0f1a009eb72ccf935c685892e6ad7b87b5f35910f1d02;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h596b2946c41d921281782911a84313af95ed8c6a1c7323aef7fae711521d12a65fd9cd6b0f7d6ea1e38c63d1f703e47127c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc69ee652053a9f92c0146b3843643ad2da01677bc160152f30d8c7493eafb8a6d8691f090a058282fd28c688fe4538f9ea5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8bf85612368d96f26f703c9e824ec44fcc5a52dd6ad5fc3e4b782298c13010a8912e8639330a7b739c41177008648187608;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bd1fdaac2802ce9ae02d4671fb7f7ba5507bcac8eb822b3b17afc7fece1364642d6706882d90d27bacf2c41875ecd746f48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76b71f2a4cfcfe412819f3506eaaf7f2073bacb66817211455cee6c86014af48cf6a64ae8728d803d155408a8f354de9df2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1029e5a87eef9ba029af4ebc0d9db5f7c05dd4002f9386ba76f08230c95d16e061f71e480cab0a79aa770d765fb2963eab3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85c85f3de10e9f9991660ddbbe960ec7f09278733a8f1ca3e9d790c3402b280b4eef0c54748ef814436ab5bb1e551a089146;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b593c66896368537143fa8718950deee12597969a2fe868b4938b3f1e2eea8df1546a0c73c4dec8e712859f706d4e3f6e70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d36730585e88407da65520c4a5a7fbb8c47f86121f4f701b38073df0de0ea5ec89afa170f638ae55f901fa8660a2ede517d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9fdf813f74903b48824b6a1c4449ef0f141940c5251c9bec0141aaa32f626b5c8e3aa2dcd7f8e1e1bdfc05169af6e903905;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d237d03598eb40931c473948716c306618abb816c622da14086548fa8f920582cc42ca18dd57f238abb735ef6f0ce507c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e6b19c350df59a84f6b97a5561b18fa9d73a88dc48a08d305aeff3cfeaaea21a78b8a94e8473b695df5d820b0c7becf0ec5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54729329a6bf4e8100ae31591224f5dd53abc5d8c32f266bd146075611b7c3dc7a57abeb0a508ea35140e0a5337145ace399;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe18e7af8efcfb81ddd6cede551068453f427e22ab142b33c8fbaa6200cc0531a43ff5c69e9b6ab544df2ab93142fb85c2cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90a9a90922e60c278536e2772461d927a5808f74d6ff6e493a25b124661e23089231c7480f49c2c178e69e23770787e044f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1b7e8db27786f873b24ddc65b9842f5aa277de13fbdbb4d35e0eb19cdab1b3f55861fae2bef1bf761fb66a406b267c8b818;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaa7af132f57c02019a25e480e068e00e5bee6a04ab78356a3a929db13e8fab1a63388ca5ec8289e18858b853b9540fc7102;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5508d212b2319ad2a5ef7ae7b8f83762bc77c3a6f0e6d52df3c3d6b88eb19a6d854370a935ef2f1297ffb7b1ba0cbcf5625;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1a7c08b6706676b52c3d8dd5d4b85ef425e8629e276fd086e73b1ea5bf67eb3d760f0571c3c42c27bfcd3f03bff6ee80920;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e5ee568c7dbd279a442cf74a2a3e421a030bab15cbbcbc6310dd8bd62669c2be38b4608c5c1646b30e365712a1690589e51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc855c8a9c755c33745629797810e475aa97db2b7708799ced3e7f452a5af86078e3e8a52f0cb25e38c734c245dea04ca1416;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h211d661756659d8e298e3f2eedcc821b7c67bc792ddd94c1a6121c918d3ee0573ec1dad0561e4b6f68fee13df38bb8eafa2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6106edba5f520c51cc3d13f41dcc0890be0d6b819d190c7e50c3fad53070b2c7e68d4c4e9a63cad3086d10f58fa1bba49ffa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc207532dfbb8e477a062fd68ace7c623a33611fa7d58c30fb4f1f669cfdbddb6bb6103717e999eff6e3981fb48078893b55;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfe239b0acbe82bc76d66e47cb4edfa05cebcd3db60e2eb2b23968cc243ba9264d1dd81756f83d8e49f8fc669a28a436c3e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed7922882c002bd2b4e85d5e6454317631067e98298187c0edbbca2ef1008fdbbfe294da8a2942d00971ff3e89967671ba3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc28c156213bc6e117a1095fef54ff04f19654014032be0b4512ea0b10f611b1d93005a6b9ed6dc720d1f42bf661f439f8bd6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48094bc45eb94468b7c943a3d94897834e38eb2a6d4d13a192e26ba5e9db42b98180d6be30ad9586492b7779d150e57e599b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h437e0eca2219ff8a2c0671eb852dd06d8f3b77cf9a252fbf7fc818aaa04fd4383590090e740b90323c72c66c45042df760e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf10f5ed49d4e22a76b147a17ab1a1234c8a4bdb47c5a33bedd80ddb797f7c149e99c5b8429fae19447978257f8430e590a4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35ccfbd8e06fe07831c08e8980483060c45032325b0cdb63ac07df0baddc64f481d7fc0ffc8214ce2cb94151ec0c36ed0de1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9b672fee5ea3eca9a4609e028934e46ecd72c217241c6c263d424998bb9b3adad10638abc67f76ccee671d10ccef84ca8f1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h794b728d0a9f2a7f64778461d993127cd02358a81c22153097e09cbb9ea7ac2d89a020085ea9094bd46f50fc4b43ed1aa43c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h468a21d641635d6a77b5ab544d9b7a5aa5258fdce16f8a1215c1647fcc7ccb8164a6f00b181ee57a463c7d250d00bb5e49c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42b1122a1b38b118c5505add178b9ac369614f072f60946d158b76c8b38d02501be5d38a9217e2341b1a6fed22fb963dee3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda3bb879aee3275029a13d278afa58e573c313900141d359f8e028b485957bead323e56cd1eb235ad25e8674d9d37349435d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf02e8068c44856e8b6ffa79c1ab9fa58bf3776d902cffdd3535f37ecc712192b706e312cbe5e1ca31149e573c2b10b75cb1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8e76519302afd37e6d1aa12278dfbbd460bcfe076a0811dd9136713870ecdbe2f638338dc96cda99a77a2f3002daa5531f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec7293507b6e6c5e1aeb4a680e47d8ef537800f2f179bdfa7e5f904cc8950ae9a2c07c2cb858d905c9da57e227157a3de049;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb05eb78aa85ce6ce7e1bded031333c33620a514c89ef5ccb02021729f839ef30b27c0b3b7c041bae779e6fe5241c4ae141da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3b11d515a78eab39c3d0ff565d32aa965fd2670f607b8898345dc42948d92130333ccd7faada7da633132bd3191df1bd708;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e389c0a49118641d278b9ba51f494c7e36182273ab8aafe80e24364d5f3d86abccb3ad41638e62ca561c3a79a30dadb8177;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb78ae1c782680314e458c8ea728c84e51181f1d1f420a921f088bd3804bf790dd031d625b8a7e74381b75e5f6e74fed2c1b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8ecb69d3ee9233372f52e6e381b3bab603b8feaa778720ac6231c0ba5410bc23df8387c60424e5bb05864b9f61098e98037;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c2ca266ae6c2311d91e13558077f9962fece1cf7b80fd3197630c37c637663f8d328c72b355aa7840e4110398f748089372;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13e3648cb31137c95ec4fde485f524ad77b201d969ffc0ea8788aa933f723edfd59bbc244d223435e2f0b16246cae777260e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9faa89deba1918172e86363a30857bfd6257d77893e99a35b8fc7553bbc6f508836b15277fc86793d1a4b672a53c9f8245e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h982c843c6465e547cb1d354659150406342f3e8d69db4c2b9e10e319ac309dfe4e8e7964889362d64953d8bcec8e9d1f88e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfe2052e246a0abb7f219e0798b7cd27f2f7a6124085b378c8311d8cd1fefb6d3a4479d722967288d6f905f2ee80e0bb46ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b5faeeac6692cc2dc399c27e3a42ad7e3ba181a78dcd88ab523a77e5ea673c2b4033d01112c7f75158bac1d53c763c4115c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4c3739725693d8e4cd0cfa8b4bc294c85c061588d3d96b038e842b708375ad7a83e4759672b43d775f81e9efb53a8172ad2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21e7872bfcfebcdf24c1d737fddf831a83ec9d9684e921bf5d0e8e1af168ce8d55174a4e8f866a5027f6e3b8e754e5901b9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4aceb47e52c7da55ebfdce3760385e6951fccd4946cd1a9c98278ddd09ed700b0e6e759a4de763ec0bc42e5a90627016d585;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c167bbcdd18d9e2cc583d449f6c967a6ffb47377eaf4953cd10be9f75aff64fc7c2e4b13be661596736f847cfc93d5983e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c1ee301a3ed891a75835b1cfcf4beac630a05123f1b8a62c319caf297fa7fd20cf244b087ef284e73b793e1dc253377b7e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h880d86d74668942c40b5eb6ed040e4b328f353be326460c4f1b727d8f23479ab811bf8f23739f7bdfc555548be5686d0ff30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36df7e77136ea23cf55d1c3595b2e62b4450ac41244ca9a169e64ca54f93b16e6e1e2c6b78a2e36fb24c24a8b42ed7e697a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd897f7cf5023bc881b94414810d0f9f67b0a8deb058144b57204a5aa70fc7f3e189a8c7a943387d4e7a1ab9c86aa767054ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bb55b8dace52e4f4976502899642431f1f285c5cc1ab2f681221bf8f89e645595f67363c556248105abca34cc94cbdda46d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc730cd5b8642f5ee06166be7a137031a8c86a79ae2e2ae00eddf92245d662572b69c9040de1b6c5e6d49b3e81cb11157257;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2af57905a610e684d1dbb25d37c27272d8693307b57f83301fdb0f242e98d25e2cac24d70e63cb4db16bf9bf1964b6c0b044;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37015eb2d0ede1c6675db892a0328306d3a1524037c96b6fae66140cfb83294233f8f5b7ee5baecd48b9de11a2e1c46fb514;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f12027665a26a69a9ee376d73d0c125fc2819061919750f32edd6d36ef40ae8cb039d5c3444e4ba6d59010d1b36f0210496;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9838ce2cdec534fdde52a303010e99d5a21eac3cf30e26ab2b00178f652f1f885ea626c167d615b82a0a773bd59d9274942;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7d82a5d833bb989a5e70d5c8528ccaa5c718c63e11048aeaf9db9b4c617cb7eab403e99428b9fe97765406ae59b498ed600;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31ebe366354092a2b24ae31577e3060007fe929f9a9ff2af251b63452e43006adc37668953f4ac8eb5abd3b8fc5f895f26a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3c475c81c12655438810adf66114d3c4636d0f2b058f7f991aacaa15724cd27f7b65b6cb80fdf20fc0078d8fa71c80a12a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1880d6928930d4232a568a791cf4a85f21de6b79a73071bc8cecaa1fa8fa051b37dd90f3bfd5b260ac2e658d90f4d4cb6144;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fc02ab2323323ea25f57e387656d9c9eb79a85ac236f6b8ca79e1967d55d8d10359edb9af147f965e9afbe18dfbd9c9d6ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdd3ed5779a5ac43c080a89d32f06830a56d07125abfbaca1dc1e23d0b0c5a50c5516640590e6aa1d85a7397dd8402d5e757;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1037807d934b72c5b202927473be87790a4994a797986ed6601d69458b7a36d3c04688c04ec13f6b02a688473db612c65893;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f62d5ae706747d073fed965b7d70da92170a0b9d5c51d3901eb5ac7aa648870273c284fff1776091d153800978e8f0675cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaa6f98158d9a61f1f23ce68b9a50e9da5f0efd5368e051fd472e51f0a8031c1b660bd5acb8da571914dff85daf80b057991;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h772a6f30b7c25b66783a186a1676d8ac4ab3a09639e881ecb5a970853a3d27f3b400a22b339f701ff509afe01b8d13fabd8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bcf4be76a3a2bae5b5c69dbbd0c643c350a2a5c4649dbb90687762fbca6b3aa08e3a544dfc640a18200fca34b7fe3c087a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc5c47c9cd69d5a92e226149710a83008d266399e78bbc170291823a6e8c5ef87c4eecb9e0274571c7a8a1b3a0fc328418e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbdb86ded58a889d25619707107b50f2e8ffe541b31d1dec29d401a1d49d52617d85e5263f9d1d60607e43a372c996b27e27;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3690e204a4a519721f2a391386d516c37f1b8902eff0956216b95faec803cfc08a6ad9f8b151ef5e00173b60a62a0acff3a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd759e5ee05c7fa97db1d7b242e63a635c5e4d8ec7e0c88d157b87ef69ac98aa34614c1489cf4390480a0cb526009baf687d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7b3327e7d5b9886cca266bafef826ef482eced85acea4bae5b7db506f8077d901d55c9460b35bbe1b5ea83e6e74219d000e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h72959c8110c78d773b1c63a695c28e04b4ba7d2e99ff8d10a40a1f213b25ab868919890bb34b70b81a1b1cf0ea0ed1dbd1fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d17509eba6cbdae3dea90e933ac50d53463ed36fdb8348001de311be5612054cafe0d5794ea71fe4ab1dee734ff99e5de35;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8faf95180140d29d2951b0689c237a7896a1ee299601f32e1c0a1cb6689b52f975778733d93113a65b92d3ac156cc3fa8656;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he718a4e90c15cfec03fac6575343e59a230dd1c52367e188b0ba8746240ad4ccfbc63e677a457a672ec920b37d2f2733ff1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he20b4ae2bb1ceacd65759e8bd817fc0585470dbdf3f8a74ad8cc6b2ae34314535a58977c683f1641bf6a4ffa6971bde828ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54f198085e96e35d03343ec6f2e4d56ff13675e291d521642fd0d83cc3d0a2ff493bee180a6c44e9f4e242c4a8a8219b352c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heca7f4a487e71dae8b9b53b6470fe9a85ebc4a53fa2c54a2db2bad425abf98a7adbfc35bd4dd7545bc6674f157c20657fd7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf146e7ef3150678e35464e3a9ed3f0119ef626d46fd12d0d89083965b3393101a370fec0963afe715bb8b55086f0758b8100;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h225c9eedcfc8eaf680c95c07d17529252278cc747336a0f3e43d14930faa98a1e0c530d8a2df026bcf3ebc27385555745965;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h565e81f09ec1adb509321b01ca27a4c566c1f18989997e40e0eccce4b3811bc60f87a978c044410cdb30ffb7ec64b3213331;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2cdfd937d1fae82c79052ac89bc0b20c660f7a19fda8fbd1b3c334b927ca96c7f01999a8fce22a52f4c4268c07edb7a0b38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4535d07deab957389062f3b75f444eeeb7f26ae3441e8924fcd202d5860d435c2c4fa035418f8286fcd8aad155215d21f07;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec0326a37b89e3e53acaefd6ec27a15d58eb16aa2ba5faacb46d7f8907c1901a3b19e5d9f695eb8c9b3cf93f1a0ee09ee330;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b23ad781e289523f73db677120f1d37e52b1a2a9c7fd3881d11de2e667dd8daeef7bf6d5b08ab90fd89f05523c6d5227ff6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c301b91308ac7a687e37cc659a31c9a0f872dd11e99376b176467a72edadb5430ae203b7fadc48444bf5f4733f0799b1daf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc143bc2e229e4896d05b7fc34e5a4d458505db78907a2643ff418b93d730ada8671f8b709c325977577ed878af9432c65902;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19538a6011b333a79af92f6a901ce8166f7bdf00ff02cfc869cb6eaf3019d95ae848e45a784836b659c0e96478b400d7806f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb272d2431a85fcb58dbb65d5c2712ce7df16606f58f9e6dc3f8aba8946ea9a9bd6d373fae3b2fcac4b25b3844e24e935b928;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he232125bbf87ac023a2d3fb1f51363ef0593f702cb6bef2fbe59c92d005cdb66880128603fb2ca4313cb64b3b653f1b731b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce778e7d31451ee88a9ce987c3ba864081f8f0e47fcf8af1bfd097932452a49c249f8f972a3592ff098d16bb3bfe72b314e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36a7826b04bab281322b297b8b8439005fa3e111311512317dd7e3b93dd12a8342ec3e51ad3e55fb8fbe237f2e865c0fd7f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ce65bd37e6201c350832915497c07ea3829645e10e9867ce82e942333ce9a386cb49cb32709537a3e7fca0aa025746a7fa8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h859d34aad923fb3071d96dd88c01268cb498aa20b3bb862abb76069ac29fcffedd117abe3db11ae79312a846df957c081198;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf85b570d249f949093610168aa66795b292c6a14c0d28f55dd9d8a20595bf263c03adc93907a9dd50c51271deba1e76a14fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8aa06fd9299aad271dcc93c06e84aef31802af9270e3c95c4f86ba58db7b958a46c0325703353d05abac9bf1b7a044bcdd3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5544b6a58c3a1409821ca43f92ff5dc4784f5278c343cc0a29c24511035aac7793bb35aebde062c0a0fce6fdb2ec86fae011;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9688a97c1b9bf01693ddb2c532c9585cc2519c340de42d924b3e97340d764dc43e820e90690c57d87954c4d8830d1eabecd8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcabb7a5be0cabc1ccb289a289176432469c7f5ad53966d0e15cbd855ddd06ec5cc13a991da028cd411386b3365d8829ebb7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7444f10607fd59459ad1a989fe3d8d3fd2307bb01f56a1e61ebf29f870c49a9ab641c2aff5725c0541dbf1a195e22757b5be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5813c4e38a9228e56a77d22dc37de2af2def97ee7ac64c5d3512b723c34d943b17888dc9718b520f294260c362d3d1f343ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee32e4ed71daf452f090cc770ee5bec487b3af5095dd731899441b8a54c2ab1207eecdc9c8255ebac5dbd78775115524db0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h396f1a224084725a9723835048a13fa30b3af965cdda6e4325961c38169cc3c43d751ea3120e66e11dd270fb1d72bb0e4f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f60b4551cf466c98b95511dc5a244c2a8f6d8a37da73dba7d1d9deaa8bd53e824fde5583ec12fccb1d1f46e6f18df17dd70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf50fa07eca2f37e9898261c14b6f14e65dd3cbe6025a6da154d830c10459b3da9c80d46d3a8456b2e6b6ed9a256b9fb9c0f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15a718d07f554699b7054d51872c000f3651c0ae835745a57466e996cfbcfec202f81e8b05fc828df63e8ec647b68078ab8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d246b67564d97888f88cbdf3954c37ac82572cdefd948bf409ca426a3488a8fbd3d22a42fe9cd3d2a61b7292c63f7216477;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf07387776fb631684c56226ad64f383a9a2de62e7b8a9e549716cf5ce78ee87615cd9061c5952e0b5911edcd16ffdaa1a1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2611eeb47ad15ee8466777598acb7ead5a3dc8048d4c0221b24318404f4f0f6a0caa70b129e219b9fd24e79da58590c6b6da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf94b1ac6a8342a4ad8384a35f8b9f468220bed4ce2b5fdc9b8cd29d83829a93b7b7f5bda3e01803c8fd43ef8f4d27f6ce615;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82a2c392d7dddbc961f6fcc81127bb1d386722f4996976c86ff60ee0c7209ff172c2a5ca8b6640ac6e91a4f8271cebef67a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24b682edfd34f0e9e2aa5499c36d64711d15e1bebce799123278536c1ceba10170233473211eac5d88a7163758264a0df373;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1482ef8965b3e90023f6a721a1039308032c705b2b15aaeadc648508ebbfc27c6fdc62ec0440855d6d1e7298b196865ea3b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5af3fb6c2a870c26c324e6ea5416d3064bb17ca6b7f2865b33f392c4d8a54f7614b53ca958acd450bba8fd72ae72728a560b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53303bb1285c7d16470ce4d0a9fc28ee8e50f8aee07ae592965c0988114b5967e4f3768e94a9abf8f9d85d0f332b4a39bab3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73e8390d3847b2efc057216b1d05e10e0a7c4db9d2b999ca9ec6aae7cc30b8292ea8369c5ff6d8b9dac048654f2646a3ea1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31512581dac0bdced85b28016ceb66d3f22e608250bccc57d05cf801d7d9b6018df3efb53c53f3bcdd0da0afea3531c8c790;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff9c8235df7f9839bf7f32f840fc5ce1b6bb69db727eec8393d560c68a059836e32c001c2f843fcaa2bd5f80655f6f3e8740;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77de82fd1abd336822420d31baa094eabf4a4f343d322c211877f0c4e3b9b37431c686a21721c564028fdf8b818a8be3fd56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfffba6362a9c0d2dc67334b3a3d422b5068e394d8f2057da07df2a6bc74ebbc60cbef4fff7f683d763ce48818be0f31e873e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d94b1d48676a88cea34a6acf9405ced808685db4b182636c96a5ff961ddb71d20ed686fbdf81e8c67527dfe50204c385950;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f032e780c4e5b0d776207b9889331e32fbafbf17bee64edd84af35f54189719aa98ed8d3f722733210350d2d1b25e1fabd0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7accec8596630594c88325717fa09cdb8a72c7eb0e1cb82caa937a5490f13153d1e09775bda5548bb2834c7f497dee356755;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d8a17922fc957c951d1b6e2d5e7e3a86d29e463b1635208555e67ce1c83647987494b3d66046c65eb93b32ca371f363a7cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae2fb6bc4ff3dedabda84eb8d212167a8aea6187401d65926745a819ea803e105cbb40ffae5546606a7bc24797ecb96a2ee3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c46261bce2c6d24b3b42bcc916c77710a02b172e958a4f9754f6415a0b72763120b22bd4899389aee8cd2fed7cdc75cae3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h969af56cb16383570ffb83f2e5c1d12dcea289697ea832a6d39e38ee7279fa7bf582cf777f9377f8a694cda9335bcece577b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30e3b9b5b8e13961f219d0eafd318bfdb5e4ac58ffeed65e7e4bb4ad7fb3bc188b9ce75c452403f566993c581a640b85bf9a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h312ac5a7cf32a3e6413f700f5903d0f61011da251ecdfa4fd571c1f38b5f1658d1821a2e7db89069363fc20d48dadef8ef65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cff109cddb9ae06602772639d9cf1c8673b56bf5c4bdfa37edb52af59569af8667ed4076033d69907250ed327b159434402;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d68ca901a1464de50721a496976b1a76cf088039fcad6f41f87b52b860ef89a44585e713123290101868dc7dee3ab0c6425;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98d1e9a091b46599d1330dd0366aefdfe62e8091111fc5116a6973cbaf15b55ed9256bdf2708aa608cab7f927af597fb5b3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cb8b5ce7169dd7a8dcb8896581d8cb2b0e1238f1b5299e0882a370d8cf5c9270cb41461413122f2516d8167817cb0d395fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bd1202cc55bbce2c4d7e9773e8b588227238c196e231d0a99bcd60bcf17e7e1390674bb228d3f1e30108902550ad5c588a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha438be8eecc51181e24f4aa6529f8b27c1fe034ec4d6710b12875ecb0ddabaf59aaede8f834ce92cee7d0d0f1d11507bc14c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h105b06d7fac0b6128f8deeb61baf91942630c170969fae3c495b599f285351395eb4965c63e076a621eb711cc99b4a5c1ce7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h171e44df943ae0ee8b090d8e65085a4a8f7afd16889bc112d467da39a576c3b78dbdde7e1f18d4c706dece555e18d16d1101;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0711ac1e36a197f160eeb2e0a05a08a1f66675270a5d4f42638bf7572cc72fdb7525b170c1bc65df922cd2fef897569c286;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d18b70a5377b52b1768626c000b156269b91963c5d3d18bec41614516415db9a9d08d684245caaa76fade7a363188a05a22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h281c745dc277f9a4fdd0b52dc88180bf240df67c5cd2a33cce99c1c44aa018fe693722c2beef74fcda77437fc6ddba98327d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0d5111b7f2d25a6ee96f564fde39b8288d05a14ba2fa76eb8cb3da5b77a656b1a493c75fbbfee92a1a4360f3aa1badaa466;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53b5796601997f4e5b20df75a4bee0af7564289ac0e6b021eeb062c9490a18b5683eedec52d9bfacb52b9488a8e6d35935fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb80d92a998ac435c0568be0aaaa1b86c3016c209f1c734e2e14ba74be3f7b6188be7154c4a1fd7d42c8b55b8676f12e323d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cce25f4085f3f6584a5a5c9518ddfd84af91c6b1bc1b46dda317e6eb0e6f1f67771638822e86c499f8aa9010b38b95d1201;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31e79d2b287840fa04a5e1331c21342aa989bde362fd164d7c7648dd4a792811675beb0dfe6925c5eea4e7b14ce3cbef9087;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdff73ce8beff1214e9bf7904a13b21d9a9df347e4823a45a208ee11c1a82a6ab0398ff801d6cc80d5058e539e70345fb07af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5a07a84df21988ef07853775dfb09b1b60db3a856ad4d27a74f16b07fa3c2119fe8bb6f7c36fc2ee41edca5b1185e6e0558;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5f99eb98a027e5314d857d40446814e064a2ab03bf91c9300fe9a2e71ed41da8d111c70221c85c54224f402277d197b1a86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0b12060b0b4f8f77c4f51bb489467a76c5dfae6233c4ed888dc5f8582fa88ccba1ad4a8bc7fda07e421c99026c4d07668be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d73a66f6d66baf5da6577c147d8b93779f8d2f84b1e02e0893610ddef289fc5fadde50d609264bc749b2f3dfffe73c741f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb45153d4e834f498b0d5cdc5468bd35eab1476ddb7c3a1c9091db065f08944032dde5bb7aca0f43408234916cb440b74fe33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha405884dda0a6eb4fafc8dbb3b6e49146ae958489bd26cd796cd7daa3b69497f075e154d9645dfaad13f03a80066d7a78266;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc7db6f62e4ec7c1c988d2c030f536ad9f890c9ae652ab33997a5337b648359b7d598496c530373f0f97f7bb2851ebaf9a52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc48c8697e57711cdcd0e019c1b188f9443f4a2ce2ca0076ffb7c299c07ba462ba413364124d6a56f6795278bac910de9084d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h211fa968d9d892d41a33b56b9c5e9d90e8607ad2267c723d405ad68cf400dc855d31860f9c1206e2fb16dfef7a2cec46c54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7decdbb228ba0c20d7918148c7063d0cb76544e2bc13ecc678fa9f75ade0cc372e03795c96e3d561a4142a50b46b639489e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f646e287d685f7e8f6b632d358dcca481ccfa6806f91dbef596d20a0a2fb42ee01205b955c3b20028b071532f33b4a1ebfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64d51bc2de8b596fdc31323264cfa28eaf9915131dfb773f620f2d32c06a35edad134679a45b57b9a10f0d515de84b1648d4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6770ae74e1abd9e879cd8035665a5e0c1a037dfa825842980719f442844e2801ff5f22a78dda2f258f114cabad5f2b6fced7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80cf74c0f4409aa327ff1e7796b51cf4e57d99dc815839942cb370121cda866088db1423e05fe0153b748705466064538e43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47ea805a5cb64235d7c123f7cd2cda00caac4f9d4be50f8443d73ea9408a2712f3a590a073c63a54d6d582c90cc2acf9dc56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d9a09089eb380cadafe49ec128efa2a039737e1367043fa0af5e7db0ad7c902395c151fcf931f72b2da0aa06351412f712a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17fffa90ff53408b1a9219adae84726fa0b2d0058c159824ebfe10f1c624e5cb3a04e9f8d30bced48e83646e60940359661e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had2d4aaf7a2652d69bc3f5ffbe9a56aa23fc3724599b8230dc6034d201af6fff5911163dfec85e41379fbfaa599d9ca1490c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d55d0adc7db228f8abb9572966962e84e12627cb1687fcabb1195ec049e5b2a19453c397602046e6ffb4db3ecd224987644;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb64f07fb65bda0c7e72856e054669f943eb2d23b514258eb1041f5bf2e26baa639f338206f28ac5265210fc17cd94c82f2f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9248d4c126ace9afcffad11c47ec6db75c12fdef5feee1b14a682ebaf36f7e0cd8b6c2c679851e7753ecd655cc009acbdf1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5258580c73b6b6336584b9eb26dc57fcd93ad342340727d461c85a6741c298bf6fb1b0391893fae88f1bb84eaeea5c3370a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea569765d97871b72308f42f100995d9db19ad104bd50b9daf8f197710ce5faf069dc6ff82ae58aaf9f19e32bedc994fe0d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28c36c08e6903ed9b4dbbffcea2c5ed67a4519198f196cb89ba1f728de83ac93ab19c6620aee150b9dabdec686107f130bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf855d567c3195056597a51f9cedc745cf9768e05fd05e20ba118bb69cfd1917dc0f0826d1331670e35415d4d6856ba2cca7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4e0a96d0ab38fa8eff9d764d48d26d6ff802b5a0ba30fb80ce69c3f1eddf488fe47c127169da25d28f61f859af4d55b48c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h139d82d25b49542f4609c1ac536e7ca9df2e7e2967f307891755bbec0b2b5bbc62a56b62ce51c86ed4811e12391826dd67f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8934c1af2454ac659b40bf9b824c727fe32f1180cc92af4aec1359438d307cd5db45ceb932e4ecf67c0b9ffba922912e348f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c3cacf033ec7a26b802fbc0111db5dd377a9d61f8d37410e23f5f557098a41201f012f11ec79a191507d37a60c839413c42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe2ad44bc1f30efcb3a94732ad2afee31f8fc3b0d436b005164e469581f1a656172d7bc6ff6f615ed26f0e8edf19ddac82da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd83be3fed4ee97d8c058b168dd110e02ee533a7cb8730baa3d2fb42a1a4fad2535f85ff8eeeb3a8837eec1e8e8a69d2dd085;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedf56e6ba2a013a7524ce476c75651a3243befff4d05fcda21c99970197a7ccc0b2e2a8de2abb911820620faff5182cd44f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h740f159dc21385641ecd11be3e5f19ad68d7f18b0f17b46868414f2e163754325bac79e0122116201e7d83744aa0ed96b227;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf68c04c5bd8ea254230749bd7d2932f8b86bb58923643332f71439ca079722c04e5a6f6052948582fe7653af9800ed4e0195;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha497690fda29eda3a2a4e97248f6a474e427f48e78abd3259283f63f139ea2363972e1dcc4daf9f07aa106cc389b7e8b2253;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fe7f068e7ea3f702aecebea97bc95a0f9b9bcad768d6d3943c178eb855ceb2a03f1d40c2c2632874fd8f19bb8b6807bab1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e534666d2db4e43523e434db5dc4c9416ea8a1e544ceee19cb1388d412e98c7ef391cdbc2547f316706312636572b7505cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12829d1c64d7d5ca03dfc01c7fa37c2c4ff0aa1eb0f8d8cc20575c9c9dc0bd9ae5bd2c968a97c223058854836d9d227a468d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbea7e3142ef19ffd245a0703cb93706125ea60d00a819fbd66587f5631a3a263300ee307b1a471eb73aa2eda200e4d67a2c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d26abec7d9db299c8fee8c0aba7d6dea99cc33dfae7fe000b9825d6eaf6d0351eb4d25479ca945b87702014ec46a00f0e43;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1806306b479e7f7793a237803d9fe1b9530548b3b6c8190c1344a14d049d9c286043e3e1410d17433ffc3d72ed6d062d7545;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1a6c317281d383f3e659c34ce19aa8d2a18754c35683f8a2268cc38976cdac7ac1b2fb1471bb1b1e30e56682ec42ca68340;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9835826ba60fc49f50b1d6f708b5f5f32020c24531b12465d9fe0936684c29c59903f83c92ce739c460971a3a2cabf6ef54c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1a77bfa36d378be197de97ba945b7a67e084e9ddd070172451ec66c13bcaf2d070cbf3eb9ef06d8eacbdc521d1fb7af7465;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd2a5a40b789e9e255d51ef99566dc823c08e30df2d8bae6634a8758a4ddb31b0d2e3ad776a0d392f4e880cf0317da911ca5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cbb0687df4d46cbf4da9d6c5417f55624ccee1664c8e4706734185abba0afa612b7b588fe11955beeade447fd67a0da3c66;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb493b050a7840ac848c30cb08bfd9d5e1df566ad7476c1161bef64c3bd01d8156c923b33ccc15a99ee405b095362604192ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15802444ea12ab437bf62cbad9c841db5732153c012435c37b636d9ba545b4689411747338ab0286a0cf46cf8ba099d90d7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he80cf6f0df81f6e58d5bb1bde7c3c7f3aecf721c6165e257f4f31876e449d4b2c6c6e2773ab9cd3f3335fcf49ba41379d9bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8afb1977c3e579f7b06ecc4e8a4f78efa052546aed770423dd7b2f080681faf969b9137f3438fee331b3f5600d3a5d153ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc64456f64c5dcedd1c3a6ca1ca66121e32cb59bcfad00ae79c2556d3669a4a329217e1f6eabe4ac4c8d0781bf31b58f56476;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc8d314c8695eedcc2440995170c9b8d09adc704c49b3e7937cd45196ebb7cc3a46a5d14e79535a10aba8ac47709312c9443;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd72c6773d06ad7f3984460f94e36e98f90607e540cb63b284afc71ec1a1ad9589435758ee3c8888c2d789a37c8449af22c11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7ec91eba2965942cbec64463a56ad066fab6ea8a3e3e0b497ecdf9b41f832f03ba23905e27525a9cc1d4bdb9b83cce454ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b7001ab562459a527bdc4ee550f072c13ad2b7e2f65b67275ae1573ce029a123e718bc09959f9acdacf124ccc2bd442281;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd512dacfaeaf3a287f6063759175412b3ba7675995ccd11e5cfd6d2c8e3e257dbaab2bc80fb35d7165e04ab3d4f46cb3833;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ded66726fbb19eb1c196fec28bfccd911e2ed0c328f64da57698d73823b28067278b8f4981dfe8dae653735ae6c3d4204;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h873f93fe54788d249026c5730ed51312c6255ba56ef7b09d299bd8e428069c7bd715b9775709ca9fb1df9e09f116f8f56aff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h268a5a81b7f2c19337d5e461b32c7c487b2d053601007f1e0578a939bf0e53ed35dc637b5dff50c97bc657feaaaed88786cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cf4d433fb8917492787b18b371935c5fab57085186b4f24f1992e2dcb1c848f20d2d5842982b8c73bd7028676ae4e128e76;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he730654c60fa5282564fdcfc543163f43b771ab093c942c139a5da2ccc10bc14449fc4b9e1a6295cfbbe5d7b99fa92b0e24c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ae941f7677375ec9eca6928fadfe31837887c8a340d4f4389b91240dfd72da35d9a40921dae9f9a7f3f199a0a6a68718309;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e2852ebd148d4b476c2155e4861d8f82039398071c5d75c3a52b6923cbed6cee732fb11a70d08af19405133dd3d22e94c32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf64d05013e98d5dd0f8e02e5fee23b7cab972823ab474d1bf9067e66bd560ed45becab0ef49a8e419e376d7bf03e09a0824;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55d8a3aed838ba4dce53d0c14481071e58398986ff547d0b8b01590587987fac6b877f97021d7f9deaa8f38b19de0c8e58be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc7add771a883bd6054824b2020b292f475d09ac92870d634e1f08e047d902e937fd1a7b19049a3d116da9e0002399be6f68;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5999577a06a86efcedae29376ec2d6f0672d3bd8ed52b02fa99a68bd5313c602720dd1408d08c25767140800e24325a99176;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h489f0356d8bb85f41fb41c853c011b67f8c7c9b7f36b9015c83b846337a61a8c916e3cf307164e359cee782d3603dfa63315;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13326b85b3c3ffad0928e97509ea72cb44ac4d031e23d68c70c46acc9ad384f5f1275d5b0bf4afb25226045d2e5095af6484;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h166d6bdd650ed7115c10670ce27437e8ab7924aa8c1684b8ec4384a4dc0a68e09a19978a465ae0b1fb81fcc895a589ad9beb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbff08b07d3b8b077d9df0ed212eed6bf41161dfdd4b3c83b396600f8120d1e4ff56d948c78b172810b9c32d72b026a70b99b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e83e74f8333c04fff9dd8e48395d8d4790f2824552268779bc3c06bc92cdbb50cbb2e64d956c21923a6d68a7e0ccea45f4a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he557207e8cd46993ebec08e2e99ef528bdd15b90a9742642a8d89d5fe4554e3746744ec206f273e992d833ecf3d44e2b6ff1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h956ae90b995c43cfd3f967caae8deaa5d17451ad106f2ab6701ee63439c2ecbd3e8f3e6f0a876bef1bd474328654ea974cd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37738f2b1ca01d839af1ff34b936d7f16f6c29bfa1cc13e240b4fe231ddff497b266069a72d5356e2e9fc1c54c0e64f32eb6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3f3225921d13b63119e7c20affbf80c44226825b6e73793cd41fe377866e08c3d9b5bf7d8efcf551833dfc794a3b1fb07b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0c111a076a5bd6abc94ef74988ce64a75e691c97a743c7783a4f14c4707b3aaff676d346d3212151aad4328982fbe9fa0d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcea9dc5061685fa52f688817277d2ed2b0381859e6edfef2bfb820122538b1dedf5b656fd00751bebab3f38b87fac3b1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd522e25094c4579cb9b2a26a4393aa170a878690bb7da7c2bc90ab15a2ea070f1aeb7b2d6930384b0ee6173b5c2a752d0af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7584eb4970cd69b34bcf911eee63269bc94b09d3271548b9fd179e3ca0317f79e2eeb721578c0d3194840cb07d0b091d508f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf2604da4dc3166cb057fdad52612f0c165945bf6bf3c2e20436b60222d1edf897ab49f8c2656c85b961a56ed03cd83fc54e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc16bb5cbcc166dd1e4a21aded53c28156b4996ce71575df90d6d0c6c1535546e2f5f73396600f6c8f8476306d2683b55ddf6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb65b4a4a11ea5233987daf4dc927d2a94e8f500f5f6f2fd336dab2795227a292d1e911e3c73cd8eaea180905597063676458;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h619e7e2c7979ffee7bdd1304cbe3d28dcf1cc1d43f3ce77ac062e40176bb812f64d852a08d7c241aa13eb9b5fef3b9350ee7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85d40dc364ef471a382b7a434dde0fee58e3a6ca3a8c7d3183fe52e45a6fdb7d229ab6b957713ff184532046dd0d5f186175;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4f7a2d61600daf70186485f7889143d6888147f0a1fcd9cac40e89d177cc30b04bfcb71a86eadc0867f82f9208ef43b707d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ebec26fc742dca7ba0fa5d38d7ca36afb36da563b3d8f39e31660972111ad1cc32aa9c540ec7a49771307965222b61f8d20;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf772cfc8e3fb165c6a0a8037515f39f7d954c90345853587f087ed0f7b0deb7221c0db4c00623559284ca101aa0838d793e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e5389660ae0283463a58a4544d715a8c2e980feba32e12c4baa9a7f8231d42992c7c59935de88badfdce2ea56f114c3b773;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59a4271dbf9a0448d7659db5bfa31a650f1415f6ab1d9c884719ee1e29257a5f1e6f920c2d0684b005cb8489c9cdd080d644;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1b86785fdb1b129afd4d4e90f707cc85d45509006709991bf7dc2882a70473bb4f47d1f02855e4e3a699dc56557b6f95db1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ddcea2762a32d3986af0a63c336541164cd283731fe1e15088ed7c78a951ecc9867bff4803a2f301bc4a3990ced46478563;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf086ecacea8a81ad8af48b4b236c1dfbbb8c453d853a44427dcfb1867057d87f31cbce2b87015bb8ca60347bffa1b115a5b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c50c4b95b19733212b0228a7538fb23226ba1d1250aa8bf3b7e804c2fb7d5d14cd786b22f9f00c7650bf777d9119c44e8e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88caa08041d50b8c0952e1b1bf6c9d92a97d12d5dc803dfc8ef194d9a22c9348e23ffe54697dcd353feda12b39282bd58624;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34220ef6c4039a6fd096011b02c7c6134e87253ba7a2367d5bdcdc6dc4f9755302cc9c64ec5bda906d74e92df61ec284bde4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadffd64cd9d81f839014ece26c8e88d1ec102fde0ea1f593c872b6d8b406f410700a90af6f7497e1ad7d40efe9ddc0f20cd5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25718cc2cdbb93f52024eacf642d0080655bb6a744ac2ddcc791ab376c9a9ea67b58a593b670a973c372393e065dccfc6a2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed0e31c0c9a3dd81fea5e9d23719d4ec597117168705e84ce4259dc109f2f9cc5ccc1f740ee4bec6983baee5d9418e7d3cd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb75b6b71da2e4e717591272de340252421fb42af6d5730d67818210d1c52152c9917782ce1bbed4212393f2b27b140d8a77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h895a9b1761e38560bf1d60a21c44171c28bc5fd07d1fb550c23fef5a8321db58c79e99c635103c648af64c576c3352cc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha218687a6be099cdecffa09852cf58b3a8877b975f432eda7ae284f197fabbc50456490755ed3dd87398d59d39e2afc57ab0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he79cd8101950204598f76c008af3f5dbd95efaeb4022e17134c8b20871ea0faff6efa730d1a5e9db9c98cce260e4fdc929f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28ad5b3f3b95410b3c6d1d84e441fc98d967b131f3f7f8d89ba8958d8547262a30dfad4123ab9338f6b73f6e80533e21ded0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cb41d3de0c9c4787e1418f1685b1000c0845534e87063c7c9d8ee2b77e3297a4e58c4d5a824b5533576ed275f405adf4a67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha063e324392d82025ec184db8e6c2ae4175b51bc15943a3b46dde9d19a62f541c9668438dc09b9b645d7adf96efc0108707d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57d8c445a4d481457d935fa0f3141b33008d26aefa802c9fc769432ad5531d29fccdd8ea5976b9951ae2b2d0cdab71168603;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2ad662c191b06b0e48c2e98e6e18cad9d9baf71c75b1b7526af136874bdc37252688b84624133c2074d5d37221914a9635d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65bdf1d7e80062d9fa351a3b4d8ad2bb1756b39bd3ed4c3a0d2c78f316d435deaa984e474747e60d6b663e6c03c658644485;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha66b1de792a52dd9a067aa4e5fd7d254a31b759ed182bf80f46e7507ed3727afdb897a6042cf4a03fcb8d6569510d9cdb4fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9d76b30f64b67be665c8e0392e107292ad545cd3814b70afa93700b03cd75fa8db1dd9d2b947e0b99d80657b5c723ffaf2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16a62fcb18dd63dbbf6f66d7b0aec653deb650a47cb60621046d12792aedac48489479662f768c27909cc4b5e63b76037303;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b1a58d4684cf2a7acfa2061e9525d383da45bc156a428919ab0c2022aad4f870b87dda661dce95856a532508c2fd1137176;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7890693d9224e03a5b52576bb5e106366f47a4349bca59b15715116d9e5079a6a4169590af34065c8514fcc409873e86cd3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8def8bd8c86dcbd1f9e241ead417227961cd446e7d270b6a97f42dd05f625f292598fba1701740f82950e51cbc9846161a81;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27ad812627f59f432f7eab608c1c75064de6f9b0736c2fb9ba9c98bd85a5f936239d5de134e08f6d3cdc392ae2a23cf6e56a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c444b6ca9a6c4775803717cd439afb4b06da29f54368178c98ca79b2e2f040ba2108fb4fc27d39473e261b842e4dce3c49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce558dfc2ccec94c4b41fafecd688231584ad81137b310b8a75fcb09b6b8ef6f312eec2111e5d92ec5c85a4ed2d8a4753103;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab7ac1d123c0dff65a2438f0e5555e0a2517587e1e48b40dadf6eec25c970c0389672abac5bbdc6b72b4d30f25cdc40f27c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a7b3dff4b81bf4736540f13285d2f6b4c7d3a7b5c5ee60228e834772aa39d7bb2ef42d0065ead603a8579e298a8a98cf767;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25300c5d5e68113c6bac20ef1deb75472e2479cb05fd32cb9c42518778be93f3b5794a85fff2050f2d169ea7f1862bcbfbc6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31d4210d1120576b3b1050c66ebb935689d9fe48eb0cf5b62cc1e014aa2bc4357b3bde5a0c5a243f2c3c0c6f29be2d1fe87e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h111acdf389a6b21c79d888a8cbd955cc64cb80153d118b33a3df3e23002d925fb4baf9eb42bc7d308f3d2aaa69577f03c055;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b0c4aba1c05bc524f4683724fe668ce85360104c92dd7ec9aeeaf0ab6cefe286b795b27b78d3f416bef8f52da958f38ee58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdee7fc2be0af6afc105afe8b1205a6f56a79ef8c10967d2c09935dba797fdf2ccc75efbe0f98321fb5e1af83c7833ae264f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26c1999aaa2f68e3186a9fa3c0f1a5242cadf0209585b0c0bf311fcd335a721b70351f9c8bf2d8244128041b69028c4dc0fe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab8c77c4ba045f751ae11a3c5a46d19b4aeffef183127ca2efcfe829d87890fb791bce708a787b872c05b1f1636f0fc9c7d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b6b75f5019c65ebc7bcf9b44983297a001811340199e82321818252e312e16ecdfad50e11976d97c6b6b022c02825f76b4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7f72d7fa64aa29d8d55224f9347db66558551121e5d41db2a632eec26ad86069aa80b004bc5f4dd09dde88a03040b0bd07c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bda82eceae9b44aa522bba6ada16edcc2e38ed4d799d1a095f7facea4c746e6762fb8eb9116f9bccebe50f13b0b7dba3025;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13df1b24f4cfd9706f28ce08a1a5ab39e61180403c3c16c057c5c6aabd14f26c9a0bf9f4c7e2b6828982a74ca19ea8d0938b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bb5aa2bb84b8a29feb9564ec89e4b41bc79ee4c66319f02c808da9b95fb74a6802f609730be3470ee3c1615aa93547abe21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70e2fb1ae185afa2d34b31286a09ec1a7115ce0336c206139ed861e7f69dc4e944ead650070c6516fd91e5df1827af317974;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd1318c7d26a16d56247f05619402a49e22fad2710fa5fd4b2cb0575ca2211e10993ff431d0e8f6534aecc8dcd231d88ab1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd07864dce13cd074be96d0ec37dab2af9807978282cd42e4a4848e1c69897a4c62b63cd574c9580304eac776ab0412711e3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9614aacace8b1e0b0c9b191bb19e75fe9aacd864ab65029a1592016297a5ff00a8516a5b1edaea48137f52eb175e1e6a93d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5859431e40140dd4e13e2bfee071b95d21e645edf4ae40090284c60ab792e9a86976ca32ed392ec5a58fc70a3aff26d541d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c813bf6cdba64ef5310a8e9491eeeef6dc44fce5add31d385b81f98d53b75118d88a9cd0f9c497b1683a32473621fbffd01;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h708567ac514f77ede0b9521b73e62a18f030a06055141e2a07e357a1c148948f75158d7904bf6c5ba42a0f8000bc221add15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e34f1223cddf4068dc85ed620ba3761a10f537f877b7c93b1b2ed6b8d96026ac2bf5c56f07dbbe3a307f3c180d52d4351a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bccb8b9f2d856bcf8a7f70cbc5582bf7defa53f2ce130bd788b25a62794d556b00a30d1beb1db9a63fbc190aa03cc6b2459;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1d88fb35131d50543693eb523a4ce38f844252da4dba5e0611407665b9f6d9b7eabf32aec018e5f1c01c0a9be90e7212de2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb037d1fc57ca95f3b768064beece48dd0185115ec50d5c1d2219c1feedca27ed96fc256653cc0f5a6c3a54904e8333f9c4b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h788ab99886b26d70f32e2a386b126e5d6b2068629f2e4ff1b2df08450173e383081e40d177d691d24f164133224f8d52370;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70d40ef0dc373a39449ecbafe6e4a01457c5dd6f977b5e9905b741721369cea7b9b53abcda5da3cc43df2bb09a82df790ba2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78b7b25ba6f16d1a7c5bfc528ee7028e8492e60d5cdf6519a4cdedc26c413a0369df016f40d21165d5e2d1d08542f44e5185;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16d26d8d65326192f1077544072445b03c0583acd5f74d751bdcf7c6212e73d34e87724c0fec17c2ebfba5af2ae933671ff0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67140678c0fd2dbbaa2d3f547bb82f8540a9c387f821ae22d5ebfc98485d7b0f80c4b879cf80198619af869006463cd4017f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d2c0573a704de30db13a239874ce2e33e371a09270b35661069273f7501d083b781dfa16d84e76529880b46f36a34d9d28d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ddfe8c26a7f48a07a014927ba164d17074cdf8ba9b875564561afff1cd1eb38b57f62a704f22d7949c7dbde251f36df8285;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa837cd3962df2245598fb9e309b1d16076c83d9c8bcec993780162a395780b3436f627ba3fc20fa9b47c0fe159bed0b1a74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79fd92fe6a6e039ae27055bb59cdbf7b0d070f8de2d2aec74b9458681c32c195965ef121b34099d6618e257b2a2d78052892;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc68d072be8f4d8137f8702f34cadde673bb56638b232ed3c549b704ecb5a89a5429b35ba725890b8257996dd938a76d0274;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb058ce2b3bbccb5e1c645959a624e697697c55d5e84078fdf8156f9d5b7af9468d9fb9974c03ef9ea2987eb3e2fe99e6b1df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca6fd7421afb43e0f7eb3463b0df27be4c9089b254c79de07a74b7315ddb2219cf429364778745f3f8d8361034e6a2d6372e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec65c807b831203a1cba3efc365150cd148ca4476ebd8761f28cdd65bed062ea7f78b402c59a8ea1bf8300be87bdd4648a89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c6c1f5cfa3e5174b6f3befb8fc5692584093810e27ed1a848c3fcd8d86d3523e7e188258155b61cd724ce01e0d53a697f69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca5de183a055143fe4500e3e663233997c614eda2793374c2a7b77a893696082bd8c1db1506c9bea253b4a95d66316739558;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9cc6fddb5024c964bbf8b9397c73b98467de9ce1d652a135c87da05194e70581e1b7fe14e55f804666d52b558091cfe918;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha69de6befc936b99b708725b9b9bcbc9d013bf9f7fa965fce5c13dbc36034d8a6e7163934d7ab3f386fd5781e64d1d0c6fea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2a88b8d4991691e275fbea34685eaac2c5e85132d23b615b25279d4d4ead9794fd41987189608d641d71d14b226333241e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3f32b0f23b8cc3e3f511c44ec0c36f69539d27fe60ac37a54be952fdee08a75b68233b4bba2fc1a0945ad5318b7e21476a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6d34106aa3466f407b911542530a8978b80238ac99532ebd6ec4f525878456a4cadca58250b887bfdb76b398b2b6e7cfb21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77a7c595060ef3c076d76c89ecfd23dae795b00e0230010d17fcd414526f8e4faa37ceeb4bf5eac8409a953c1923cc4212d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc279e8b4c1697a15add5e83ef20d48474c244636f23cfbb35ad03778e4ce0b85ab911a17d2cc173c15b0fd8b1aa05d13b11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef179a9dba60f6b8f7d8e794d3a59b9bcabf88be43d41f12acc7276f374ce20f81a13754c2beb6299387232919c101a98027;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15452c4b154f1a532b7b5869ed52190e88bbe31525f468e5f78dd99ad29c8c50d53518f0ca97fb22316128e1f1852d289b85;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0e59ed6dd3e50bf45096a8d29cce1ca49936a9faca89ff032ae5ab7fc386cdddfb8c0c39e13cd566fe41493498eb791fc7b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd31eb8e246aaf61e9b27db62d732b9924f796c61a233bde4f86261db22ae8e6ba4e5a89c51630e81888bd8f237078bf9c2c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h946cc034f31bfd67f004694c1e253b5a767a36cb86761902d46478ae581c09914bcaf168f2e895c0a85f9e9e2c1f7e338581;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcbba8861e6824f582a7246c2fe20012b33d7b9c5689d84f98d0ab99ea187e0ae0933293ff53f84ac7437b4782232d15dd95;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b56a1feb38fd6418a7135a256a6c7e874c3e3eb893efead26a613c29772f7e4f47b7e46d16e70364790f805e4cc96db3e14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe1df306ea85a4da0b5793b8770d6809fffad4b584a4dc2427661fccb8a9b9895ebf1e33af6dffd822a4d730a1b59eab1fc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3add778f1f2ae379af08b5a268ed35705f9a3de086fb129f359cfadd2cd7896ca385319c2d09b43078c1ee14667d879bfea9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a46d2b6c80c02d6fcdb49f5c486f852253f02f7b8db5a953d23fb6d88f900169232537a45ef280715045d3d24df4f76214;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefe368110864ae3e6e09c4e2538d57d0c92b7f76aed543352413ef0a8f651a90bdebf14adecffd3d411d81c6c6925dd07bd9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16b7bec13c7e493e424df804a59a9e0b35f38b1e1bc1c1bb193f49dc7f7d29e34b3e8029c2a3a85c4be685cb701008b98f7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4303e8ac2e2b08b8247295e9a39f025ad42dc1b236cc9e87b7d5fdb5b5a8a0cb69d4044256336dc6d4476d8c83d09bf21b97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bf3212f2d64e0fabb6850c7051e723098269bdf93efd28d59ea4226ad86ccffd76c0d68f5ff93d7bd0a3a2af301818bbf0d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86a4a0fdc277d9a796ac0d0ed07c954d7ab1f9a5506f5a1d982ed8ac69e2ee631e208b866e78fca57ce983f224248d751466;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb020f5eb9794fa10bd20dbecaa9833f5cc231a650039aebe5fc510bc3f677db05dccbcb6f173a54b4623725ac53345780b77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5289e73634290cc07e066b04472f99a5acff5b073a6de052957df98d64575cdd004a62f3941143839aa7267e21f99ec9efc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3904cc7938121644c14727bc9889f942880bc6877870f350e062adff3b826be8eea0706482f86900373fb6ce5d5edec32f7b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7ae293d13919c505d92c2f77f8d4478e7e93a105559784ecd8ff56ddd6b84dc44b1e43fb53bfd478c76771ad6af88007652;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h843d113d8173804c06a215996d303fe53eeec5bfd693a598eef045c0a5b9e28bc60e35e9dce05f278a868dfd7bd06688c05e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heacb1309f838eb8195fcce0818cdf916c2bf27ff9eaf1576bb1f8e26972aefc937b1ae4216e5029c1c833794902ce35e6584;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ca6f33b1b50e9a1af38d507e027b26966f7c3fa561f2881571114c4dd279f7db6983e87ac5c6f7e95959a2aa4cc0fa434e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h81494c6b11a9e478c3add4bc1668db909ba5938dd4297262f775f62f902ed8559bcef5c21b98bd6a425f8ff8e731609d1dd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc497b1ef083c5607eb7cc909765d8287697c945a08b704d132448c98e11ddff954a24121c36026b38cc5d6c582efe172ba3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82eb24ae85c66224857217a99fa0f5bcafc085e9cdf02b31d9955c2b8792f22b4c2deab14d3752a0e1690446987b15950b40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd8fe608a371d4f4b77a68b2e19055663d722f08e84a21969fadcdb2ba71cec614c36d55f13588000a4abda7373621acd434;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0f628b7ae4297bd8553842f260e006cb0b338312f3ca20626b8be5aca3eef24c77b2311e8e6a7c9a046395629041fad0f54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a2eec52ce5ca402eb796bcbc48146355ba40084e0652fd7ad298594f96e991d87f77a773c15d329216f3a86e5f06881e2d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe126240dcb214af8551c3e2b88b78d18c2fa289c8188e863e06d74a2f71977c72ed1371040495530fdfd0af3d5178492f46;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cf649a0ae9cf4db0e8eece63588db69193fa650c71ed3a1f115e53f9030ab0d134de507eb5f7534ab3d6d47f2f2c1f2abd7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4b958ae1501c1367a5521a02b2bb7db3c173c79f80e4b16ff30cda4fd6d8b3bb93d0b4f9c4ccd0fb823439e86b5c456c852;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5a24824efedef84f93dd47f6b40faf57e24658e57f6afda4df93a054fd0c68048f176116e0eea4c3251bbfb81782f75a738;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haaa0169aa2b3feebcc5c58f548f6f0b673d973fbf8b76ddb09af0bf155b25225ea4048fb004b583eb5105d10b6f6dcb49766;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe339a31f24bea0c7f25a085c82fe6f0913eac8f57e724a0359e05e18a2ea8e16dfa7cee65a4d0331e44322bb84f8f2c5152;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf22390805a360f9f99ce3df1a460b15367fd2c34f56d33abfc260275b99247f8c6b721efca4cd26b4e5e77a7cf1601bb4572;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21d9801757f8d4da3ab75b3c258b12373911847f53070d4cedabade76d4b54f8e890f5e484dbc6ae2855c7f0373f3b40a6b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83539a59440c4341d6732eb4adb71bb16ae93c65062f1ff874ab9e75c444494626dfc59eb3b8649225cd250e5a45fb213a48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dfa6561920b8dcd5c31416d0974fd3de8480366d857553a45eb503ecc2266998c13c5f4d3cd8e12578a385a9c34afd6ec10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcca9c95c6cc7ed265b4ad19963f4cbfdfdccc76626dfe4838e7c8e91bf26035e144132c2beda0440987e6695342d09acf1e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2deb3f55ab3a301788ee8e0e1886bf92fdca7487e7268ce61bf62e05e71974acebe2307d63ed727b5bb8fe5f2527bfb5c24d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0f6cfee0546010b59ac349ba9da42222efebf9f6b7bae454e025d3ad7f00960dd39cc459281415ab407e2344d61fbb63fc4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f7e2a32738b5bfe1ce3f55b22d468714bcf5e8866d8279ca5525461d98cb37dab8b8137498c7b225f81f4a7eb4b4523d374;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd19cf7e6702a93027fb0891c96ca080f806499bd2037c893f50b17acfcf7eb0549f7dd875bd64adff23ad15ed042f0295ae9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02e5db8fc5f30a3a5952b6bc2f3a3f2ee2285661b332038ef5869b3a5652997cc9ad7c449baca63d9eedbf7d105b52bff3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb87c6499fdd04261306374b6e05a63e411f542cc25237eff16afdff0e818cc65c4c631b5b9c1b10ee89674f7861b02347b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdac6d7499ed00fa285d51139c99cf750f2c16647c49427ead054f280692215362b0857dfbc65b3ea1ebf6dddea735bf2932f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbcb316d64e4f9c6691aa59006a585d68d06793faffe3a00c119fe2ef0f8614440e00358e72a381720af8b3e41759ff996673;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h585b25c52dc9c23e3da435fca3ca420b59271c3091f9230ac97246585a93ccf83c86b2efc4c66cb740dc0d62178e045651bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcdfb1c877dfa4fb68fd8c47485c0009dfc42d691abc80379725e08a508eff1dce22097ff93be49b099e6d9ea12aea516716;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e29d63c01ee598c29130068e6bbbac82a18645f2cfddf5f5ce23cbd178793e9c670c92349d646c0c323798bb5607bc1c841;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h437d0ae23ca32cbe96af3f24810ecfe016fd1b1bcf46e5244e2d83ca8e9c140854d0103eb001646bcb0e8237bc011bb353a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h223b1e58e6655b5f7b19fc851b694a25961d51963a3e345c96a631475f978fd8895599e4e8ac7bc6df2fb29b021baafe94b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12a3e7e30ebf0bf5652f4c8aea19c09e1fd361d9ed2ce7d9edd1cffdab73fcbf38ae7082bb9bf59b3cabd2ab8d1dbb9cd051;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb4c7f637994c05bd92f122449a0ff699a72f74e54f92a6b8835b9163269ebbbcf7811f62eeac58667a2febc236feafaa63e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf43eebfe07b1f2b3de168517961f40ffedfb221d88cf7b0ccee577ea91bab49f103307669cf78805ab70f6494899a6636a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha61e016c374c1a98d73a752fc901d4344c1c19f1c62a468045645754760c23c40652faca40576f3520d86096b8c1e6f1a578;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h958a3b53ff30196a78c6fa3d580af21ca273f6085f91062a2aada5497523d60d267fa3e3164bda3dfbddac4f238012addb54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7f3c098b5cea1702605bbd21630bbff8c28fdb700e2f35638798e0429578a5f5b90b0b7b13141a1ac9c26a4d0a83749f96c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31f4c21f9bc8ec4e26ba563611b4c5d53af976a48933e59494f01a78c5fd9d611eec26700b1ac5d2e856b1fb2a5147698a8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fc8caade9a028fa26c17b7749443be4e6d7c6775dbb9b2ce218f992ae76e43fa43cd120601162ed7a8d15edff7b193092bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c2b0c2b54da8efb4f2cc0a2e574a1c09560b3718a542700d46e6feaea05931f43c3dc91e93b89f8023d3082e50db6efcd20;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb18fe6971a087c75553cc2038554ff9c8204b9c624a041b204361bf805d56d7f1519bf36e67ac53e23f83b6b3b7a87f2826;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce49bb4f88c9dfc32e8f3649709c1e0f7a8c5c9bce069f3c05ba5485dca00254332ae5193facec420168e95e819990907e6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba9f1fb4550173d3fa96e7f52ebc5350120615680a8a54fd66af85b7a68fa44e5be2494c9f0334cf2f5f170ef19f54c04530;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9a48e16a4b6804270c449f924c7ef215cb3f2fbf67c85464744d94087eebf5ea2c0024aa8bb578b1f7a0328deb5ce18806;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4071f4fbc48a32339b2e5b1d896357070345e424a08e6157e1279bdb93e4f67f2ce8a6449d032abe19e624c9a0e7809ec4e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha72ffea8f893b0e50263c568b466a6e2b2cd76fea07a8b6de0cbcaa0d7dcf1acc9b5c89926b7f72238414791ff875014033a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h312d909d87c3f3c94f79c5ea26e72216000330a07282819771ea0902c6cd254bcdcd0451a7077e5fb3056dbd413e59696913;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacec57b0036477c2bcdd82e1a78b1719e9c9d3f5d901932de7064b521bd4d144c0cb5557496c7ce9d39b694e12b59d30e6be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb27ec0d62296012ab40d563e9a656c479617897519d9a02c4646834e5f3a8ce1aa6053b3e0c42d59a8d0e33734a0c7d4f282;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a472a9952e620e6ee77941307670805bf1138d58d35d44933a77c7266800585dd46bab8c2664ce9481e3759bf61529fe443;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3874b1a954f75f2e046d71ed0b3c5ac6fd93511a4c5cbd03e5e254682a6b92d9619b8ea36412f6a2258dd95b9858ebf3906e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a2d9f678901fb6cd5eba688299b846871c8ea469ebd590286bc06d6cb584f3a921239110e79226a2e485d56993175704b04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6db18d7d7d0f0d85fdc8fa2c71ca7e6d1959fe668c9678038b2885713ee9ece4cd0269f88d59d68f738f5c27788e1d4e23d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ca349247fa51aa300b720dc3e1a4133a76671937f3fdb32c29a0db5e7871daa6aaaea03bfb11835c13b6941d1232cefbda6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80781bc32873ac4e664fde8aebc15ec58da36c72c284627a07f13ef6d2415cf4e2ae6ba60a38f09dd5d092b9990bfd8bd438;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8838b13c1c7ad2edb8f06c191dc90caa7de0fe23ccbc6e92be60fabb711c08e98a8bba5f7b347f3e82ab4411f4348a804074;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h499ab3baf7582602929532940690e70fce4393ee20b9122d63ca568a5b9304432d39c7b2e9e7e0ec63e967257ee182b437b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb13166dc54d8c17ee63e3c449a97c0d7e45d02f9ee61ee534190ef07c772228eeb2a663f6ae5933478e96e9bf38128fc85fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd234d7a8982a5ea0ad7c948f5bb75c3841393fa90d73217357f70069795499a951b6a7650812efb698e3f9675de6ebb33b12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d8bc9036f008427dfca1a84a2ee2443e8e1b1144775a3dad6074380a93037697d9ede54f101b20da07f93f2167aa52c0313;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfbf7c76c98c5425f443db2e37e5e7badadee01da7867a6a0f8c9371342a8fcd62c23ffecd22c35232748b16bbc4f5f914a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9519594cdf6b9f062b58ab83216211f2186b4fdfe0041890efef5cf030994d8427750dcfb28c7ae6c2db9a7aa46e53d6b1ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7609a2d5e007f9f310aec1bc73b579bb13315e1bd17a5dc4fb6f600e69101f34180033d0dd2397a662dec0544f711c80e68;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f6afc8dc5c0e05c86d40126c41bda3146b5c0ef4ace384881bf5e940a2faa94a0eea40cc6d82569f27054b98271f1228146;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h429b58ec007a61518e49a85dd0bce562f3229eede939e101c69c57a744c46620d285c93b2b0864f510e424fbd25c70a483ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h565ba14ec7d68f0ac12ba9620be7ead30520871fcde8c46f6e915086b2902c46d45e7c24ef6386f5bde1f6dffd4759e08f68;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94797d09e953ce08f124279a91aaf77c7e9ab3141d0d4b24c37d858b7a3758463f9ccc9a100937d252c5e3bef5604ae54987;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b2b5198e6840329d28523d3dc1cba1e9149ca476aefc95ae5bafa636095bb80ba0e1a9d35dec1feac8e3974ba2fb6fb4224;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6828e0200b792e347b9fdd5e29760cc8ecea200ec82180b9d0b305a071a729e8df23005864f3b346668b100036bdb0459915;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab6b9bece7133b39251d251b054b80dd2a32a0b716dbf00318b9c376cb516b54b1e0c50d0a91da06d4d9c4e6dd64eca4e09f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haceac1e48adbacf7a4d4b657d5d4fcb743c889d3972f5f1fc03d0abd917e37cf63fd52a1f117a72a31a35af13d1c4c289cd5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfeacc42748a2fa215b5141f370ddcb971796364d61e81a2b1230ad00d57a23e861f72d37d62159dadd446518f53aeab6436;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31cf2b3c1302cb614ae99a4b8ab314b45b7100e981769b5439ae5b3337b12c479d31af509e7856b91b90635fa0692fa72f27;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99da32d0cb381d8a8cc4b81cd385a7a0e20c916b08c11c5e5ef1505fd43c4447cf47ff5a546390132f4997f2da23dadfdfc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h951fbeb494a60abb26068b7d04b0880ca39b61ed08dbc3f4602616ee9b4b4a4db7d928e32a6ea4bbbb15185565dec06296e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba19cc8f7f1c259757d01029f1ecdd6137ec5cbe16ecc36b6bbc12a6c183ae49a4a738d6a3a994008d80469af6e160c1ee51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86ac584fec2c446d5bf2972df73975e53c9172ec6dfdb6496c708d70b5683284c4e0006d014cccaa51562d383ba864c5aa8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8056d50ed23d8c074b05e0777659c3e05cda3a7867faf52f0bc47b68c8a4529fb3e1098e2cd5056f94956ea6339eb881fd72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd46d048eec2070e2a2c5dc2297cb492303d07c1d183e97be12ebb32f0f4bd9c983b9db176f78447671145bd0b32cbd743f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb97ffdf14c252b23a27ab21763821ffd8cdb4ba6bda5c07b049a59a9d85b798ed6b87d5a686650b89efe419b1f535beeffc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d684fdb609f4a16139f938584fe9fa96542e30016c845f9ca81680b533c07f55ee943821d4f64c68aa4bbc95078b8028e1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16148bffe3c9cd9903b2cc62a80cd8aa383c8de3b969f106c0b9cec07c95dedc9eb2fb17f2a9fd39cbe0b0b32be7a6d6b57e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc76650f911cba6f616fbddb7dfbfc91986b73d6f538cb7c8c8290d72b77c356154ccb25f2e74f9e25e45365a6f1eefb24f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fd2a9d90c91aa16f8ddb487dda081d152f4160c2d5658752dd674314c999d601d0000318e741e46d3e5975bfe8392491ac0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e3f6e21c21ee7a384b50063cc19e5b6f70255025fff9ef2eb14bc2bc229ac4c1487898f1fe1517cf7058510dbf792ebbf90;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdd46fee8bd591155c2ff31c777ed21a4c4f4966cbc99e19a6244ad1113d23687e297911c29edc9d217d4c0b28e58cc7fb31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cf1398eecab62a34760912b66e6fac1e03a6bf51721f8e245875c10a8a6ebb91d5a5de2b8e978a2e3db5f34ddbebe521f1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d88417f379a516a0c492dfde1678879a4feed730f6f4f21e239ed144f418006ed233ec8edde4f0e27ba4f19817ec83dcb5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb290d767d2b30baaa79373ad3255a1553f869fb7e16b0a73079815c76a78af568f7c36ff16f4cb246da106e519326fed248;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4164a1acfbed1c2cbfc7e738d87c7d8bb4abfbe231ecd173d37f3170a4e21d29136f39ff07b9e5efb0b4ebef799a8810336;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae183db172accf11dd8ca059de143bf663d67c355b644f37f9a50b0288b025d1252c839752b75c09727671b653154b6be271;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefbe4098bc935c87aab2e8cc839dc7dbbcdcda327abbb8bc39d8c09299ada205c539c9628ef625405d5f1846b75a55c1ecca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h122a4176c70ee4652ae3980701c967c217ab7cf433320df3be724dc22f1ab598cdb147aae86e48bd3b39c7b90b09e7c49801;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56c2afcb1e11f72baf9623e0cb90e305ad3908bb0adace8451c5e9a3904f3f655443ac5fa7e05d74c1a1ae102c28f8e2e1dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d93522746d73ace7f4d458f8e32e0937cc9cb2c64570b33505e17a8ea745e50ec0d055635def7600e00e81fe53507aca3ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65913ec992150b42b0675418de6f3446f27c7a812a92d3834e5db658c7f01794b50d477b4873476a7081eb15c25c7131d117;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h353b8ca8d2f1a6c0e3f24026e5dbaa689166b61c718da14b2fc8b267e281f44060a6f5cefddddddce0032e29039e975a9545;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab928b9590b0f994cd56ae7cf96b1439f8e4457fd795418e33ab5a3e0d13ca29261deeefe84de416eaaf9c0c5918dd077d55;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f01d8efed8843d0358622fc8b7dc8eed18963e7ce78fe099d87a8b1c867832178333fc98d33330e3fe0f280b08f7648ee2d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc535c3a1f42ddb39183aacb3fc523ee8f75f73ca64e826663b555879cc23701d2628b3ded52d1bcffe7e3ca09d2b0e7133d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd30ff0496bec3a23032347bc7d95220dd1ce4752c77e97152448ac9598b78e52b60b9ecc2bd3d3eebe71a94910b497d84e9d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb9e95b4d1a763b21b6244b1c8a32ce17bcc518b63719edb80b0838683246fc4b080c05b2e34f348ab8c38b6e5d4d6ede487;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ddf00064ffa7175c604858feaaa1d448abc4b20811c4cd8365af63f56c0b28766faec3ba69023f1d9c8da4965583703508;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h270239eeee5893e553414dadbe9e430a3d1cd2c0814e8e205534f662f55fda73b52a8fc0bf0248443d745e21f439a57a99c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb98b4767740b2c33ac104c4cea6f9a7d2dbb5edc0a06fa5ced8b4cc8092959cfea1dabfcdf5842cf12d4e7875273c77acc54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h872a0cfd37caae006e085cb5d9e08d674793824508eaa2c0950db611704c73522657a94e45f5ec806c23db22fc5c754eab83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26d42cbe8bb22b0ebd8436d216b8bc44387a03287444669c7e56b3bcc043a3ada23a398ec76243a10783ab562c917b58bb4c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19b7bc265a99009d852a88bd6e86902016c0a3949ae66e2de076bd237e3c60a2ffcde435f6f58b493b4e219732149cf6bb30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44c80a42a567b1b45078233719c9bbfd90375dde4c60e3fce30f1e7e33c6f33d06423caf7de531cb6cf9cb45061e24e34919;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2768c595c6581d6d4fe8de44077269b66f8267e7b26375b0889b1c1af6fec96703227ece8f984cf2edce304ce0d5a110298;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb02794ad4a3ecbf3bcce6cda143374750d3d3e914b3ca10563419e16fd9fb17f5e2ed5caa6e9e9bfe2916b983b1eb767bd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h750ae0b8e6f0e0eafcc19cf4aeac887cb6e179fea57b6b1b5367c25121826dab4adfe963f144ba003783f433ac0ff52bbdc0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2762490fbfc3d16061ce2883ca684bae8f6e54a76de76353056c05132090dfaf344fdb7658c619cadb376c7788a731b97dec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6189041e37267c1b19a1fb97d4d2c71be8bc0c63cc2b4aaf7cd4359aead13c5499fc3f3af5994411c3df96b8ae719ece92f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb08971e05a8fca712dccc9f9dc7359481133a4459eb3f09f699c211c39c0f74931eab0f6e70026738c5faa385d362870880;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9982e1abd4ca352e313be231f39d3826300ccd75bfae557b1caedd8645c3e9d98fce228a4d3b91ebfab22579da7aa7b804a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62b43ba80473b33fbcf288c263cf01d750c06d5d8f47adb5fcf52e79ccc73b7e2a2ec98e10ef77ce5c9a4beb1ffa05164993;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h444846b994dc91aa295ee40342a9de65bdddfdef7645060c1cbd3ce6c1146a83c390ac5b6590b82350582d4c6951b6352870;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19f25d24e3b14306b27c7045e97ae3e4d4ddf3c4b2122d4d449879f3be8e3c474b0d1da2ccc1217a126d44675ed7b33170e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf126762d411be2f1cadbccbf24fe9295193b56b0d4e589c0c910692efb406daccdb0bb92cd12123cd7d063b13a34a78768;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19c41175f26be1aa4a13079a2bf6d21d4739c47fb838540f8ad5c68c7298d66b2cc5c7985fe43b5b190f15eefeb9eed26a94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h568759ba7da678c6f358115c96127fa59fd2300bbc496d8d115b6b2eb70775fc48b331438dfe3abe07ffd93a0183bd40c5b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h817de72e2af23588f8528eb13a78f41723e3f438c182816374947f4918dd432d1735ddf0b0b1576b90aabcbf37b5bd2b8750;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b3a21d43ff9ec2998fc8646e1d30f1fdcf70dc86cff303686cb4ca23b1aef31c31f80bcd72ded581fcbb5b27ab9722339cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1585c22ee4b9152ff126b091bcf867a568edeb114f1be55a34ff50a800a99833bf27cb39a1c9df6f949e35742a695977f93b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c25883956343a9d0fb5934310538c987593e615053e8153b2f4b370c963ff314704b09f607a8030b13044a640fe209cddb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h951ca64121fd894515062c53c3782de9487471d4657a108222e9e067208e7d201e0a95cead7cab5144437ae0ce1b619937fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he90b0a02772e8f7f2ae84d8f67fa238e1d524bac03af21f00c6e8b394f7816a576c2a6e64053a072f19b4ca99dc5f91928d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96941e0405b7eb42380ed328e5f62dbed8aad3454a21650c729d81462fa09581acc9aea3a5eef54a1e8e73ae3cabe97a4d03;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb917c2c1934f460ee4766a6b02964511fe8b382a262c1a272e02a92b5dbfee86dc3a12e1a790183cf383991a3ed89633450;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a6f74ef39f502755610290a2ca5b0686ad9164cda44a2f902462fe48e6e31a4d43f1797ee15c748bc6fe840fc11a3428b47;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc61862556b92bac4a7070ed50e2fa686944529d245c9b349645d8a19151180b089d7ea2a14aca19b47da85bdd2a1a238988;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1142ba6c484ca01e56c1324713ed1284a4e005cef7e807c7098ff8f81b5f2a709dc4b3ae4dd113c6b2682aa4f2dc00bd83e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h861bf97c2d84fa3f0488d3f91fbb69330dda8d7a4199cd1dbddf67272bea4368131fd5a5b0b391e88a397977802f7627b181;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb6da0cf898cb169e378915fe3bf08e9b0eb102b3f9342c54d022f52df05dd133c4151eeb09134f5de48677254752115397;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8c5885e213b8b8f1727032cfc7141f9cbed52d7a180c95bd3515b324ba4e316fe1dc22e381c03284bbace3bd582c6afe81c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a0b698282c6e3fe2e4f111d84afba09df66c4442a840c19cc28363b451774511c1c3d51eef86f864303c3851f66bdd5a20e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd8bab3520432a7aef43b78da1f49160753463955367fa9e5e46228b89d8b6a7436aee71f302efb156152cb0f4713187ad6c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf229c4fd42a0c432c29580065d0a85d4dd9d93dafc66a03143ca5dcc2406f0a937b5720fda2d58fa3582bb005d4e762d03f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1351fb7bf6234263cb93c7438529fb73e5d6ee3cdb4d7cb0ad4be26a4f78feb5e3bbfd3159808c83e8f364148ec4b7de07ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h937330eb8adc834045dd1d074c225080d1917e458c4ad2a7bd26fa3806dec417fc4cecdaa76e0b9acb53fba2369ed614b60f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54a27e3afe1d263765ecf982a073e6d2f7f451187d940fe52fa4667984c7c94261923513c8af4e9726a4a4af6da8566f6db1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9abf7511f3a436d023bba088c98affe2af3a6a61db6c1991c8188d10246ea5e865e7b26d4c90d40841aef0e951b5d5b349c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ccd63854f0b47e5ee3de2f78e447c5f1085dfe0a12f1f8555e3a9c461c8af68c051af4ff46c420f8f40c942c45dd3783466;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96c4556aba19ee0c028eaf9772770b2c80be6cb2cf084af4aa0efccb9b24b2d24669d65fa0a2cfc7952eca1154d74de45649;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddafac17f8ec23a53c2c874eb48db3640cefa4764a35cbc00d02555c38f3b140144b16b6506f0391bf02eb0ee77965a9dfee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdad7af0fa5caead3099ea17385d198f1da2ffec5047d7a8f3a25e401a9039e17b69c611f6a80b32cef28677349863cfc64ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bf1cfabff5efc1e67c666fe9446db12afad300a62d7ea9427bb52753b2921ee7586daf131a8e948efb97a20f4989e467460;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32551ca3a171785b3c745a0e43e1c637f7d2c6520e3d0fae3e6b0971b44725e3424e8f197b2be0294868d19633938c29ce7b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cd004dbf8156dc080213ed7129d72dc7866ed5f1cf53252f1e8f6f7a4e95cdac9fe289e9e9b707d4e6b5907bcd75df506ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7afe7cbd22592176566d9f459bd041c8c17f651d42bc348d847a9f03fbbf8b29ea82a9334afe72db541c4042d6e4cd5656d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfa91e3e5c5d681cfe13f1a0c41f5e1d943073cd0e277877428a71bf7b997560fac32f7c783c86faf3535db6bcadd19adc06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd49ed20de332220adc5c2f2ff4e97e7e2c1d15734b9a13c72e58fbc7aa349fa7074defaeffd092555668cc390536f8b8e17f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h296f71847bb425af20e04c7c26fe8891f1591a9a0cd4a181403993f2cc3d748d68ec265f7126e3be1df3d518e7ea70ada8d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58863f0323c2eba77aef4c3947eacca1621acfa766c410a02eb5bdb014c51637bfa6e4620ca419a79b90f9c294de2f4f6221;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e1e4c6ce38a300e9d48050a8818840eb31cb104f46cc5f7138c2d882926543b609bf595d7dd7facbc8bf8bf575881bdf575;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79d8c3e6a11222096949ada375b0f114abb4ee423c53cdea806166bf4e3b1f4a7ad3903eb1e084daf15c8a87ab4a9cbab04a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5301ccb1dec671272333d06b300f08bf2ca802582fb825e49fefbdf22a6c71914a0257b8d5ba5124e532a203e4f0b33a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f2fad75d133598628516fac76064c22e0151049019d4ed69691a29c6bf94e6c7e7408078f73c6902fc7cf0edbc2330281e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h168b4db518f922ae9acb20f406fdd4b4187fb15b02798fee443a4462fb457cd05f625d39df7bdec6c1ecee871a545046b0fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2e8c9e7925367cb981b6d6f298fa8f7aa57778bca3eb3edcc7ae54d16a9c45841666e970efbf85a0893f9093e6555ae1cd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f34d813261d412bcade8acae5b1071eec90f537d1dcfd1260cfdca65721606a632498e093d99cdf1865090c1ae58165fb10;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae9cff415a2eafb1dd44fe0f5574aa59273cff8e5a1b1ad7149e07a334c692ac11cdba4b42969bac88bd8d24c544d701a91d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4632dc3fe01b327e8453e1c924a04a301e589eae2f4f3f537ae0f102a3b2a23555f9ce0c1fba925b2cc21ba3a474606c7785;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb922a21a7f21175dcd62c50366d927ea470d375728cdeb8abb5b393720f07e45b9d7cd87767c2629e7a9af595d75a588f3a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6054460483e03a7a8fafc7a301a935f3f13226bafd71fdcc37d59a2c407bf47859eec3022fefc68a3ed17381f47dbecb1905;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadb91a37b5c798fd1d637c85184e1cc85bc4dcc1dd6f89ac852d189b932ab434e13b05645c6858eaabe39a04f952f4391ec9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80908af5db502b012288cdf1608d09cda9d7d6a78f8c92e8e01aeddfb02632b2a865467065df52d711f2ba5c37dbb7607466;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98c4728153a97d11616d5a9edc98588438dfc90b3d176cc1eb156c46dd87cd36e80cdceec637e9d3e08ad60a52e7b204b3b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h332d84ebf2e7b47451262d0229566bad37ca489f259ad0306a3e4fe6a4d8a1092b6fd98d910ee6e79fa0925e73bed5005080;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e3b34c28c5d91fac250da03e453b39b5cf2d759319e8afcdff1492e40c55f4b091d6a72efa61ee06da11d29609ce71487e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he964170c70c636214d5ff735a6396f096fb8a82f0ac17400b1e7b33da4cd28037f8a5edb12a7e5790dd88ffb4a25ab7a4f89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ccc918e49ed66620314be0d64e1b1b1159540d278dc5fba4d542ec027c30956a9eaeab774a25ce54d36c76bb4b0aeb35c9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18a6c6af391a514f5b02987e56de408c6a46dcca9608ebe702f31c04fd6bf2782bfa4545331cbbac4ed689a05b0fb0df9d69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c8c9a546a376d55fc0b3cc6a68dccc01b873d948aa7fad71f2e1c8f207d1fe34946fa063c60db8c9826018c6dc4a8f2d213;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habcfccc03919d5c5a02e6857302eb755d1f7c6476259c2e2af159ce680d663a991b94501723599f2a24513805dd1f8fbef01;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b257da861a0027be3775aa036fa2e0f3ae653a82f773e39c3c06838f28320e33f8881526ff6f5260f7bea33f360ad5fd1d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9789c1823044daf8eddc023b8b3181763421ff9df4e7d70b50ca4209e78d4200e70645fc552c965dedf2ec45e1c239bf2356;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h938736f9ce6667c9349c25c0bd0fd4c6a2d00d559d87a18620c64eacdab26eea3093272e9cc5150f7f6441d669059a11bcce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had8a2db9f3b5c9d572903987088f704dfc31865292a47ccd6c6ca38a60e3e0f41adfa35fdb76985f94f2afd3598b2af09cc7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8bc1ae8e3d3a9af40ea538627a6a4a21862054a0f6e8cf5bcf24f50f0a983500262cdb13121f70f1bdfe16af03857619f44;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haefee4bc0096685e2c582cadd98ca943a3344546f59f98de01d2236b37cd38d0282f9f0a255d342bd61a98f874d9792ee6a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcc9e9bcc93dc079629965ad25464d776aacd947bea4ee721ddaf5cf60463a168c6d14ea80465418a361485153fa601fdc94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h445764d426d9849326c7dafc944580d1eaa2f8788c911fb0c0579bb959901b377dfb9ae07272efe0cd1b928ab1890f014401;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7be465aba38a5064f109416ed2275035613bfcb3019deba1b261a472076ba30e46d6bac9a8cec1cfd492c172fbf82724ec4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h895f6a46b0d8cb0e9cb7a0f97beffd5373b87307e6069213b7350283d32f58a68bbf5be5b94a65cda0e86f422fdb1e246b09;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a3ce2b2434166764607f1a702cb213bbb0ca14122d1cbf9c764fe8f3caa2d2a18038fdd64604cd4b34bbf520150cfc7e807;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26f642fc60d3a3e967b077f8fb3593b38eecad6019e8dcdd6605ec4adb8b1767e940cfff138167f5fa5adc8625086464d76;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69028f549a7415abe1fe6ae480c6872bc6f323d787b8078a6c3c6cb549dcaa5a0f1445d417cca5c9f79fe3127524ed9e7632;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ad47441d597c44eb1cf9196e397e648eed0496ae170f643482fe26e908d8ed976dbb9f9dd631ed6919b795ec65b37fb5f5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb69c12f87ab7a4d3526c628445d1f12a102db73bb10d42be5afab9167103e20fb7e23926d279387315883ce96ed3ef41662;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27d6c9a0b61c295e519b2d3d851aae5b3fa6ca5bd6898ed5c88f1c7a346aae3ea9399eb420e49bd141ed9d5deaef5949497;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0ecf8d242ea8ead62843d0e5b2d5a82235973772d6b32058b63606a92341b777666d44f251af4258d74ceaf26ec0b33d69b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d9f354ee1cfaa95447d442dbdb473c2a797f415f618d6fa3449d969fbdf1f0807ca32ab84341177328716f4c07eccde0d30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc119947e32142ccf331370f8e2e0c396a98f3d2052d8b9ccb6a1e6aed58e9c9b779939450b821c451f7734ae5541071c359e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf53e777405f8dd8efe742ed31f137009b7c51aa3c7667d1c706c38cca5ff820a7073949e1814a8c4402d3eacca11c1370866;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb800b607b3257180887158090ca9a7709bfcabc99d0948b7240dd9c4d6b6aa3832375595c508043619dc15487c44d970f463;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54b0e1ef7340cb822e943a4fa7f4841402416042e8fa67ad13d3a532fc8cfac63c391d78010d232d65f326dae3131eb027a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h786b554581e4b45a240621868152caa549b5507e579a1f3da144e63991699f0ac2d7438a5f63429b497631018443ace87770;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8e8ca30f384fa0646f9afce1d57eea8e1270b7d7f14e80cf6988a342242b16bc336af3afeb25388bfad75d22d803ad90c3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69104ec9cd6c69fd1855b6ec27a94315ae93a93fe7b63faf8477a07721b5fd7c0b3a9b0880b0971d650107a0fd29414ce281;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13bb7079facfa7e0ad6e518ebbb9238b5e3fa12e9542f42246c110a9396267329db692558e572e62baf73bb659f31707d9f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h807dd17035d69fb3b19cb68d2ac1981ef854bd9fd3140bf9940362b36971815694a84468b14176cf437332a95bd2d9671f49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7dd1afa08aa5258d9419275d6b022aadf1b36f98f74f9a8a46047785202464c01e2c07efadb5709bc997a25e46466ee0d307;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec5c587a4641faa0958b7e0f7cec394e52b921a804b6123e37f0ac26b013c618e7ee271483ef9478c8cbebbf30c7fa8732ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e43cb358720c7a28fe66c0057f16a9670ee0dadbfe28075c373f49967c2b68c75a61d19f06c9b42cee73a0c9fd21354a0ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c248258905c6576f2af7686f1510e8f94ee5513aa68fc410eb3865c586b191f7bd5bba736ad668a61c37581356df5a0983;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he19c0a5e700ff5a62be06bd0531955808787ee765ab3f81737eb32a8744e130d7c46bca9fae22b4f4c1a0eb82096ab0a61b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha96832dd801696922dd8398a687857a0c5fa974387508a9208b39f043b24409967643fdc080276424d2c3d31d7f34d4bd811;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb54e458774b2e42bc613b64b6de6a3eb8d133cf706ffac25cc4e1f079d34b5ccbab32beb72a0cfca2a0eb71cca84364cfde2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cf505a8217551dbbcdfe195a73ea1248c6b71f88812773d6dbbe11ba509eecfec28070ad587e489c5713c4a6225d03490b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f0ae1cdfa74e1ca7d541b4683a9c64129f963c4697b67d10da86bf37938c30d3c7b16cb0e4ffe8f634215656b757d0de335;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d49b65682a2581e7042baab3bf340a7d51db5226d5ffb400b2141656fec4d301a06fd01897162e9e17673057fd4c3e1e694;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b0886badbcb8de283eb9e3a33708c7c6eaf0277a14d86e96ebab2ab0a4a85f23c9cbb3e7cac679e8dd52077c3cb7a13ce1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13f3cd3053294aa41ed050317785cd3f895962e36d390e11c15d23c32c58314b22667982329eeb39b2541c1f0c457f7242de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha58e71d709079eed2f51e586f0b2afe590be8335b6444925dcc751f194f5fd919385b74779233425c0ab294e70775d3ae38c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8812b2dfb34430b74663101671ecf235c36e021339971252dd924d3b0e908d1472d5e8321950b3d1288f7b5c4bcd90fed526;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa807e2eef5dfe6cf8736b4aae18c03776b82d5025c5c65fcd83a0281b41f202bb7bcf1185685898953d30aaac985359d361;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b42aee9b6550757a0f7500b18dd65e08a009985fcfc6f81ddf3f553f654731c9340634ee0d8fafda30579e09338fb4d1853;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7f5117c51f7d11ce659db4b21313ed960e08b800a70ab4b23ff2c5ed029f9ff41d0f96ad8545d16c2423a8f13afde01f0e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e692e8f0cb2f99b014a991189c7507819a87971cb1cdc63614b4882c2b7fa625b1d2d4e4e71d6cc51048e069405af79bd3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd3223641ad88a06de20a16ac6b145ed0e87bc847e24b0824ac34e5b3371ea2f37ceaf686e2de15826ad8f52f29c4bfc3c98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha20ccf96d52973d77efa35ec2f5af2455afbc1bb9207785f82b37595c62317210925bb80c6a53b05dfd44f05db40c2788a77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31f3d17c8c6fa577f6276c0c885aded4b84038876fc6951033cc2e4aa544990f525a64fa58e9e4820d9a47d67799414165b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he507e68abd798348379ae1004d25023f1bb1df14c6352cd740f6d963245bd7426af6dff20d50b99c376eacc9315276c94422;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf7bc21ad11ce2bd5d367f0b31d38d1459f679e8f0db9d539d03cf2d90c53a1b9078d6c53bb9be7e91d2f4a19af4ceb5a7f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3575ab0cc23098b1f4a0a4deae61056bfa07edcf635d6fc1bb83d300ca403730c48797cbc16864aae2593a470c8ed705a039;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h194db51167ac3edce075e23317bfccfb75b56b01cc69b16cc82288c039059c433fd5cd8329ea207e8332eb01e3a87687725e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce10c1bafe21bd558cf7427d3797296e9e10a08e8af58f05fc5d029a94319d9fa063f8a50ccc0017cb7d7d312aac5814efb0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha90bccab89e9dc22cf11721e55b836be813eb8baee239295ca7867e136d21a9bf4bbe2ddd5f4faeb58fc724be3e10a4f25b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45600c95d9d6f3020ae560fd49dbd744e1dca4aefc3b7a8132f06d2a709d783ec140e8dae46bd80bafd0a8c6bc0166459fc5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3832a8a61630ab43d24495fd476cb6916d8bece7895c302fd48d965d5b3823275d1d8f80f70aad26c8cd01d522a683ab4ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h600be2d4a109e0a915fc142ee6437cd8c6626e955e735b959e7aab33b61f70a57b184d871e097d496707282753ed2d714302;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc048ef3416b62ee89ce7cc8113a3e20b912e85ebfae3134239809cb576302c32304ed324e60d30b5ac4141f6947f4969a28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h922d5816b511d58fc8a8d606ef84dcb07e8a3cf261fcfb81f6c70a886ece340f8e359c3b06f18b6dee3c7f4fe9838178f54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d558b2d6de046d4821e97046fc8d116f1256cba54e02162bc88567a766a741b0eb229ad718b26f417e920eb1356be79aed3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf095b32a4469f37df827f9300c244972cb455df03ffec0370760fc132420c0c318ca1151a0ac82353df6651d89c766fbc2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf598cda044468b128d9b38025688ea5907ca53fd99a242797a498213a860db3f0a1a4910308a4c56160c9686e945589eb572;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h553c8d99b9b19f152925eb634f39d3b4ee24aa1b3776523886571d5785152a0e6afba983e8c0ec603fae372fd144282b8648;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61839d9cc692ebd031bc1134d2d9050aba6f6a21d0090643db5a6a5b4e5ba8ca7648248dd64278f3b1ea765241a15a133100;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf3cd4845bdaa6ef873e9eb715d4be6643ba3259e5547124c7b9503a8a2a94f2801c133bc66c9b5544cf7e4b87a6961a9cfc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb82f5a17afdecf9d20c1a0c22f8e1bb0af6d6d3505327f09d58b81115d27c8d3ccb6783ae2cfc10f7b3d9120fdd70c7598f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9626facb85930545838840f10683ce41ec38e8a13e5120d66f5d9dc2060441c3b1eab9023cb6de397d785c8c0e1fd66838b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20b4ccb6870bf76a8d571625114bbfb8235cb3c032c89c41785428a3f74eb49e4c5afca1251bad2a6ae8f5114042e74575fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d8e4053b475a10d70d25af5ab56e8c3881b265268eba591bb3d17929c6e0520dfb3a62ba7c238ce27248d8f65fd9448093b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha743500290ed0dc3e2e70f1756ad8dd7aacfb81f62f6eb439e049f58884618b06b6bfb3fb64f5d4a02fe63f61144ca2f3bc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haff89f7c8dc3d8337284952cd2dcabe9334e6176bad1137fac3a74396bf52c6b055a4e2b2efd85f93738c645e1cd1e366867;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h281f237ea9cbc47b2882a0cc6e3b93f63a19bdee134e8abb7daef5999acd1036eea637864d0051ded7f233a1be9ced606236;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd0e0f0b389ca6009c7d487cb53dd989670e8ac66914626f41aa5bc121888ce870e8727f8cf930af9fabd8835e44d7d33971;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1cb5d14661b5a9626c594ce54ae4ec5ffa2f442fb2513916195cd4b7618749bbdafff2829892b09719de63c07ec9f279474;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f72e414df14fba0bdc7d108d56df694b4a7b9d819779ed659a80ec7037ad9dd11461a72d621b543d2d6677846afc154594d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf227f092b596b2dc7190f2e6472ba85f91ef4d1262f6e2814cb031ab3da3705f1312e3e9e7c98b223f49e39be50e92639a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15319f4d3be7bc1d9a889ebdb185d5625fcc57f9bf7102bd1384c0ba40e060b055a38fa67b594121d14d77d486da4517f475;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e5f67f0c4f4c9ac65e24d95c5282883e6cf39afb8cf7b94480a96d86ecead2ec09042fb2f9b14f4f1d2899d1bb4562beeee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f32da1524b0f47f056470051da6748e0f35a39b95d9d31d5adfe29a21c3305b8ee9c2ae67a169d6c1f1caa173e8a300abca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56d047f1bc012a718b159d0e17fa1a56b05e79debd6679d23c3e5bb655689f4614398f78bb20c15977eea58f9bfb2a220505;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50c2a5771c060f619c251cb7332ae4a5c6e1345d2553eb830dd00b1d237cd20e57f894c1b7776dbbf836dd0d9934f389e999;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h721e1d005f31ca71bbbc895ba04045cfd48ad528d811200a745a5c3cbf2694703ab5c98db32778d718ffe8b9261560ff8b80;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0e547f046340458044411e10f10290a652050e81dbdea5a841acd5bad5e3c1289fbad525b75db8624fcd1d4a8282a55cf58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h590949f9b36ef07ccf1fc97a66e9a7747fa34425b950d69e1cdeb2b028e4da6fad227ad5ff3d6250b4a0e64c0a6344b23254;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2e2b0b36ceea63705f2b40531c90f6dbac5e2bf7aea4280187bd70ccbc85724d1a4e274f6c727c7b0ef3041a0fcad170fca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h426360ab1af78178de2c97abec42254d4efab336e4c5777ef24837d728dd7959c2bcd4218fa4329088c92cf161923573bc04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba2ed7aed7e2a2bff024fcc0678e9903fe6568535645165afb3d4bf1e941b28c678870ea9a96ac4bc120bf0464b9a23f99bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h770b5c208969b88d3b0c1f0feee4a3a4ac33a2fbdaf546d2bbf89ad1fdc0edb5afb22a395ff9d7165fbd7852906aebc97ba1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea227c0107e98a7680aa84e7627b6e18ccfa33366f0947bad7ccfe901a3658835d41dac369ef87b51e61504161cc5b563950;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32d412f39f7cc81bd060349f5a48b05ca445631c0b1aa4d3c10b0ce304c65421aa8820dac0c6df407b96008a96a9f1ed2c57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ae779f5a33230fc6c4487db35476ba432f9e92da20a21cc04e23ea2d0ef85284105662ab9464903b23e3c64801758d78140;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc07508b6ef3ba4d8559bac4e717b46eb10e83787f1dc006b3ad368a0538b421cf3f8d528fe41d6b47e5b65f715dac63e48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hccca2efa600e1c9ba2962a89e4ed9bbd2ecb8d27ded612c3c12bdd00a7006d8c9471bd64fe7f8117dfa599916986511758c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h348a035c7b2944c40fcb1d8616f5e97b185695ad39d0231950443a7f7f263c73d0ab226cc675248bce542fe8c2bb7ff4432a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ed380a5483868533c101829809622064a74289746dd1cbbf840a262d8c3d349116324b5275b5af031bc42869f678672ce65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37abb257c6c7bfadefa7ca16e7b15ef56bbf52371162bd7d061f4b28945fa6d8ca437b914f2d4485e126221e7214a65a1f81;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27ed2462a1df1707f2c7807a4e7bd3e4185f3b9269fae8f27c1d5496bf47fc8d3bfd66f342548fa0ad44a7c9143ca71936a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5d1703bc47c03903d6580e415d7f43abd5625354e8e51117fa819545f1b079939cf335135258a44e07b081e38ae9eee8192;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5e721f3926ee1c0c6b27df225d9e420e6ea837b09cfac7e806e0164423db8d3a97ad19f14799a4c67c53d2e24bc125fae25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd993d9246561ab930132facb82d605877838f187f3cb5a88490b371ba26799b9fdab934f4833de273235bf86d3921a159183;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3401ba2f25312349e234dd37509a486a9b0f5de0fe87f346470b0ee8a6f94134667d23e43857688e5f0fe845cc6ec4595c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3f0e75c2337154e9a4cf48ae6fc4dbf0f6424ce77137e1bbedc0ded48aa83f1965a17210a66bb393f3bae41887dbdb4b085;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b3ac3910a30f86db29735d5efa220cf53ceab6ccb70bb87c64bfaad0d4fc901aa464103fb9cad0bb4c5f7ea1fc4a4a11197;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7af2b7b690e2c0d7ece738d32bf04cb468dde4b06d7de239bb9d1daf3d32881958052dadd0c5f99a9d7a60a8c0bcb7fc790;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a4e5329ea6bf48c344f33770cca1e9688ff9e8934b36b9ec9a7444856bda808e247781488f7710ed6904064f3634d5e5c4c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac939d78ca6b0c5fae5940cd35f6767cb5de351dd6b7153fa7cacbde1d720f7c7e5c928381dde72d2d32d93e64f1d2762783;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4b7a023993b27b3e2f7508aff2c7797744dae935636c5f8e16b0722cf3d75fdc9674f5956e0f58810bac3837244fbf24beb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h755b4a1421ebcc16cb08429d268ebc8211d86da60a0179c5109a6f34b9f250de95a23b4cc0fd4331418e88f60f4b5a0b74fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h457d7dda4eb9c43974e768d3d1edc7ca9fe141feb6961988d9ecb165e7dab4aa05f206f03e3d27c7d712c56361f14ff8442f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8840967e8d2e8d3f3c18f0dcb8819fc4172086aae4fb520c709f93ef17f82c3c306439f76644327c6fb9854a6d5a98c493c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e27eb8c4b2360d3d9e297a91c5a48559eb35b50169da9297c47b66a348d79fd5a7e7cab5a2b5a1d72c8200c74e715106d64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93ea35d6b112f4fdca36262628800188b96de642ccb0c4dc98d6ed8c1fb02815ceae6d6f281704a96ecc82344cd3bae98494;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ef3630082e2dfa431f9d6d06de3f76ec8c92b6a688dd095bb9e8ab6d2b4f385f4b3aa670806983f0a31c326f3143bb404b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc748cecaed1b1eed3a1b43d61e960400716ff17d29db907c90539bed5a43806a6f5aff2e904f143491340bf3d3b2041d559c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4eb5a414467a34c375626c9b969a65aab751f0942eee0b8e5dcc0e4b65a0a19699b18cbf1861cc227b2d64946c7d9f4adb4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea7c20c772cda88220128cf22a9c2d0d975d9545f6e7f242a6282b54d313f379f2bce5d7a972268682adf2fe058e8da860d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb618dfaf3b79b9b562f59adb6d36a5a0b5e1229b86517f31166c2919aacf18b087fede376e69bc1a7d3b8e319844fe7a0e98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b6844518b234697fcecbfae15077d0af4fdb1a6aa8281681b9770f6b3e1fcf693bc373d3dc959f506921e404c17ed0c7bd6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f777a826cfba3642fc92d57f5d3d9feb8475096f0d90892abb719b07b871318e5d37275ee248ff26cbe4c38417c9f252813;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf3658f27ca567761fc83ad1293c120a204b975852513450b484d214c785099e04696053517f462eb2dc3637cbffa5b46d1ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd758c1de1ed5cade868d1e7a3c551ec489d0faf5a3cc33a61e2a57e3f38204e25024afe29b9f422ca40ddb6c2fb674a5757b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heee0a29787b5100e48741a3c8aee2c3072117f94b43531b64874dc9c0fe4638dc042a35a27446b2bc49fb12fa7fdb587e49e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cf0d90e31780964b6a5809374a6519b0f14c0226afea7afd6e1f0a51528f078de1f0ee25ebf3fa2463476ed2e58b43ee2ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c3cca8dd7a814ed1a68b4b903c103774f8a20e664aab404feaf35c92e08774ce0e68579b2f7652f47055f6b9d1d4435a544;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb7f7c917b2fde046c842b9bd79aaf1990d48a537a0ee334bb43fe9220a2a62e6b90e7e958afd2a058bb714caa890d688add;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hceae3e46624821b33dbf907ce6f40e7b71728fa208a783ae211caca59a8b8c2e09ff155c07594b334cbd85859c0459540bdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd423f74aa4e475b59f63b28dc8d3020a51a2607a55e111b803a3f6ba1d169e942ad3c5d84c3e0b55717623e9dbac10792fdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafaf1a319b8ba0028ef53c60b3d8de47f58746c9121ab4628e6eac3097e569ab8542e5206d88151058f66bf20168c7c35ffa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44c518855550e37b95c910d7fe746b15470af3d9ef84bf524db5e5e3c1d79758c5178176c423333e12a06c5f6749e4352be7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc114e1263ee0c4e6bfba95198c129eb38c357c30114bba03e300928c1dc9fcb16706e804d9b5e7cad98bbe53841f890a1394;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac57e914b5b4f80cbb6ccf2629e43ac1d64fd50849b099588dbe9f3cbcc4323efa87e20ced56ff26eea8f1361a0434d98aab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1e338c3b96325e1ab51c8e92a738a931faa30a3b1aed2802d5f34d7d04f97390541e0d4a22ef6f0e2bf1c14ea5e12b5e9a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f59d64d5cf23a41a78c25828b1d69019a0f2577c6bf1bec30a71e59ce927c514b4dd9eef433235cad092f9c84fcea304289;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h527d967e6acd83f6b670ac117861378564dc8f1772dfe033aa4565a3a09e47fc76188c113d5158ba41dfb0659aa0614825cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h233580837c471235d3db719bcd3bdf867594b34f097378256dbf86529d8e378101f75e5bf9e84a2e0d6d0de2ec061f424a0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67744a7c055492fae8e51422d1fb246aa4c82cbecadeca0cab5251174cc4e28e22ac3303cf94a1666a412cbca9a07e8b4e3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4207fc96a3ae99255650a9a8c91cab8ef82e068b96bc35451b50879671408ad9d1b712ba5b5db90b89b7c293e190328cf6f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a4832e031a7dd01f3fa853d47e17b4841435a21d17bcfe5af20a402dda996585ab7c8d7959ee6e11172589ba2ecaac76a8f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5d5d17019456a78291e5c3808ff0a69302eb48948b1631374ef06de3b06fefbc42e2da4955dbaae7d28d8b2e8cc912e6312;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cfd732f5bbdc778c74e021a4082a3049d9651d900205a2d617c78550fb1b410b645c29fcd3b29d85f9c99f34f8fe8788662;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f01888fd110bb641aeb7a2411eaddc5d52d6287e48b9f7cadf4a461feeb86f7e53aafc599b1bf66567050f234e60405d43a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4934863abdb665406a922b120d2473ae397080443ed9f80ff881b636886dd53b7a62b9d30b37a843b01d8c73cb37dcbce79;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he11221a05df7b453c655decbace8a6ccfc766499f2502dc27519cd2bd178a30b38ecac2fd7a53118d7f4c2faaf328d1a549d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7e0178648287e1d5692541d2d8a013df832f90feb075972fcf72308016e1a34e586a0eeb5208a0f6c7a9514d9794a3fc706;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb60b3c1b05f832abfa62e9489ebfc8c75544cb306ff4333095627903bc691f640d9aafab431b626fbf29d1c42f09fff3f285;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a7f18162e97f6b12258d9d0a610cb00a1b288be3901d213924e07c18cefe9c5774f59e6013d55af00881c7b9ea7f174e49a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c7919a0905c061a1808be70ba05c550ab40c8e92eb5a9a016b730cb6223207605450b4c5ae2b4c8d59da8f98404ad747691;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec0ff528f0a63988ac5deeda2791482378a326426e21ea4bf059fd89b3fe7107c61013ef950552758c9a2e03dd08215c43fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d03b6da48fd7e84939acabe2706a77017c70c728e0f4264126a406c27f8979dd916f4cee53f89d8da60bfafa522ae4dfdda;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d5debf14e468deb3350086f58231982b88b62f2c4b962ba1c6b2fb83a093d2f98de4e7bf72d5142e3a95ff7ecb2b6db662a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he166b073fbde4a8780238067fb65ae98a4c369f94bb485eeb102dc9dee64d60bf31775bf8d32420e25b3347282ef1a59818f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heebb5b5c110099ed172295acecdb864c767b2903ef92069a7afb4cbd149679bb92e8e93d80add822eb2c9f100c5a17818aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7399fe95008cbf2cb09c0c05daad0938c78c50f3db6811eef958efd670aef25956d7fb8ae98dea5cd56a81361b5f86094e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h753e2e21d8f3f47b9017fd45c29336b044b0cc6f77988aeaac53cecda0e893cea385bdad38682acf78a8ef1a2eb8bece7f9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7808cd63e21c558d3011026ea19d75e4919c966a1ae16f66239b2b53c4b4986aaa2625e7fd836c315d92e4ab6ef325c53c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7c82b4b83538cd82851d50c088e37d724a0e1b8e8cf394eda84ba62bf8e5661e377b00fce4f19b3c7020de574f328a884aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d275d83781cf08d07272092ba8f3b233b2150af5eb485d09f8f35e7f5927c016c0d7461e5d27fcb26a30201b59937b25c42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30e5040c515332a170f7401823e31b7b0785a8afcdce19908e072973ff8f8a22f21c0d5401426dfc062820ab1c6676bdcb24;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha18380c8fa41dacc2b00a8e993a8d63ecd451aa7cd3803fc62f1ab7828a3c8968ab3c2b390f5e9aa53629ffe69f934a88856;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94051d7b9a1d8c760a6de8fe36a89ea71a2ce1884694bb82c1f431606579807025fa11437f3c74f43efbdd0efeb3460d22da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88cc416c7fcc0f351b804b6024809e2fa348b5e03c25a79ef32e908be2fd83172cc93b34a01bbe4456d2abf93f31ecb5ffaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8641b59168cf37f5c070c886ea8b31341cbb7acb59eb326f79bb4bd0d5521510293d508d7079d7b1d54d03cf3b6c3b08f8fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40a07481dd74604f53cb8f7f8558f627c513351418c98661c212d73e77d835bc6abd7510e63d99c1e15f8421f4a195ee5ef1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80be90debc994d7044cb552f9bfd4906d7255affa96cafa553b261340032056c60d9b85173c1c49653e6b443d48499e5a32e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80cde57bb20dd167c89073331d6a0a248e3c8c76c7300c92b4c94ff64ee8931ae212733b293147648664c970279eba5f4880;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha31b7dd8869783166de73cc469f17c383e40893e6841b666ea7c758c1a17f0ebcff7997aadebe247d050dbbcc7980a8a3793;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32207b320fd33bd047b32948c99c62672246456b84a4bd3752923f24b56112bdcc358bf9c4111cc55acf81fa797783d30d8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38193e14aaf820e7d8d93b6837da36717c8297b0518bb284c6ad62fc20b06c19e96bd882bfb622f41e7c3bf1c0631725d2a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0a1445a33c30b0b27092a533b075e1c99456e57a294163a098b990f10f22a430cad1c10e3bffbc8a2d5fba698156f6c305c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99f6230d0f077f920aac08a1a84e478826d8c15fe9bd7d13b8a85ca71e8f6eee59cfc64b705a4958740ac86e219ec9f1f5de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21db6e29d149adb545716ab914290046a224b6bef8b4b0502d2c56a7af6778a5e7c6fe7210a030b4577351bce9274f2202f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb8135915a56ed6206df5045ba7b32c54771376940c389c8b4cb40214dbc3e99d28627781c9fba75e2eb43d9857f64c7c113;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20c261a998d42b71999710470c15d80b0b7df53c50de6d3328dde1a346b129143107c789f0b53606af808bea65eb8db580c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6c59d94f2e5178130f40eecab974265815ce988e89a119a9d78bf41efd73f56673f69583479b64771ae1b3fd090539ebedc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae9abb0a68e178a85823e200bfb689b7e5626c7e0924a43c7540d5fbed66a30630d1ec7a208c7e7118946dd2f7a7c9f01124;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfeb65933e036720de55a9a921a01913754d44d3a42d9aec66e90d567f351552ebd50133466231f6dffc84bad5a5b322e2f0c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb797a31d6c730db25cfb3fc567e0a0738cb6c964ad7969b703ebcc2a7dc4ca919fca9aed05db331f24881c8437cc56d646df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15de2c0a02be579c724e15e7ffff05f5696d778f9d3e56bb0b9cc6ba62010cb2f05f207e0b06d44bf15ad10e0812e52108cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39d9d1669178e64bf59ac3c118b0c5bde176c80f1d9269240542c52253a5fbc987ac841d81b7c17046a1af9fdec0fb257da7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd43fc5ff6bfa0f38b1751c545e9ae54b35bffc531f7c80878a573eff8290d2ee1cd3cc8377f3f466d0a8f36804c9519ffc37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedbb989171ab55d7355c778112e026bb0878e7669b13dbfc5f0d5fbb28ce4829b86605bb4d446022487e07f7a29bb9fcfc1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5ecf55a6ae9d8757ca323858dba80f08400957508372bb374caff263d9734e077ee09e2fb3692f3612066a25e8445e6d9a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd23f0c90ef6cf9f747ec54da4a921872f83145a3c0c2024fa0c3b0e72af6cad639fc7bb845ee67de9332ec902a241d8ee4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h199b3abc049db902290fdd581fb56ef64d7bdaceae91786d065a3c31ff8c150eb839345635f47cf9c7de7c8c323af68dc0e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca33ff86f5dbd996c8b88249a52680b34910a3c056c6a90a00a054bb71ac0f4cead9e8f64c00886fd5fd998865ab2c5a515;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4433cb4f22466a455ad7cd754278a437447b2b448510b6333a66f92f260f95e1b247ac0bcf881d9f3ade7adda570bd4fd5ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cf45ccb9d71105f1dcf1141a718c1b0ce69f489abaf8f07d1c1b24e5b930e096e7e76a48007b0787acc009300f61c949e50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1843598221f5c9b61bc71fce4675a8bf41f3b05720a62b9dbad02b4fdad17d8467f5dfaf012735b4c58ff77659bf0d23f22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h993e32b2af6788d1016b1cb0c90a82b0ed5545d852f482d62bf86853b4aa8e3d6f00b0c12df150344515c9ba0f5a88467511;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20b658a01b5b64ed7f43ae3c6c5faf4311d6f138c4607d0ebc7749cdd8276d168db10fe06852a038533e82e32706d2d91de2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12896abba989beda608cf6045304c441818de116f00ae9e7711b9749893decd4c4e1a84130ecca0b485bfa347f7ee1ca17a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h426392631162fbe9c15528901fa047f092f013f19c4022582ce442610e86633a337abfca075a7345e4ad9ce4291cca724d5a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40dbaa0711abf42c6de12621fe8751f8f44b6dcebcaf32ab681548f20d48115b02bbd05f365897e024cb6c3248998891f3cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ceaaf5249882860139103d51c95f7ce0d38c64f810673e882db77b2228e3983c7886feb6f6cb6f47fbebbb3839164b5dec2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h351381ebf4b5bffc7c24d3a104e66225bb4d0db58338aae0eb005dd839e49d5e49a66c7be700fa1d40ce624d48ce5af092f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he73859246bfe94a8aba9254c193c5296ce33216854db0978278151c212891d3f6380beb9557d91e97d436c397bddc284bc42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9116d0c8b404ece68acf33262c52ff3de7037adb4d29ce583eec44797b8d63bc1a8d808b7b2b477ce772d9c516b15f0d439;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc48e7058cc2e3362056cabd63af2a970dfa0154af6fd473fd444d077f6ee6a59f42cee4594b7a3943b63bcf09b17d2e843d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11fc8b4bffc92647bd1a74d1c677774ead7a0f9522154018b8849c8abd78ded90406da2c9c8190d70fd1c509a759c09ba24c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9985a6f39aaad3b92c87ccce542a2076b09f7e1be279e1aa7ab0e4b000dbc83c0931838c36565b508cba940c128556c065c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbae3050f88db4b066366e673ae761c36ba708305d4315eea6fecd3a981a4b887034f5d74105edb4289c3350bf4c3f6492c95;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd986a407e1e4c7b8bf38eadaec411eb2909b18b038c28fc5cab511bc6e0811bfc52704112f0d95d1c8eca0366c4d4221b1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd8f6b96740dfe2794ee5d4a952ff4f2183c62c6984d63c68e2304da08f6ffc94b2818606e3d1cb071e8ef4d36f52d81e637;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dc54b204b8adb9958a52a5d533c348e61a06367a7a8f2c4ff5a6df9d088f183e3a278efb3cfd841968f1d82827245106dce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe37e6b71b041adf0c32bb77b95fe7d62e7f76a885b06a002013407613986534277fc6fcf784f704e73e713400ef157745a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he591eea6d8c15b0c6036e31e0ef57115e9d6b1bea143f7c499066e732a5ed8f1bbc48d94047853b3a23121bc2949993d59f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde90752889e93576bbd5872ee742fbf95a55c4ca3dae497ab2f1d8250be89449c4e61a5fdc9c06172b31b6ce4fbee9e3c0bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80a16491d9850dfb56ee7db8c276be3c061e523c5a0911b656bf87c2de55ab80ae71def0916f38f29de687d79db150559229;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha006f8d923553d81dbbe994199e37c11c35072cd660bf7f1e1c9d1a2fdb5316f3ff40c6cca7770fb6269f0b133407dfb70c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8085f18d0711943471909e1ec981385716b8476b5d4a258a135f3aa8ffd72cdbb3aeca701873d9f0f745c35c1d49fa874a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9e58894450b90b89ef68154e6bcd5ef76af0c308e59287023713328fd8161084cd542bd62c07dc47099dedf546a8ce09ed2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26e3d149f32f3adbfe4a440b990d353effabb77fd5f46a939713e2e47fb713c8acd4d0f5466216bf7b30d94bc0e694564614;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0378155aa68dcad226c09d8fbc0cc6fab6d0adbd73271237f17c742a9ede23d8cf3701e283fe99c42cee9ca189c151bf88f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b7b0c21638ce228639fcd0f025ced827eadcca81104d2fae8d572dd0e4369bf40ffe9cdcbae6e16a04a207708cd93a79d5f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74b9e4d7799d7f5735439b4ba403448ea894fa2eb95607555b82d4093624441543dcfbb0f78810a046fb620e38d36b5affae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d0e3f7ed0fbdc1a5b138ed9e26dcc5ba8d97a3f64de5427754757cfe0fb29f6e025bff34b880acb3ff7d22d7834817e5111;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a36cb6781b5987e3c5cccdb643bff3d72903191497c286770dbb1227bc245f7674fb509d1ba6b55f903edd36cbffd74e579;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha838445d94648d1a660528d92d9b59f21799992e67e24f2aed5833db0bded263d7928cbf3df023dc75d5fbc1cff37699ce6d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf83cb459f99a0d920dc5c87146dc856ffff34e7d87328477a212eef83a9500811e66435e0c5d9e615b4bc5a67d525c4cba9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8984d0982adb821a08ff69ba2df4c2d18b0511bc15b971731c3d790f4cea17cafe11f9757327b8396d0b3ad4aec7d33baa57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8517172e2ebb30a8c5bed18db01a0db9ea38edff5a924d20c9b80f56b4455ac45735da87b9db3b4bd99260ce19d503638704;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5659ad6c362d7f0833312689afa0bc19a5fb58fe76f7da1af8f3d0b56b03175d0f8f2ef5c3d6c719e372eefad0cda6f65cce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e4b049657296a9b52e55b487c6ee54a6c256ee9f6c5da56687d6a720a33e4e1c8277a548d392adda3a4a48c11d889c097a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he36db27274a78a35b11c4fa67d52a90c99e4b602ebf37ea8f2c6844e38c787b18d9ab6710c46847b42f1cac97307c18fe8aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha867ac2a2e8618c58447113d38b1ce0a685e0e77b1891f970380c060a5754ac34fb9ff952fc16cccc2448b1fe4bcbc4ce69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf656edd0f0b5acc27153217cfb2c57c6739b2ee415e8882c8122fe94559c7f991e6634a1583f1d4868427c3458583a841a4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fec458ac22aa9ea1410a4a2be83b2fed19b3feababa3c4dc9f73709fa0c573e22593a638c923c4a0923f5019abc1faa833f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1dbc0520a0880b6392b4cf0a84e3327b8a0d5771916d0535fd1fde5e7c7fdb4c9ff1d774c2a0278bdee9d89ed6cbfc6b0a69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1b4b494f8f0042ae91735c425dfd389c6b5aae6e73d05265616906782dd99655bb9cb8444a835a0fb71b17f81a6441ded3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cb792a095364e6891f71350f5eaad1e529157f45b4473ab4b4eeb4b84996d21a446836a2e5470e0c253c0ce14c4ccef2168;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba4a4b84d8c542702a52546714d7198821ffd13bea6ef70975b25627bf1ca0875f18731039812adf34bdba9f3770e51fbd6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd45576a28b1d42b75426d858c0c4d8a212e62bcf852fcaa520e974dd63f16ae09aacfcc5b765dd16ccd50b19ada259ed0afa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaf72c48927b2703971126500714cb81d74c98aaba3d928f42c4679fd566bfb33901da3b4366acf48df06491e5f34fa13c5e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2e4bcb0807228f244f4a79ee8117d185d7a4d080b5011afcea9e389c30f2a733b9f4ad1ba40aa59000380cec85e921d9c18;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he29969a7ca2e624d90314935c6703c6e7394ba803c7a21f0a30a6a825fa9a9c4394a3c8bbd97d6fac1ab2f012c91c8e8d8ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71adeb76a7e0f3f5833f71a0fbe083f426ad151e66e91a3894f54b5b98fb043d7af1fa75a20c9ee6e5d6a7bedb17b0fcd0eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8edaff3ecb0eb679051a738af40fa8411401845e5ea408a73e1d09f0c97d89982a808dfffdd47e050579c835822dc665c90;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1310821e7abea26d6b973abd94b9a5c5020ccec8314e991657ed488a2e31d9d432d6792f72bf948830a0d0d2f9cd9a822cce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2aa5d3b192c0165d5b2d6bf55531ef236eacdc04f7bf639c78361635cf98e6277b095c87d6c8ee5e00b1b67a52f66bde9e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8127b7c0667c6a3f2cff850e5a48d9a157684d1aafca2bd2f5286340c80be451cf362c295c33ce3ca4fa9a6e1b4f2abb3f29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32938aeddd83b729a2b0c80b1dde6d8b3e283c016b967a3ace85dd28fdaf3eb28818dd55cdc8457f5039b435beb04b2a169c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88f47207cdc7f944abce9e02fc89903800bdca7fdef246fc94077c5a6867bf29401d8250c0e7b68e60b18bddf524c8d71e86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45ed281678993c6ce1400ddd5fef27d801dfdb61cc2db0688bff52fdabfb96140c96a819274290a17790ce5b2d2b5fad2b63;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41fbe295f77a77fc85b29e11198b1c535d80f088f98471c474143d5e217dd19680532d14827e17f19c45705091736d8cf4d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0fe0f46609ab268cb2fdaaa14b01ecc959de6174bf066b972430a7c84020ce0ad5b615d36b9172febff5aea01f9ff12805a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc70187221ecb9fa63eedc1dd9f072d7f0f0b06e773ef510cff4b5b8c27fbf628cc2de314d4cbcc83c7dfec0512cc0805d938;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60dd88e32d6f2b55c32c13520203c7510fbf8e9ad71630f9970f355eb74ffefd699a8cf0379c9b99a83cc3b434a1320e1647;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ee1333652d9341e00b68922ee9f5bd0698ee186abede625c8a664b616cb264d298397113b48890dbadea207d03a1b48e169;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb7031ebf68f755b48e1161ddc50e6612ddb4ed2b3ac0b16c597870d545a3098d99426ef34994b47835ab1d20f981f83c361;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h466513696a910f44b5e4f33b82472287f0bc600eaabd40aecad714e415383c3cd244618cfcdcee9b292fc95ce0cdd0ed41b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4b2d34e24a5096912edee2e317af7306d61fd97164a4a6ff1fab38571ca5eab1a4a3fdf8fee2ebf2d60e200b70d9b3bcdd0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92b59daf8824043e302c45f9cf8f3644fcf0124d609ad60944508d7d946d501ddaa5043a16d8e9f84cfc399f5f11b7ff81c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h679917f3ce506a815ccaa12b3ae4c86457c0410e3925e8cda8030eea22174f2893e8c671301736877047939d8990630920a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d887a058d6b9f85028f986ddf0533959fbdb1a0d7c96a1987696183f63fc12b9e9230a99bcefb1bd8aeb79354221d63b8dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ebc5698853dc4f76af747da3b67248d018e798c1be06e39bf41c6f4da5f29ec9afe067ffa818eb1b8099e3990d878db0493;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf631233bf09396eb09822ec86d3bd50d7b856c3d484c7e95fb2160b6df2286eca092f467c91517fff9c863a700c2dd2ecf82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0332430614de6a617dbc4209a1c5e89a6570e25c04196e62b6b89f69ff9dcee940d484051635d9444104f6240bb69e06ac5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa4990511077eab05b2deae23487cbd479822e7728f00d6c7d842667327d98c22c963770458c76fe44d7b3ca23a4b311b4af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7797e207902f6820bf5ca56ff519aff5c56a08c5880ed521ba99f52cec0ce8b005e52d0e1095e9757cef5924f604ecd45e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e72ca35a249446335ea29484841b3e16314d71984f6d9aa8a54bb8ef7993d5081b22e7b77bd074675065cc77f905f097526;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d02268da99694ca8c7f828c177897a2e4e4cc60f8973116d80da4ec1fe267bfb9c186e31f81631c410a1d26ebba32930fc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63409bee70fbdc060379b99012a861541e7d96f33c192020a96a35400a9221ad5d5258de9ac6000a9ad49a860f8b5a458a70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53b439b6b34bd930a67fa1a2589be803293a80766c38449f410f337fe4ec924296ee324329e7d2476089ec1b08ee681129ec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0788743705c099e994ec3ebff9289bb2643a702d616090fe56ef7e01ec33253cd31e26930309daf9eea6a3548cb9f3a5aa5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h597efba5ce5f236c70ea98ff88c3073ed1cbfa99860724bcfd0e83462b8f8949bf4a7feb85e8195ff0667a2d79868660866b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h227431a9ff7528b6c9a27d294459633be0115d99a5f5707c7f61fe7ca15e421a849a414a5c435ef975d424f1315279b7a55e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha14c94fe9c79ea016e1a8e8a7e309bc4d85d548b3a25ac5fa35bd48c26568550413136caa6062f87332199e63537b4b94413;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h812862904e87234d80e8d98e8e3ae00e30cc5d3eeccc6489e9beb7d42e306fee82d930fdea828eccdf2039ffa5f420c02261;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7678b29d7743e78fce0201513a9c7878e0fe3582ce1262f47d479346f7ffe4df1363fa890300b0901232d6f2bf3eb5f3f3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h695d4e5ed438be9362d482a49820888dc8a4388626cd85cfdcfb10a8bce2d4498a593adf5cc8d37f25d61bc24ebd4b73f175;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbee07290bb68e6c10aab5ba64801e2cdc72f967c15a5a0e43904b755c348796aff12eac1e237baedd57a64e33dc7e34dac75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51d57fe14ce4879dc7501f06bd41438442af590f501f4fc92edd2c34e1cbc1fdc30dbac541a1d9a276155feb2dd04e1bb3ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14cb0308d9afc02b4d284f24bb898691bbf75745c83d043227ba9e4379cdeaf195bc4b015af96a5e03ee704f4572d852a134;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda7d99bbb4f163a22c77e48506c38bc54b7457c241e1958b5b67056720d2e2c7e04784104750a664f8fa25db5076c87bc772;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf712045f945d06e401392260131d430373362c075c6734b376492c3e7682f58c6eb484f317fb36d3230464126de2b1719a9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcaa4182d5cf9b6a5829ff2aa52dac3b5323309c5363c06eec2a011a5d2ec59212302be5912e9367ab2c1628562d9260568dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc702a33bf86c2c74cd1f259a07cad465fee163e40b47f39fc79e9572917c4813d4f2d149d0eb421616529f13cf0470bc481e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc943eecf9a090855a719cde963344060a12338ef5859e54c260c4b821951d16fde907c0fd451eea22f7f688071aa2042d1bc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb69e7d65ce7c502be9149d7e0ad529854ffd88111423ef95f16d9b19e4669acc9627146344c49738cbaff4bba202b7729f15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a211ea877a5b491d876aaa3634b7be98e7dd7b5a2a358626294a4c1b6d809378c56482d067b314e0c056cc24224b04f59bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d029e41163a057ee6149c08ac537208527e4bee8238180da9ddf0e6d4bd55e3afb2b39ae5799140dff5be0265528abfff57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he22dc95607863e70eab4e3cb3e85c94d0c513faaaeafb6c0fdbb4fb404951ea92a8e15968147cac0d740a7d542c137ff7462;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd25b05491c7e0df3075217d7d019cdd731958c58074f58efe504eb17cc47b8f889457ccdf728b084c02b620a6a0f65e5f86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d4e9c540502e4e3549d189bb20a1bb15f568957f213c310a39d7197af3f8792bbbc2c4fb37c71edc7c85c1ed440e8f10375;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h253cd8c55c4bcfc15f08d20ffe249955676baa8c9be24b9525865e8b67277ef126d0a49444b3d9ce6f76aa2ece332dbea5cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h897230758e5c2e2015f205539c234153039c3b16f2f1d34df12ec7f63266e316d022ac44678423ce42644d85c48e3715e82b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97d30c4452efd981b2669c261a0d0cbf3861989ee9b7638973014e67f3e86e9e783c0b896fb13f939e0a8dc2f1579150f8c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5d605bfa892a39f3c651088c94ce45902a730bdb9f8ce982f9855f9680911eba7b97239c91947734548cbbf81fcfbf2a41e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5a34216cea4d06346d68410d148051dcb9f637642eccb555a07d47614f64301bcea2c063ffbe01587305348deac07cd632c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h290e70ce84fe25f6c585a2cfa8dc43d228073e6fb616ec4a373d7bf2cd0bd3f2c26134f5afb1c4075892c37b04fe2afa7bfb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc8d7e82ee175eb44a9a8b205751c075deded256fb0998e753ecb40a4416920eb0002050133272db83bc94e1a6f46d23fd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c0043f412ad3bab44934673f1dabe3ee23f57029f3ca3ee25184ba7243a37fc0b092c0e91f3a593993caf8d6e44e00ccc3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc135c8f75eda7cab7b689935009d75a04de38fa2e267660a5eae0040cdf0c06346a403b19624fa283abc02e8cf2f9f0f4da6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haae0fcbb11a3f48abdca1ce499e8d34d865c24c5ee708dd98ca8cc9b3dea710aeee6c7b59babdc584d9151e9c609ff3af9a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f2f1016f89c9fb4f4d1857a5804642898297ca69e8ea3976f7b52736d2dc42db7a7a48b5d419496b46dbe481f9fd881cd8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0da7627ce12cb8f6d52b4b1c279064fd0e7c9fbc7498410497e37afa7bc0ffa4b702b579326e81a45ed858f56a811e11d9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h604b067d577f4f92892e0f607ea6049ae5a2ca3898cbf4200518697b2b9c4a30ff711255865b4d6eaf8c99d6a5036545889b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37cee7bb80858c5cdd501d41e11d4fac608d05098ae5c34009d0abfc72da9e57c6784572b088ae687c1fe37a879c8a1c78df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff246e82b782dd8ad2a626b71ebc876d210523fb5c0ef68b2e0f1b1a9eb4e101f3890b606752d862112c9c2cca55222934a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1b3356ef2cdb109994177c64d36d0eacdb818b114e5ed8a0fb69dbef101e5e87a70340576ec1acab5db7f0b4e328e6bc9c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6d04930f4278b3330f02d997da2a434b31de4d4f06d1dcbd9196335cac6e336af77d315eca5148dc90013a73ea09388bdf3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f0fdf9eeec71febb67194c3f1c2cf12c8c90c1b737cf0d25743cfaada19bdc509f3cb51372a2868e7ea98dbb7d4b07a6e48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19e86544be275d90a9fa9f1bc071fb57cffa1c6cbe127310665bd6e33b41ca1911007719775d0195bdf038de80b18e2482ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56e3cd0c7c77c4493f045e4d39d047ea2947f9c437874d2a105a917d751b2c88ff8b0537b799736508495ef5c78a419269c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h441d241dc8866b6541b54c0e2fad2970f481826fe20dbc5ec6622e4babad9927a74d9b71023c45e77e9141a4cfd673cac79c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd16ddc8b44730cc3dd6166b5caef1a140fe7758fbc8875ae451ba7af46aa73f6a8e8cdd86a7b4ea84d94a213ec9078d57264;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f67f52c2ad8d0d91e7fcf0ce1cb16e7fdbf38e959c131e659d5b6f469a5c924980d8f9ff10c5bce144e034ca09fd8d6e4c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he425b0083b75621467c8e92e8467016db17f0a33ff13bc77342d208d62a95b7700493a529a1fed929770e1d875e05481366a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h145fc35964e4a62a1c8b4e8c84a716745b4ea6096515af2822eddc0bbf99c7e94979201696df742b72efdb8350b6e763705b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8ea6e7ae19313bba622f96066d45cbc2a4975d91067c4e4d1afa41f0d1f145de52e78585ee7f718bf5ad55138611d73cff4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b56ee3d05b71037021b2f25fc2816a25f1841fa8550710be058c876d6cbb7ab36ab05bcdae3b3ba6f1380f45f049e89c101;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4532a037df8a0067c0144386c91a13423bd849182b9ffdf3d9b9d7642947954b8989f08855bdca1bd76bb37a19fbf2d1389a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0ce74347d43b462f77c1c8cd59a58dbf758522f2e7f08956ca879cfdb439ea8763c481c619773c053a9c8a4a6c3afa51474;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a3944077c31d2e333f1b471c92676b19dfb5349d46d50c65197138bd9b3de3f52dcc704933aa583faba4dd1dd292bb08904;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44df08132ced982850cbd6a5fe5dca246877741d38c363312f226c4dce5cde4e9f5a63836b84eb900644f96e456054254d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1246276077ad4a58a077c6883e83e61357f6f55f10f25dd16d644e5aa5d8f44d743eb9f1f6cb120f4755cdfd80afd470ccda;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68dfd27bc61b07cbe49eae2e11ce79bf66b6b93379cc1a29e21823439dae200507701796690fc6fd144a89b14d811fd13024;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15b5d930139956697e7b4e8b85f8ff4887cfda9a8e7c902a7adac2c37d6d3da5deab442744e5765cd8d6785fcb1767f7a30c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8c07491cd9b88e5a9cbf7c864430bef50ed01ef2068be80dc7a0e46ffb73e020bebda6837f597c00303a852787bb13f4f2e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55c400b60365ce4da729c0c3f745a95980e6b42ab7e412e269ee582373f293f65028d55c20c240ed587b98c4a835575639cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1a1807a30792c137cadc21723d5ef4360266630bdfe7f42f2730239296cc6ef8eaa2cf2c536a86ec964b2193cf04644a559;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf320409ae23dc5cb6d53f3f0f19f3695ca521c3343792c1e4e479dec539b0c6df0b4b4f67237595d2fbe56e30a4aec22fae4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb16b4621acaa5689633b357338ca058e5fff3206aacc78150b850af79bcb55b1fed9a1e551ea02ff4ea09d38840cce1eeb5a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32df26d9563fab29ef199fa571a45877f2100976a62ebb4269f33ede099a168fd68812ea32f5eaeeb0985cc30172036f3cd0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb88d96c377cb56866f2d2a6402e2703b5ee30e5f9e2ca0f38e3a41086971e39438fd86f745aa8b22dbe3f231ba5647d2ae22;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7434218882c0f8009078a450a293ad03747172b6ab01347c7f74050cb18730671f4876e1ea2c66ec81445b6e056254b1ada;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5b59cdc3dd8df2fef7cd7b78b554abe0ae333fa2beb7e596e1362e58fbaa64265b5376ceece82062d1166ba7668660de206;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22f8436c701f5bf3df9ff17f6792be7653fd6188441aadf019b828b151ad732629ac678d83c5d25e965d342b8205be879f2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15a9569d5bf08e837af2b9d567d7305b663dd6c607208c6e0164e9c300d3c1430a5b0e2bb99b226826b0362c706e297e9536;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he41685af1e2431c63c393e8d533a1d149fa54c41e651f5456d5d7e6dc3a663bf5906eb00a653862aaa958925fa1f09721591;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f792fc4b4167830884211c3ef4ee78e762e59d7f27dde2aee1510d5e3b335b8e8fb6975cadca5291969b35f5505c662b841;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5632c6baa7a1836b620274acd2ffa2c78def879a567ca8571f612c2f425a026f25c06aea0df24a1670b86a70218491b35eb3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce6f72237643c59f8dc170173322aeeb7b579363c6a9b7bdce77472b79773282a1f9d895e7848ba3e2d40eeed39136e4463d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee2b6a5f124f855e9eb0743cf3f1307ffc1e3c42dbd665dc2319eadd72730645b9e75c3faca2c252f5a8a96d2cf78753e22c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7619f04daf1f71e92b83d9fdf48b644120199648abd65d0750e379f2925961ddc69545649511fd623cb4ebd941781783ae4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bbfe6881f9126cd03c3b8ba4bb0f48493012e45650f4f863e3a448d9ad765dbfa4de4235f503336daf50f75cc36396b0215;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h704b25a669aef0a1dca84d7dcb0519f1cfe214f800d52a0c6bdc0759f05379dbd809e277eec655ea72a2df159088f0282b66;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1df3b1c47d49bf3e2ce3affaa0cef7b6ee1005405b97fc236533ce0aeea451acc08b57bf28a5700dc90d870380ca9b44a94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h789d791a7c2acebf36da45165de7bc1483be7063184f0d017b6402589a990abc28802f82eb675645e38b2b9805276457c83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he85e76e0b1dfb8512aff66645000f455c28d0ca71881d2e693098cddccc66402fb00fafad428d6fedd47f1ae317814a577ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4713682bf0a247e0f9e515faf4c7b853b0baecd5c0876c42c672a3b38c65f6143e155ed494efd719906658de33eb7474b0c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34968b96e7e66db67c6bcd6434f445fc10bd38b8acbdb6c431e002cea0110d62b019245582f41cca716e958136efc1bf5909;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5c0b1e2bf096fda6628c8a68425a4a28357b31412190e4effc85ec8508b03310f4b3fe121ff7c0f0d15943f7190275c227;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d9f59dd16dd8c80d4fd7dfdd8f37b86e9a936c2697caa02dcca20c4e72fb37b3cb18490d94b7d05ed52379f3aeeadc4901;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h157cc5486ef5d100a39bc50d01c59d26de6b7a3095d0f4ee5ea0f38a0471e0dc34e682cde2277cc88cb429c0ff8c2470f0c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc500992136cf6cb42de966b279eefb5df898d94b92d35c22694adcc5c83ccbf0d8416c510d98d01b4cc391bdcc8c15effbf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7132d289182c8b19d2fc0414007418ae235c6b512cb01819ce2c258039a3120d0a94e3fbf9895caa0cf5b1b1241173fef308;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb397091c1730fcf134805f878e5760534d090b581b3791d67b769ee103a3ce923ce0810b96028c57b840f51e667527e19f74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27bf5f54b6493c8d438fd6d65e11e81e21e235bb586c24e95f1db908a01c2c002f70c602cd1d6300eac00adb9a9ac2343544;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha84b932e300547d23ef13ee1403634bfb60774a4eeac5b4a886b2a53d65c0a4792c7ea13878d99f005b3744d8f6c9d160930;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdec71f7f4c29c4b1e25fe388f08ca80a8fcfb69cfab4977eb4c9f30572976a202ba6d5d6273f868133afcbdeddda237888b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3396294fdad8f6f0feea06276cec63642fc4ed45415265b84f1a8960f9b95ac08579a2f60e8b64e246ff72b5b6ec41972f26;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c575c013282538ff780deefd06ae826f74f43c72ecd04851f6503619240136d7a5a345c03633234eecd5063ea549a341d8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43e6b32ca4bf64af6ed65e1ae156a00d2d4f84029425b244dc6bb804855711e2cf7121468ed504cab4bcdb0bc97f5d8fc54f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1380b9f04e8ecc6f94ed7182a353ec87be21c7caea12e0df279b026091f6390518b8d918138915af5d0ba0ee8f790e89e3ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82ec0e12a436c6a40c330b7a7506b6cc1c3486eae6c3543830c18e8a03ec4663ec528b23f375025e16e06a037aa7845625c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8000347bc46547aebb67a6f6d947519c65253b927c0a4b3a171e0448c104b513d75981afe3a20d8e74db945a662db11e02e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b5d19dc22aaf432d0deb953ce15a34c962d6a8632d7ec0bb50ec79715be58980a567ce99d56c61064ff1b764456fefed82f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c0eca09061577d1f3df1bca45c58d63dac8f2375dbfeb4e13ec32b4d372d06a2c0d7ee544919a1d4819487b98e51048331;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ece3623c1965e696f92afccbecd61daadcfe6a8edabe4f79078747a3165c5949cd4ae8696a68d0b8ff9a82b67d17dacd7d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h972f97602234cd3bd3f4120f4e594f20ce540616f785d403d60d1e9aa01e08e1cff3837a4e9edb84fdd5787ae8e5cea3d376;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c08718d17ea1d4f39c015789766c0f766691ac62143b9f26d3fb3ceb528c87d907cf686a60dc92d72ceb61f0e7e31a18fc4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h399fa4efbc18e675abbac976445eaecda333f2294a807d8a4ea13987c5591a134f37bca69f7b871f4ad34bf6bf03d30f642;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h929e13370a48691b3e934aca4b4015a1e8d9848644d66018b87a0325c727ff3b3813fc0c0d57b3d43e579afa95072c9bb84c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65a813641df1411aa7cb3d129bbe5388f92fb6bde5aec5d952df7b75d623888c038c56b140aa77aee2ef9f98b5f736ebca1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92453f8c1a1aa537b4485cdef96fa9e160fd131471f165087b28daaa8ff4cb30f9b531a4ef0cb6ad859eed954d0ef7ce8d25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h299a7f1c404bf44201edd35881f320efdcb06667d26db9cbc67aafeddf8bbca820b3a97f2e25eec2b487096c70320060bd75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5eade9d1e9d5ff483547311e1cdb0266f50b4c898238971c8d1c46b19daaf94115ae584ca017c8461026aacf43d85d305f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e92ec7b7aa743316af8f9bee68ae76596589ed72dd5b511fb17846e150bdda52e4d7b0aa74d924360da08a21373dc20bf26;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e40270c5d35df4836f8e7b9e3a34ea7f8ff21df2631b00d9499debe9d2aad0bf475c33c348239bf662b2b589348a1124833;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ed2c7bcbfa62e6c1b2469170b039dd16924687ebba3acd087064efc4e82e539fe2b0cadf3dc5853ece46de1f0b27050ab0d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he81a8086b90077ee7174f3065520ff97d3ed68d16ca727f3cb1ab5a5a5ec2bcca158c4c8ea6ccd458e084cb1283df623260c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7968abb25227a0180c179ee8a0599b8ddc7db333f3cf85b35769c982a0eded8318ba15f82fdf496282fe1e34ec939bb6350a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0036b7dc93f9531e1cd92860756850e479e61753faff264ddfc1bdcb4d147fddfcc30b2124c80bbff9ea158b66ddf61a1a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb38c0356e88bcf1f5419332337340db0ba155651e202ae21423645b63fa181788e49311569690cb2f7e56c729e264d73bed1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h545b528355fbb6b48f2bb00b16297fea114358c982e37b3e61012853322c01fc94a61ae71ca3f64152c3a35248ed857a97ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7bfcca75987b91f1410f21ab7aa859527c9b95fddc52a6d5df784685c1ad909b3f852c2f3403175f8789e3d87b615319baa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36ba407f0084065c408456941b12d00666d65c6b73a50900821b9e65ea20a28562b9613119b08e309d937e14c1dc0340f06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h719dece92dc499c5ca41dfbfaecba85266cd4c4605d0a483cf030030bbd183df6e2f43a5d5573dad3e8e4aa82c7d021b7e08;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1be1026a763a7450d39d4906dc9a7dba24e85054ed41a57c633a78fe7b84f193570e6b56508255cd679e46bc9e50c4651c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31ad2090c81d2a864b1a9ee486aa7f5ced62c42186531af202c4cfdb18100abaf6acb471b1a356ccb52b5e876434286e503f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99e94d57f3d0b34264f74dbb468213f321a9eca80b9b6bc4bf7a793e6d87579bf98f2bfa7f36920f241f2af01b78e07090b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he13fca3d65594db1906b88fe4819c104ab0cbcc6d92bb9d66dba1b02dbccd37cfcd6a636d5d234af3b6c0f717bd75eda85e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h921f4c6ea09d3f7e3f887b5887954504ab0a1d318f7e4ec504437638d15174fdbd7b8ee42049cf441d5927d5ec1cc2a9e394;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d7fb55803f30bb134daee12e3804e6a2746ca9ccb625b6a28c56e49da0d7a104f8fd5ed7fa630056d4ac7b602485be4420f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f609f1594cf487f7b3d8d09bb3804d7f07c2452111ec7a634a84272edbd30371f7dc1a6e892ba98adf5982b2b39252be9ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60cca6e90b2529928f4b760c4a0ca159e182f1dd54bb1622eecb667874736151182565271cc02d87c6abb540dc84bd82f534;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd2b4dc2ab74aea905fdc5dd0cfc4c0a890eb07666361c8f4328dae8b147c6e9b18141359c3f703db00362f7e3c26e295aec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1603e2f5c2423506ab4e7c5f01c414173e20ab3e1cacf9c8a0aa65d923481e86b2505f2bfe1ddb79969ea70238c8cb871a64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd59ee9ed61ba769b4f60014530f350679d864cbe8c6916e58a0f70967714f0c40e59e147b2d579da7cf145742f558dda0079;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h376b71e4d208169bf1dc069f353902f98b9b336495c7389053347b0293d111bd1830f33864898f885f4a2e3d0060d834d7ea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf193a9f5eef33e876ea61ca4c128e70679b0ec94e9c85fd420e2d1e443e5a8179825d81a2c04a82e0a9448bfe44ff7d45174;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77b0ef5a5c239742eb9b79042d5ecf13d860671ab00ed03253503c4f3e2a523bc8a5cdbf2e62d48442bc6c325b7f225b9da2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ffa3bd1d201a4bd36e2296343bba3987a7f798612086ac703f427a63ee9e4d73e0c1f0d18b001ee9e67231b5608fe76f1fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60c6c3eaec9d4aa80c8e10c34b96bd3232db842bac9cc573ef21b21c02e0ae48741eb98bdd82a9e8d3cee86a1917338da7ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cfbfb0f86752eb6d44401562537cd1c80866f148a4fd532f226f3830f8f3d5ceca159824f43992b42f3138fae796b6a71a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87560a821c4ba69d6b2e614e097d1fca77980dc48d6ca805edc4733ea3c8edaa98be8ef824ca271cb867118abddd38b19ae6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71b903a5e5287e2bb1e583c86ec54f8c04ea762a6651a54c38454b4070d9d8f54395b1253a4a19d695e5745e233b8bb0ac49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5085c3b72f3274088e631bff8c5ec78bdb104d204e7ca2847e74080078379ead346c493970ac429b3d14740ff54fc2444a91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18eb5e56722cfbb2e093bd5c3f86b2bc2b8de6827fe8e325caf491937d1c946afce9d25ec39bb647eac759ba1044ca03931c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8314110b1db1e31d6bf34ba5c49b198e14ef79112f7dfc7179a2627327d712fc6e7baaeec85941c65893c99ab51291c7f305;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a4eb0d4bcc00184b73952051c1a1e1dffd33f53984274917c0ec23756f4f374cec9f34daf7e418637d9f68c424424086c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27fa9994346b2e4bd81d25e7005d0700c1a12859dc8a64b1ebe6961ae47db0d6cd9e189d17771d41efe3535d10ed2e9b39d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f4e25817bfd4f01b4f7d7512d649af4a8921ad7a0c9859c0c6cd4974db1352666126dd8af0d48a84513fcc9aae4f66b9ce6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6deae4a6eabb9a93cf3d92c0701eb56d4e0f453fee13f22b23bb584ca59559757bd756f372ff82dd108ae87cb7b2137a93c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h533388ad757dee72c56432e604bd55f93abeb02fc8b20de2713d6e9de2da96ea56a8f36e3c7bcb39622de23a155276d74aaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba3d12d5d5d6be1676ffd5d2dc8df165c60286fed5a5f27085c6fe5b036e3c97f8a6cb9bd422037f7be38bc685197d8819dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84b7e70960d06566e0c69a5b55dbba60ce91ab0c40ec57535156a2351ae779311972950e34f2f5fdf6f856fba1d610996260;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15dc262d430b333d6c2f10d21ac48c58ac49a91d5d94945e2463328b5ecf4ca5bc39eb285118a1d0d1b5f0810ca5a710ea3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e93a1d6b36258b0571f10a96f8bba3dccbfbbe0e268b98240d98877dd1fa9ed43ced7cafbcaf8645845cf533474e36b5971;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24a15ebb2c75e4f2618fffaa74ab3b96580589b45e384dfdc38df90aaa8c1eab5bed929545d2371077c779524a797fcc5976;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he22a05467dd174036513359a92505aacebcb907a327883bed8e1079f306b93ccf0f47d67686a5336aca5ab7d6f53e1744cba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c43e4bc6f79dd7a58d0f1c449bae319d59804fd44adfa9540c98faaaf723278653fd8f13d680afa98c20305497a8b006828;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83b6bedd6d532f50dc6239b7e3e8b47b8c828e14511bc6156da6fbf56f3471bf3c251011af08985c55ff86c08fd1abdafda9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb623befaff7ab72a3929d2f4ddc3cf9063233883a277a607ce9f4fda819d3910feb569e7cd7d0a4e5730d32932c73dff2f25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3608db675456f1a81490628c45d53278ea459a33cc494327ad37b89670c9a7e379f31ca834e770af04b5b00d391f47bd42a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87b9c10379400988324eeb477747c1affa0cffafb60caffc579469c8fe4d7c83aac44120caf454732a04e9591cf5b44c9145;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68c573c598ce5c9c739da9926b8839f025dbb3ca0247763aa868a77e351201a5bc93eeee7ac906be2229178ebfc848650ebe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6366210e1095b0f03ac7ec19ed31afcf07c519dfb6070e3ec06f6f43036f0bd7076d5c2dbe1bf844fea32997b91c0329b8c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9228e8b191cae81d254aa55e306981d1c158a4a12ba4ea9d9b878821596473bbf45953978300336497bc14d41bdade4cd288;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h30c8a783680dcffbae50c57c8c19d5bf3da4128a9b24ce655fcfe4f5442447422c75556c967fe8953cc09ce829202c95623c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h815466319cb5c3ae299e6f129707cfa5a656c24443e78177ca4983660694a3d965e1603f519a9a02047e2fdd19be6d25f73;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h485a360e2e5ea5c0cdf7784aa6d96aaa8253d8f0c6baaa2ac40703ae6704eaacfe2a2f5c1f7054ae58a7bcf5097d34b31f28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdb75882a9e059fe7478bce35ccaded0ce12717fded4280b6ee99cce8366455cf5adee36059e38cde1bd29e077083498d25b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56a643c430c8c2e71cfdaf1ad8305dfc5e9316b6c407803411aeb6f417e78339375f79ff0a96f81ac9b4244b828d46efeb65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde4416dacf58105966eee235d68ffdb86d2b4900f179cdfbcbabc7c25b292136141fb5909d349518b61e9e83f0d466b09400;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc86fdcd6883f0216cfb89ffd99eedb28a28717a6814a7a58025e98d847b6fd2fa8cfcd89638ec169a4c516f22903297191a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1feeb4d33df7da5836629f8c0d8354b743ba77181c73ef343c1d659c694889a75fda81a9829c267ff82c1592a123541bec33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a979c54cc177c49dc9c0e441680256d0abcebb9065d7e1688804d6c6b3feed811ae7723aac5d95907382a3d5b12a10b4920;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4053a8b9041aa3f3e2f8c4176fd33df2e6465b6ecedd5cef870d1323c0be2870e79be60093718a7ac443d97f730f5f9890c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1060833dad87c55213577a9e45ffaa6db073d7557a581867daebf430d399739ac2841ef2bf319d25220b05fcd4f2a6e42d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc096befd1e228d7ada37091dc0ab0d482e6cda9a06eda4b6a15b3813d860e4464f5b7cc20089f354a4e9edcbdf0f05e8861d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb16a7c518ca132d86885a1b1b15c936ffa159ecc3b9f983313234338b110a3f89a3b1be06699b9df2e6bd2abae3ca72e9477;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb54b32a084f964017b127034843aaa570af6a24d0a1bd11ddbae70e76c4a2342da9eb731f7d4dc4cbb0b9a1e8456cdba5ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h440dfcff61a859bafcfd9f74aa2427ebd691e2614e1fb68e407cb033523436430d51b337b75055b80d805e681d5bb46e0440;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab30c909e3c2924321e1d0851b1c4f70f158c7786fb82f75517861cbc353f100a354cea1366e55c5ede8ba9ba7fddaa360d9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63a7cf4ba2b1aa4159f8f379707f97534fc0eb1a64ccc8c7fee3ff8b457e6671371eb4c3c9378feaab6c7ece34ba51932d68;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h254e6e4ad44c861a21b0101f94ced547f3e9b07f3d52766d9b5dad67cd908e334b1756783f340404417035414df8fe0f1eb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd5948e7209d0d709ae8dc25e654b9196ae6675a054917a64052de362a7b0e9deb7533efef4481d9e2c6431bc8efc423e7fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h492c0d92a309f69e607953b30ae8bdcc0a7a6637aacb8db9fe90db50cd472e87e8f54152d427e600e2094cd6cddd599b6280;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e0826fffe69756c30a73cbda966ee17b8a21c957537f19a6aabf5c15ca56f8f754f887a0034e3a281f1d2d93e61151cae57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6eeb117796440484a7dcb8c9e16ffd354dc01ffe25b0b9aa7986a07da4870993b30f410177c9a9c807852d37305b5d0afac9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdd561e53c0ccd9e77c66ef206e5a6b1aa03525da061f9d59d8842f963a0b67c5ed4a01bf7fe4423773487ffcc26c3cff26b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha17c73bd2a8092f73e5fbeeb99d7f0dde89d07749ed9210d52e6bfc97408290c3762437adef8b92d22cdd272ea0ebd60304a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha87dd69c3e88a1e83f55be966cca34b24e80dad466716d2e65f1d32d977fda10acdb8e8ca855112ee6436b47130f3f7a010a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c1e2c3b3413e239cd4bf52ffc085527741bfe7b81fdeb3b8e862630c154c760899d3a51a2bfbe05bd7259efcf780670c5b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff3d92a77a6bcdf1096d6f1b695ebc0bee6ada8b2c00bf165580cc926ed8a0f62cf627f36ba0cfcf2c1fa7269c044c0affa3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bd4e5924737bcfaad3abd3f4cfbf2d23579802b378fa30553c89b495d83e3cb9ca898d3c748e0f71afd06c4724e96bc3fce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd13278a9b3ca81e63b539c1b5bfbd3d2165de0a203827a2d2a9c81689bbb09e2e8ca6fbeba9a21f5baf8fdaec87bbde6eefe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc39db4716e8f02aeb1d54d48625df1aa7716f6471ac8a32cb9a9a38a4806141dda5cc9bc51d234b393e18e1742b6c07aab14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dbae6d57e5ff41fc7d1adcaa58201635ad7acc7f26a28e4ee65ea7fe4906dfa400cc6501be6c6c26ea7f17b96d523726c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b10e8a387418a13eb5657a35f8b966b67ffc888ea6bd538a1507673b92d3acb9dcf3fc9903ba36f142fb625586b0ed99ae8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a04d9fcd6654b541af58a176ce48f1b4188973af6266b45421398cf4ccfc148311526f45c10c44543c783c3b72125765025;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6796b2dcef82a600b127f2b4c04290a0e0dfc5d3786a9cb6e670a224d19552f71731c99752a2d42d4cb8bb3516110d185528;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57ba0108c1518cbe1cd9a03fb1705f0bab99628bb257f61b6ec545916b3c740a4a50d7279f95cd4458b30e59aa599cd00615;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae23e569436ac2f4638d42277a73203c25475d921c11dddbd7f4363a1d0accaf8bd4d8f9eae1cd3e894ef5ac441ffb602ae2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaaffd47588b75104ff7a39fd85e5424a7b43728a96ad6a50c7584b292652c44f71adb5b9d4a547ba3727e0a09131c436563;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h681930ef6dd3979d500b9dbdce14177dccd64a744ea95df8ab31495d3ec1297773035422ab5f94a1ebb229d717070b1da3bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9de92cf90d2c4c037fe852378db87e54871002aa06d6b68a9cf0663b730cc421dda1fc25a37988163bec526c088f1989b8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8514a902e473a5683127487c7c39a0346ee4f4389361e4dc5bdbd8fe9fd48015bb887296624bc1c2a4113243e708ad2298b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf412d4811689889b78f5f42518cc7eb607e51343af94b07369a40c3f16aeeb760908f7826a54edaf0af5770ef254a9757f08;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf11768a7014215c33921b75ce84ff25f88e7664986a386a2cae9f4fb803f4b227ea2e1fcc355676092050c3e260b22c13778;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ba2eb70f10a60faf7fa8fb782428128dcbf67a8c807ce64e787c2f93a5759e21abf1dfc6d3bda789fbdc7e682582b84b1dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44ec5658c9c8f0b79f519c72880e7c0bece5902017bf5df79931aff66ff8d32f4b0d4818a671e33122dd2760cf3eaa6398e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f2d7c29846a1a09c7ed54c482b7e33d6cd58bba303b2d3fa9702c7d1f8cbab6ce0c9f3e5a65538576b675a016b7f4e6a15d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h60b068f22886f50846f1b144934738acac8cd6ad909b5d97c3c09ce6528455804f5574510598ce21966b774f3940703cbe9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc3105ebb8e158864a6eb251db0fc420fcc0bf09eb5e788b1e89f6fc1b144c09537efce04c4766b7474356cd52d9e97f74ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cc8384ec1cd61fedbd51d18cde651076fb74660469daafc9acadf81211db14206968ee3a8840497828d096995358810dd3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h371a4bb73037ce99af0994fd589b98dfb80c13176345010eb2ed8563a5274aa94b2b10c5f95e5c66a2f46d077b28933a168e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ca02f21c38dcb1d2258cd01ec3093af3b7caf346a8adcb267b0522b2fb88d9c04fa360f2180d06b7f4c745ba29d152b308e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h381323227dcf852fa3161809f2d23a29c64bf5113bb4d8a3e347007aecc1ee7f21240b09baa6f473b0013146fe3a5b337bc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he93a02f94ee086e9abf8d6345c044a5c60cc50c972cf39bc6197d296ff41f0cff4adb80d28807e3ff96e55fe62daeea822d9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76ec5d98b3f7f7e26cdcb35f99db1223a7f58e3b74d304d0257ee98d5b4316b23a2671ce902c8c571413824957d806e25a9d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfe5df05b468211aebc9ede570bf0f9ff3111c5b408b1a40741724f95c3e47d58470094b910aea2f80c6e263ae340d6dd3f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02b56084988dc36b6a7eae64f6a63f2683fa1289c321ac8d1de1b042c89b0be3a535d45a4d5e8afebc3df1b246e6eb9bdc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41e4af518dfaca009a7b2493f899a74aca9f2a8362a5fb142f80e031a5e1f99b1ae446dfe1eeac3b55dd2b503013a799c1cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f25a193372795a1a9c5726dc1b6c264fa89e99a7df6bf2b873d5135e59f0750a52b41e66f6d94faa9249622bb53ea360731;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9d705ccc069c3097b9d42572e5b3ce47fab0c5a71565bb9d348c78b1d167176ed24c86cb0f95cd19fb18e84a2fc8ea07e80;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ff60825bac60ca194660cdbf02948fcbaf5b604d18421d755d94a1afa2eeb749226508df3f2c7451d0388f2abb21441bccc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he909501b155bddc03c5de6004a0fbafc771e1c641f803871d22b9c4b6e15c142f032be3a1ac2715885771c431752ed44ea4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f27852890f6317809e2d9c12907dd5dcf8f33ebfa8e99bfe022124fc7f5ac348ee5f5cafbf2c1d9ba4314cb150678ca0740;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77b2e18ca30402badef27d776832c24ab44c3841a388730aa29e47f09a7fc47cffcb320ba0cd8403e1b673a7fed9a6726769;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h723bb94674712ae0f9527d68451058dca21e5cb3940083f3bc3590bed05db399a855bdf840c5467be296028db7692a2faf48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcda7c12bb933028a30b094340d143128e3982beda4b01a66d26eab7d944d561f1241161fc4f1f59a0c44d3f7a6afe875703f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he757ab03950f1a88bc6d290d3424703b4e62d08c90801c281bdde5f341a8ccda7e9bbf50c702b6e7649d06a4c0ad5e572b57;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3f7ffefc6950e85f4aa601c6ad5cea1004a14f5bc844470a14d2df42464b54385ae10968f8fc90124b9b79eb1df6185c682;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a9da8d4ce3ea76c6b4942387e8f57499a78af60e0fa84cf7c8ea9678f1b8e566716c36ac467d610befc02749b2fd7baf718;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa2c9e1507abbc084a314c49b812d70712488eb7f123ae15956725a72ed423ea168eef86071a7c6af56bc6303dc396c2ce1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf23ae1d028abe1e65e971ee6f6b5cd3212138a3bec71926ab6548e615059d82474a03e266bb9991eed773475de84142b035;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef56c96dd3d9c846a2f2ef99913b88cba54d89f5537dce0106bf73d8a37b35cd2af196b5d1bb6a178d6cd319b083482e5608;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he729551be7dd4b53bb1920bba96af6b72719ff53247d93ea3a3a3f232c8758b8396b4ec54f196433ee4343ebc22c0c38f9c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc997617f42397ddeafcc88e8b42501e41929832faa6039f924829f11b9bcc9ec3c6140d57dff7edd3b25dcf084a0aab40ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadaac4af76628d6c392b5b78569a0081a480bc4791eec86ad6d5831a78c46bf0c9b416e4979b29b444991e6f18b2e98fe20d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h358a4124bd7175015c5fba35b65703b2643003fd3b8b17ce5f13d557f0e56d8b12fbb5cb4c6d59da2b3de3f1c3cc5b6419a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47176184e05315433f505b4bce5bdd8a1eea29b570e75f3f838854a9b818d3c3ec4e49a3081e53ce195594720ddf505cf8f5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf99ab56c9cd4400f8be7cbe496bad9fe2fe4fd2427f404d83b106b08224d0ac5974cac6e547c62ae5799659f231e0a50155;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5ea4402cb30377fa46d40add9e0a76f2f8a7b515123c83022a6514f1da206b31b7d4bafa5e8478868d91420b15e971c9a1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74d1a216608173a7fe06c3884e2de875c0760c895782e2fd1bda36db9ee830dbe3030ef268c54677d9f60be59cc7a14705b3;
        #1
        $finish();
    end
endmodule
