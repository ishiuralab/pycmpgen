module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    compressor_CLA64_16 compressor_CLA64_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
        src12 <= 64'h0;
        src13 <= 64'h0;
        src14 <= 64'h0;
        src15 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA64_16(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    input [63:0]src12,
    input [63:0]src13,
    input [63:0]src14,
    input [63:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [0:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    wire [0:0] comp_out20;
    wire [0:0] comp_out21;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], 1'h0, comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      input wire [63:0] src12,
      input wire [63:0] src13,
      input wire [63:0] src14,
      input wire [63:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19,
      output wire [0:0] dst20,
      output wire [0:0] dst21);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [63:0] stage0_12;
   wire [63:0] stage0_13;
   wire [63:0] stage0_14;
   wire [63:0] stage0_15;
   wire [19:0] stage1_0;
   wire [29:0] stage1_1;
   wire [23:0] stage1_2;
   wire [26:0] stage1_3;
   wire [39:0] stage1_4;
   wire [28:0] stage1_5;
   wire [26:0] stage1_6;
   wire [22:0] stage1_7;
   wire [28:0] stage1_8;
   wire [29:0] stage1_9;
   wire [27:0] stage1_10;
   wire [23:0] stage1_11;
   wire [29:0] stage1_12;
   wire [32:0] stage1_13;
   wire [24:0] stage1_14;
   wire [23:0] stage1_15;
   wire [18:0] stage1_16;
   wire [9:0] stage1_17;
   wire [3:0] stage2_0;
   wire [21:0] stage2_1;
   wire [7:0] stage2_2;
   wire [10:0] stage2_3;
   wire [15:0] stage2_4;
   wire [17:0] stage2_5;
   wire [11:0] stage2_6;
   wire [11:0] stage2_7;
   wire [15:0] stage2_8;
   wire [7:0] stage2_9;
   wire [12:0] stage2_10;
   wire [17:0] stage2_11;
   wire [7:0] stage2_12;
   wire [18:0] stage2_13;
   wire [23:0] stage2_14;
   wire [7:0] stage2_15;
   wire [12:0] stage2_16;
   wire [5:0] stage2_17;
   wire [3:0] stage2_18;
   wire [1:0] stage2_19;
   wire [1:0] stage3_0;
   wire [6:0] stage3_1;
   wire [3:0] stage3_2;
   wire [6:0] stage3_3;
   wire [5:0] stage3_4;
   wire [9:0] stage3_5;
   wire [4:0] stage3_6;
   wire [3:0] stage3_7;
   wire [7:0] stage3_8;
   wire [6:0] stage3_9;
   wire [2:0] stage3_10;
   wire [6:0] stage3_11;
   wire [6:0] stage3_12;
   wire [4:0] stage3_13;
   wire [13:0] stage3_14;
   wire [6:0] stage3_15;
   wire [4:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [2:0] stage3_19;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [5:0] stage4_5;
   wire [2:0] stage4_6;
   wire [2:0] stage4_7;
   wire [3:0] stage4_8;
   wire [3:0] stage4_9;
   wire [3:0] stage4_10;
   wire [1:0] stage4_11;
   wire [2:0] stage4_12;
   wire [2:0] stage4_13;
   wire [8:0] stage4_14;
   wire [2:0] stage4_15;
   wire [2:0] stage4_16;
   wire [3:0] stage4_17;
   wire [1:0] stage4_18;
   wire [3:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [0:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [0:0] stage5_19;
   wire [0:0] stage5_20;
   wire [0:0] stage5_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[50]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc615_5 gpc18 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[51]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[9],stage1_4[18],stage1_3[18],stage1_2[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[3],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[4],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[5],stage1_5[13],stage1_4[22]}
   );
   gpc615_5 gpc23 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_5[6]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[6],stage1_5[14],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_5[7]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[7],stage1_5[15],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45]},
      {stage0_5[8]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[8],stage1_5[16],stage1_4[25]}
   );
   gpc615_5 gpc26 (
      {stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50]},
      {stage0_5[9]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[9],stage1_5[17],stage1_4[26]}
   );
   gpc606_5 gpc27 (
      {stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[12],stage1_5[20]}
   );
   gpc606_5 gpc30 (
      {stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[13],stage1_5[21]}
   );
   gpc606_5 gpc31 (
      {stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[14],stage1_5[22]}
   );
   gpc606_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[15],stage1_5[23]}
   );
   gpc606_5 gpc33 (
      {stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc34 (
      {stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[17],stage1_5[25]}
   );
   gpc615_5 gpc35 (
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_6[43]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[18],stage1_5[26]}
   );
   gpc615_5 gpc36 (
      {stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[19]}
   );
   gpc615_5 gpc37 (
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[17],stage1_7[18],stage1_6[20]}
   );
   gpc615_5 gpc38 (
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[18],stage1_7[19],stage1_6[21]}
   );
   gpc615_5 gpc39 (
      {stage0_7[57], stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61]},
      {stage0_8[18]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[12],stage1_8[19],stage1_7[20]}
   );
   gpc606_5 gpc40 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[4],stage1_9[13],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[5],stage1_9[14],stage1_8[21]}
   );
   gpc606_5 gpc42 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[6],stage1_9[15],stage1_8[22]}
   );
   gpc606_5 gpc43 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[7],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc44 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_9[6]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[8],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc45 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_9[7]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[9],stage1_9[18],stage1_8[25]}
   );
   gpc615_5 gpc46 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_9[8]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[10],stage1_9[19],stage1_8[26]}
   );
   gpc615_5 gpc47 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62]},
      {stage0_9[9]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[11],stage1_9[20],stage1_8[27]}
   );
   gpc606_5 gpc48 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc49 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc50 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc51 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc52 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc53 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[17],stage1_9[26]}
   );
   gpc606_5 gpc54 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[18],stage1_9[27]}
   );
   gpc606_5 gpc55 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[19],stage1_9[28]}
   );
   gpc606_5 gpc56 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[16],stage1_11[17],stage1_10[20],stage1_9[29]}
   );
   gpc606_5 gpc57 (
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[17],stage1_11[18],stage1_10[21]}
   );
   gpc615_5 gpc58 (
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58]},
      {stage0_11[54]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[18],stage1_11[19],stage1_10[22]}
   );
   gpc606_5 gpc59 (
      {stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[11],stage1_12[19],stage1_11[20]}
   );
   gpc606_5 gpc60 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[3],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc61 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[4],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc62 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[5],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc63 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[6],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc64 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[7],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc65 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[8],stage1_13[17],stage1_12[25]}
   );
   gpc615_5 gpc66 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52]},
      {stage0_13[6]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[9],stage1_13[18],stage1_12[26]}
   );
   gpc615_5 gpc67 (
      {stage0_12[53], stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57]},
      {stage0_13[7]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[10],stage1_13[19],stage1_12[27]}
   );
   gpc615_5 gpc68 (
      {stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61], stage0_12[62]},
      {stage0_13[8]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[11],stage1_13[20],stage1_12[28]}
   );
   gpc606_5 gpc69 (
      {stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[12],stage1_13[21]}
   );
   gpc606_5 gpc70 (
      {stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19], stage0_13[20]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[13],stage1_13[22]}
   );
   gpc606_5 gpc71 (
      {stage0_13[21], stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[14],stage1_13[23]}
   );
   gpc615_5 gpc72 (
      {stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31]},
      {stage0_14[54]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[15],stage1_13[24]}
   );
   gpc615_5 gpc73 (
      {stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35], stage0_13[36]},
      {stage0_14[55]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[16],stage1_13[25]}
   );
   gpc615_5 gpc74 (
      {stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_14[56]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[17],stage1_13[26]}
   );
   gpc615_5 gpc75 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46]},
      {stage0_14[57]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[18],stage1_13[27]}
   );
   gpc615_5 gpc76 (
      {stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51]},
      {stage0_14[58]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[19],stage1_13[28]}
   );
   gpc615_5 gpc77 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56]},
      {stage0_14[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[17],stage1_15[18],stage1_14[20],stage1_13[29]}
   );
   gpc615_5 gpc78 (
      {stage0_13[57], stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61]},
      {stage0_14[60]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[18],stage1_15[19],stage1_14[21],stage1_13[30]}
   );
   gpc1_1 gpc79 (
      {stage0_0[53]},
      {stage1_0[9]}
   );
   gpc1_1 gpc80 (
      {stage0_0[54]},
      {stage1_0[10]}
   );
   gpc1_1 gpc81 (
      {stage0_0[55]},
      {stage1_0[11]}
   );
   gpc1_1 gpc82 (
      {stage0_0[56]},
      {stage1_0[12]}
   );
   gpc1_1 gpc83 (
      {stage0_0[57]},
      {stage1_0[13]}
   );
   gpc1_1 gpc84 (
      {stage0_0[58]},
      {stage1_0[14]}
   );
   gpc1_1 gpc85 (
      {stage0_0[59]},
      {stage1_0[15]}
   );
   gpc1_1 gpc86 (
      {stage0_0[60]},
      {stage1_0[16]}
   );
   gpc1_1 gpc87 (
      {stage0_0[61]},
      {stage1_0[17]}
   );
   gpc1_1 gpc88 (
      {stage0_0[62]},
      {stage1_0[18]}
   );
   gpc1_1 gpc89 (
      {stage0_0[63]},
      {stage1_0[19]}
   );
   gpc1_1 gpc90 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc91 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc92 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc93 (
      {stage0_1[54]},
      {stage1_1[20]}
   );
   gpc1_1 gpc94 (
      {stage0_1[55]},
      {stage1_1[21]}
   );
   gpc1_1 gpc95 (
      {stage0_1[56]},
      {stage1_1[22]}
   );
   gpc1_1 gpc96 (
      {stage0_1[57]},
      {stage1_1[23]}
   );
   gpc1_1 gpc97 (
      {stage0_1[58]},
      {stage1_1[24]}
   );
   gpc1_1 gpc98 (
      {stage0_1[59]},
      {stage1_1[25]}
   );
   gpc1_1 gpc99 (
      {stage0_1[60]},
      {stage1_1[26]}
   );
   gpc1_1 gpc100 (
      {stage0_1[61]},
      {stage1_1[27]}
   );
   gpc1_1 gpc101 (
      {stage0_1[62]},
      {stage1_1[28]}
   );
   gpc1_1 gpc102 (
      {stage0_1[63]},
      {stage1_1[29]}
   );
   gpc1_1 gpc103 (
      {stage0_2[59]},
      {stage1_2[19]}
   );
   gpc1_1 gpc104 (
      {stage0_2[60]},
      {stage1_2[20]}
   );
   gpc1_1 gpc105 (
      {stage0_2[61]},
      {stage1_2[21]}
   );
   gpc1_1 gpc106 (
      {stage0_2[62]},
      {stage1_2[22]}
   );
   gpc1_1 gpc107 (
      {stage0_2[63]},
      {stage1_2[23]}
   );
   gpc1_1 gpc108 (
      {stage0_3[57]},
      {stage1_3[20]}
   );
   gpc1_1 gpc109 (
      {stage0_3[58]},
      {stage1_3[21]}
   );
   gpc1_1 gpc110 (
      {stage0_3[59]},
      {stage1_3[22]}
   );
   gpc1_1 gpc111 (
      {stage0_3[60]},
      {stage1_3[23]}
   );
   gpc1_1 gpc112 (
      {stage0_3[61]},
      {stage1_3[24]}
   );
   gpc1_1 gpc113 (
      {stage0_3[62]},
      {stage1_3[25]}
   );
   gpc1_1 gpc114 (
      {stage0_3[63]},
      {stage1_3[26]}
   );
   gpc1_1 gpc115 (
      {stage0_4[51]},
      {stage1_4[27]}
   );
   gpc1_1 gpc116 (
      {stage0_4[52]},
      {stage1_4[28]}
   );
   gpc1_1 gpc117 (
      {stage0_4[53]},
      {stage1_4[29]}
   );
   gpc1_1 gpc118 (
      {stage0_4[54]},
      {stage1_4[30]}
   );
   gpc1_1 gpc119 (
      {stage0_4[55]},
      {stage1_4[31]}
   );
   gpc1_1 gpc120 (
      {stage0_4[56]},
      {stage1_4[32]}
   );
   gpc1_1 gpc121 (
      {stage0_4[57]},
      {stage1_4[33]}
   );
   gpc1_1 gpc122 (
      {stage0_4[58]},
      {stage1_4[34]}
   );
   gpc1_1 gpc123 (
      {stage0_4[59]},
      {stage1_4[35]}
   );
   gpc1_1 gpc124 (
      {stage0_4[60]},
      {stage1_4[36]}
   );
   gpc1_1 gpc125 (
      {stage0_4[61]},
      {stage1_4[37]}
   );
   gpc1_1 gpc126 (
      {stage0_4[62]},
      {stage1_4[38]}
   );
   gpc1_1 gpc127 (
      {stage0_4[63]},
      {stage1_4[39]}
   );
   gpc1_1 gpc128 (
      {stage0_5[62]},
      {stage1_5[27]}
   );
   gpc1_1 gpc129 (
      {stage0_5[63]},
      {stage1_5[28]}
   );
   gpc1_1 gpc130 (
      {stage0_6[59]},
      {stage1_6[22]}
   );
   gpc1_1 gpc131 (
      {stage0_6[60]},
      {stage1_6[23]}
   );
   gpc1_1 gpc132 (
      {stage0_6[61]},
      {stage1_6[24]}
   );
   gpc1_1 gpc133 (
      {stage0_6[62]},
      {stage1_6[25]}
   );
   gpc1_1 gpc134 (
      {stage0_6[63]},
      {stage1_6[26]}
   );
   gpc1_1 gpc135 (
      {stage0_7[62]},
      {stage1_7[21]}
   );
   gpc1_1 gpc136 (
      {stage0_7[63]},
      {stage1_7[22]}
   );
   gpc1_1 gpc137 (
      {stage0_8[63]},
      {stage1_8[28]}
   );
   gpc1_1 gpc138 (
      {stage0_10[59]},
      {stage1_10[23]}
   );
   gpc1_1 gpc139 (
      {stage0_10[60]},
      {stage1_10[24]}
   );
   gpc1_1 gpc140 (
      {stage0_10[61]},
      {stage1_10[25]}
   );
   gpc1_1 gpc141 (
      {stage0_10[62]},
      {stage1_10[26]}
   );
   gpc1_1 gpc142 (
      {stage0_10[63]},
      {stage1_10[27]}
   );
   gpc1_1 gpc143 (
      {stage0_11[61]},
      {stage1_11[21]}
   );
   gpc1_1 gpc144 (
      {stage0_11[62]},
      {stage1_11[22]}
   );
   gpc1_1 gpc145 (
      {stage0_11[63]},
      {stage1_11[23]}
   );
   gpc1_1 gpc146 (
      {stage0_12[63]},
      {stage1_12[29]}
   );
   gpc1_1 gpc147 (
      {stage0_13[62]},
      {stage1_13[31]}
   );
   gpc1_1 gpc148 (
      {stage0_13[63]},
      {stage1_13[32]}
   );
   gpc1_1 gpc149 (
      {stage0_14[61]},
      {stage1_14[22]}
   );
   gpc1_1 gpc150 (
      {stage0_14[62]},
      {stage1_14[23]}
   );
   gpc1_1 gpc151 (
      {stage0_14[63]},
      {stage1_14[24]}
   );
   gpc1_1 gpc152 (
      {stage0_15[60]},
      {stage1_15[20]}
   );
   gpc1_1 gpc153 (
      {stage0_15[61]},
      {stage1_15[21]}
   );
   gpc1_1 gpc154 (
      {stage0_15[62]},
      {stage1_15[22]}
   );
   gpc1_1 gpc155 (
      {stage0_15[63]},
      {stage1_15[23]}
   );
   gpc2135_5 gpc156 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc157 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc158 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc159 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc160 (
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_3[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc161 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13]},
      {stage1_3[9]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc162 (
      {stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_3[10]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc163 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_3[11]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc615_5 gpc164 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[24]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[4],stage2_5[4],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc165 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[25]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[5],stage2_5[5],stage2_4[9],stage2_3[9]}
   );
   gpc615_5 gpc166 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[26]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[6],stage2_5[6],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc167 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31]},
      {stage1_5[18]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[7],stage2_5[7],stage2_4[11]}
   );
   gpc615_5 gpc168 (
      {stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36]},
      {stage1_5[19]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[8],stage2_5[8],stage2_4[12]}
   );
   gpc615_5 gpc169 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[0]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[5],stage2_6[9]}
   );
   gpc615_5 gpc170 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[1]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[6],stage2_6[10]}
   );
   gpc615_5 gpc171 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[2]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[4],stage2_7[7],stage2_6[11]}
   );
   gpc615_5 gpc172 (
      {stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7]},
      {stage1_8[18]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[3],stage2_9[3],stage2_8[5],stage2_7[8]}
   );
   gpc615_5 gpc173 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[19]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[4],stage2_9[4],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc174 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[20]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[5],stage2_9[5],stage2_8[7],stage2_7[10]}
   );
   gpc615_5 gpc175 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[21]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[6],stage2_9[6],stage2_8[8],stage2_7[11]}
   );
   gpc606_5 gpc176 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[4],stage2_10[7],stage2_9[7]}
   );
   gpc606_5 gpc177 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc178 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[2],stage2_12[2],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc179 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[3],stage2_12[3],stage2_11[7],stage2_10[10]}
   );
   gpc606_5 gpc180 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[4],stage2_12[4],stage2_11[8],stage2_10[11]}
   );
   gpc606_5 gpc181 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], 1'b0, 1'b0},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[5],stage2_12[5],stage2_11[9],stage2_10[12]}
   );
   gpc606_5 gpc182 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[6],stage2_12[6],stage2_11[10]}
   );
   gpc606_5 gpc183 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[7],stage2_12[7],stage2_11[11]}
   );
   gpc606_5 gpc184 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[2],stage2_14[7],stage2_13[8]}
   );
   gpc606_5 gpc185 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[3],stage2_14[8],stage2_13[9]}
   );
   gpc606_5 gpc186 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[4],stage2_14[9]}
   );
   gpc606_5 gpc187 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[5],stage2_14[10]}
   );
   gpc606_5 gpc188 (
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[6]}
   );
   gpc606_5 gpc189 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], 1'b0, 1'b0},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[7]}
   );
   gpc1_1 gpc190 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc191 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc192 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc193 (
      {stage1_1[15]},
      {stage2_1[7]}
   );
   gpc1_1 gpc194 (
      {stage1_1[16]},
      {stage2_1[8]}
   );
   gpc1_1 gpc195 (
      {stage1_1[17]},
      {stage2_1[9]}
   );
   gpc1_1 gpc196 (
      {stage1_1[18]},
      {stage2_1[10]}
   );
   gpc1_1 gpc197 (
      {stage1_1[19]},
      {stage2_1[11]}
   );
   gpc1_1 gpc198 (
      {stage1_1[20]},
      {stage2_1[12]}
   );
   gpc1_1 gpc199 (
      {stage1_1[21]},
      {stage2_1[13]}
   );
   gpc1_1 gpc200 (
      {stage1_1[22]},
      {stage2_1[14]}
   );
   gpc1_1 gpc201 (
      {stage1_1[23]},
      {stage2_1[15]}
   );
   gpc1_1 gpc202 (
      {stage1_1[24]},
      {stage2_1[16]}
   );
   gpc1_1 gpc203 (
      {stage1_1[25]},
      {stage2_1[17]}
   );
   gpc1_1 gpc204 (
      {stage1_1[26]},
      {stage2_1[18]}
   );
   gpc1_1 gpc205 (
      {stage1_1[27]},
      {stage2_1[19]}
   );
   gpc1_1 gpc206 (
      {stage1_1[28]},
      {stage2_1[20]}
   );
   gpc1_1 gpc207 (
      {stage1_1[29]},
      {stage2_1[21]}
   );
   gpc1_1 gpc208 (
      {stage1_4[37]},
      {stage2_4[13]}
   );
   gpc1_1 gpc209 (
      {stage1_4[38]},
      {stage2_4[14]}
   );
   gpc1_1 gpc210 (
      {stage1_4[39]},
      {stage2_4[15]}
   );
   gpc1_1 gpc211 (
      {stage1_5[20]},
      {stage2_5[9]}
   );
   gpc1_1 gpc212 (
      {stage1_5[21]},
      {stage2_5[10]}
   );
   gpc1_1 gpc213 (
      {stage1_5[22]},
      {stage2_5[11]}
   );
   gpc1_1 gpc214 (
      {stage1_5[23]},
      {stage2_5[12]}
   );
   gpc1_1 gpc215 (
      {stage1_5[24]},
      {stage2_5[13]}
   );
   gpc1_1 gpc216 (
      {stage1_5[25]},
      {stage2_5[14]}
   );
   gpc1_1 gpc217 (
      {stage1_5[26]},
      {stage2_5[15]}
   );
   gpc1_1 gpc218 (
      {stage1_5[27]},
      {stage2_5[16]}
   );
   gpc1_1 gpc219 (
      {stage1_5[28]},
      {stage2_5[17]}
   );
   gpc1_1 gpc220 (
      {stage1_8[22]},
      {stage2_8[9]}
   );
   gpc1_1 gpc221 (
      {stage1_8[23]},
      {stage2_8[10]}
   );
   gpc1_1 gpc222 (
      {stage1_8[24]},
      {stage2_8[11]}
   );
   gpc1_1 gpc223 (
      {stage1_8[25]},
      {stage2_8[12]}
   );
   gpc1_1 gpc224 (
      {stage1_8[26]},
      {stage2_8[13]}
   );
   gpc1_1 gpc225 (
      {stage1_8[27]},
      {stage2_8[14]}
   );
   gpc1_1 gpc226 (
      {stage1_8[28]},
      {stage2_8[15]}
   );
   gpc1_1 gpc227 (
      {stage1_11[18]},
      {stage2_11[12]}
   );
   gpc1_1 gpc228 (
      {stage1_11[19]},
      {stage2_11[13]}
   );
   gpc1_1 gpc229 (
      {stage1_11[20]},
      {stage2_11[14]}
   );
   gpc1_1 gpc230 (
      {stage1_11[21]},
      {stage2_11[15]}
   );
   gpc1_1 gpc231 (
      {stage1_11[22]},
      {stage2_11[16]}
   );
   gpc1_1 gpc232 (
      {stage1_11[23]},
      {stage2_11[17]}
   );
   gpc1_1 gpc233 (
      {stage1_13[24]},
      {stage2_13[10]}
   );
   gpc1_1 gpc234 (
      {stage1_13[25]},
      {stage2_13[11]}
   );
   gpc1_1 gpc235 (
      {stage1_13[26]},
      {stage2_13[12]}
   );
   gpc1_1 gpc236 (
      {stage1_13[27]},
      {stage2_13[13]}
   );
   gpc1_1 gpc237 (
      {stage1_13[28]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[29]},
      {stage2_13[15]}
   );
   gpc1_1 gpc239 (
      {stage1_13[30]},
      {stage2_13[16]}
   );
   gpc1_1 gpc240 (
      {stage1_13[31]},
      {stage2_13[17]}
   );
   gpc1_1 gpc241 (
      {stage1_13[32]},
      {stage2_13[18]}
   );
   gpc1_1 gpc242 (
      {stage1_14[12]},
      {stage2_14[11]}
   );
   gpc1_1 gpc243 (
      {stage1_14[13]},
      {stage2_14[12]}
   );
   gpc1_1 gpc244 (
      {stage1_14[14]},
      {stage2_14[13]}
   );
   gpc1_1 gpc245 (
      {stage1_14[15]},
      {stage2_14[14]}
   );
   gpc1_1 gpc246 (
      {stage1_14[16]},
      {stage2_14[15]}
   );
   gpc1_1 gpc247 (
      {stage1_14[17]},
      {stage2_14[16]}
   );
   gpc1_1 gpc248 (
      {stage1_14[18]},
      {stage2_14[17]}
   );
   gpc1_1 gpc249 (
      {stage1_14[19]},
      {stage2_14[18]}
   );
   gpc1_1 gpc250 (
      {stage1_14[20]},
      {stage2_14[19]}
   );
   gpc1_1 gpc251 (
      {stage1_14[21]},
      {stage2_14[20]}
   );
   gpc1_1 gpc252 (
      {stage1_14[22]},
      {stage2_14[21]}
   );
   gpc1_1 gpc253 (
      {stage1_14[23]},
      {stage2_14[22]}
   );
   gpc1_1 gpc254 (
      {stage1_14[24]},
      {stage2_14[23]}
   );
   gpc1_1 gpc255 (
      {stage1_16[12]},
      {stage2_16[6]}
   );
   gpc1_1 gpc256 (
      {stage1_16[13]},
      {stage2_16[7]}
   );
   gpc1_1 gpc257 (
      {stage1_16[14]},
      {stage2_16[8]}
   );
   gpc1_1 gpc258 (
      {stage1_16[15]},
      {stage2_16[9]}
   );
   gpc1_1 gpc259 (
      {stage1_16[16]},
      {stage2_16[10]}
   );
   gpc1_1 gpc260 (
      {stage1_16[17]},
      {stage2_16[11]}
   );
   gpc1_1 gpc261 (
      {stage1_16[18]},
      {stage2_16[12]}
   );
   gpc1163_5 gpc262 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc263 (
      {stage2_0[3], 1'b0, 1'b0},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc264 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc265 (
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc266 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10]},
      {stage2_5[0]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[4]}
   );
   gpc615_5 gpc267 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15]},
      {stage2_5[1]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[5]}
   );
   gpc606_5 gpc268 (
      {stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[2],stage3_7[2],stage3_6[3],stage3_5[4]}
   );
   gpc606_5 gpc269 (
      {stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12], stage2_5[13]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[3],stage3_7[3],stage3_6[4],stage3_5[5]}
   );
   gpc1163_5 gpc270 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage2_10[0]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[2],stage3_8[4]}
   );
   gpc606_5 gpc271 (
      {stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7], stage2_8[8]},
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[3],stage3_8[5]}
   );
   gpc606_5 gpc272 (
      {stage2_8[9], stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14]},
      {stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[4],stage3_8[6]}
   );
   gpc606_5 gpc273 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[3],stage3_11[3]}
   );
   gpc615_5 gpc274 (
      {stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[4],stage3_11[4]}
   );
   gpc615_5 gpc275 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[1]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[5],stage3_11[5]}
   );
   gpc606_5 gpc276 (
      {stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[3],stage3_13[3],stage3_12[6]}
   );
   gpc615_5 gpc277 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[4],stage3_14[4]}
   );
   gpc615_5 gpc278 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[5],stage3_14[5]}
   );
   gpc606_5 gpc279 (
      {stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[6]}
   );
   gpc1_1 gpc280 (
      {stage2_1[18]},
      {stage3_1[3]}
   );
   gpc1_1 gpc281 (
      {stage2_1[19]},
      {stage3_1[4]}
   );
   gpc1_1 gpc282 (
      {stage2_1[20]},
      {stage3_1[5]}
   );
   gpc1_1 gpc283 (
      {stage2_1[21]},
      {stage3_1[6]}
   );
   gpc1_1 gpc284 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc285 (
      {stage2_3[9]},
      {stage3_3[5]}
   );
   gpc1_1 gpc286 (
      {stage2_3[10]},
      {stage3_3[6]}
   );
   gpc1_1 gpc287 (
      {stage2_5[14]},
      {stage3_5[6]}
   );
   gpc1_1 gpc288 (
      {stage2_5[15]},
      {stage3_5[7]}
   );
   gpc1_1 gpc289 (
      {stage2_5[16]},
      {stage3_5[8]}
   );
   gpc1_1 gpc290 (
      {stage2_5[17]},
      {stage3_5[9]}
   );
   gpc1_1 gpc291 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc292 (
      {stage2_9[6]},
      {stage3_9[5]}
   );
   gpc1_1 gpc293 (
      {stage2_9[7]},
      {stage3_9[6]}
   );
   gpc1_1 gpc294 (
      {stage2_11[17]},
      {stage3_11[6]}
   );
   gpc1_1 gpc295 (
      {stage2_13[18]},
      {stage3_13[4]}
   );
   gpc1_1 gpc296 (
      {stage2_14[16]},
      {stage3_14[6]}
   );
   gpc1_1 gpc297 (
      {stage2_14[17]},
      {stage3_14[7]}
   );
   gpc1_1 gpc298 (
      {stage2_14[18]},
      {stage3_14[8]}
   );
   gpc1_1 gpc299 (
      {stage2_14[19]},
      {stage3_14[9]}
   );
   gpc1_1 gpc300 (
      {stage2_14[20]},
      {stage3_14[10]}
   );
   gpc1_1 gpc301 (
      {stage2_14[21]},
      {stage3_14[11]}
   );
   gpc1_1 gpc302 (
      {stage2_14[22]},
      {stage3_14[12]}
   );
   gpc1_1 gpc303 (
      {stage2_14[23]},
      {stage3_14[13]}
   );
   gpc1_1 gpc304 (
      {stage2_16[12]},
      {stage3_16[4]}
   );
   gpc1_1 gpc305 (
      {stage2_18[0]},
      {stage3_18[3]}
   );
   gpc1_1 gpc306 (
      {stage2_18[1]},
      {stage3_18[4]}
   );
   gpc1_1 gpc307 (
      {stage2_18[2]},
      {stage3_18[5]}
   );
   gpc1_1 gpc308 (
      {stage2_18[3]},
      {stage3_18[6]}
   );
   gpc1_1 gpc309 (
      {stage2_19[0]},
      {stage3_19[1]}
   );
   gpc1_1 gpc310 (
      {stage2_19[1]},
      {stage3_19[2]}
   );
   gpc606_5 gpc311 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc312 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], 1'b0},
      {stage3_3[6]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc207_4 gpc313 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[2]}
   );
   gpc615_5 gpc314 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[2]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[2]}
   );
   gpc615_5 gpc315 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc606_5 gpc316 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1]}
   );
   gpc615_5 gpc317 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4]},
      {stage3_14[6]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[1],stage4_13[2]}
   );
   gpc615_5 gpc318 (
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[2]}
   );
   gpc1_1 gpc319 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc320 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc321 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc322 (
      {stage3_5[7]},
      {stage4_5[3]}
   );
   gpc1_1 gpc323 (
      {stage3_5[8]},
      {stage4_5[4]}
   );
   gpc1_1 gpc324 (
      {stage3_5[9]},
      {stage4_5[5]}
   );
   gpc1_1 gpc325 (
      {stage3_7[3]},
      {stage4_7[2]}
   );
   gpc1_1 gpc326 (
      {stage3_8[6]},
      {stage4_8[2]}
   );
   gpc1_1 gpc327 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc328 (
      {stage3_9[5]},
      {stage4_9[2]}
   );
   gpc1_1 gpc329 (
      {stage3_9[6]},
      {stage4_9[3]}
   );
   gpc1_1 gpc330 (
      {stage3_10[1]},
      {stage4_10[2]}
   );
   gpc1_1 gpc331 (
      {stage3_10[2]},
      {stage4_10[3]}
   );
   gpc1_1 gpc332 (
      {stage3_11[6]},
      {stage4_11[1]}
   );
   gpc1_1 gpc333 (
      {stage3_12[6]},
      {stage4_12[2]}
   );
   gpc1_1 gpc334 (
      {stage3_14[7]},
      {stage4_14[2]}
   );
   gpc1_1 gpc335 (
      {stage3_14[8]},
      {stage4_14[3]}
   );
   gpc1_1 gpc336 (
      {stage3_14[9]},
      {stage4_14[4]}
   );
   gpc1_1 gpc337 (
      {stage3_14[10]},
      {stage4_14[5]}
   );
   gpc1_1 gpc338 (
      {stage3_14[11]},
      {stage4_14[6]}
   );
   gpc1_1 gpc339 (
      {stage3_14[12]},
      {stage4_14[7]}
   );
   gpc1_1 gpc340 (
      {stage3_14[13]},
      {stage4_14[8]}
   );
   gpc1_1 gpc341 (
      {stage3_15[6]},
      {stage4_15[2]}
   );
   gpc1_1 gpc342 (
      {stage3_17[1]},
      {stage4_17[2]}
   );
   gpc1_1 gpc343 (
      {stage3_17[2]},
      {stage4_17[3]}
   );
   gpc1_1 gpc344 (
      {stage3_18[6]},
      {stage4_18[1]}
   );
   gpc1_1 gpc345 (
      {stage3_19[0]},
      {stage4_19[1]}
   );
   gpc1_1 gpc346 (
      {stage3_19[1]},
      {stage4_19[2]}
   );
   gpc1_1 gpc347 (
      {stage3_19[2]},
      {stage4_19[3]}
   );
   gpc1325_5 gpc348 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4]},
      {stage4_6[0], stage4_6[1]},
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0]}
   );
   gpc1343_5 gpc349 (
      {stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc623_5 gpc350 (
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0],stage5_12[1]}
   );
   gpc1343_5 gpc351 (
      {stage4_14[6], stage4_14[7], stage4_14[8]},
      {stage4_15[0], stage4_15[1], stage4_15[2], 1'b0},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc1423_5 gpc352 (
      {stage4_17[1], stage4_17[2], stage4_17[3]},
      {stage4_18[0], stage4_18[1]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3]},
      {stage4_20[0]},
      {stage5_21[0],stage5_20[0],stage5_19[0],stage5_18[1],stage5_17[1]}
   );
   gpc1_1 gpc353 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc354 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc355 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc356 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc357 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc358 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc359 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc360 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc361 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc362 (
      {stage4_4[1]},
      {stage5_4[1]}
   );
   gpc1_1 gpc363 (
      {stage4_5[5]},
      {stage5_5[1]}
   );
   gpc1_1 gpc364 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc365 (
      {stage4_10[3]},
      {stage5_10[1]}
   );
   gpc1_1 gpc366 (
      {stage4_11[1]},
      {stage5_11[1]}
   );
   gpc1_1 gpc367 (
      {stage4_13[2]},
      {stage5_13[1]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    reg [63:0] src12;
    reg [63:0] src13;
    reg [63:0] src14;
    reg [63:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor_CLA64_16 compressor_CLA64_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80d751dd93924eb1cf1528062f669c0497adfd4daa1773fac519515781fa1d56aa1652de38d93d9aaf4bb4036340aa9e024415fa0bc9ab3a8dd9f4a6b7e2588238030e6d1d5c1385958ebe27f4febc6614c68c58738b86ad8df302be65c4e2548a5b04049340cc2a3cf3d5e410af9fae2d4ac9cf53faa657a49148f548359a7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53b3f8f40a54fd834f8aa2fa0f3d0d3585dc7a0075bc37411bae356e5ad8075fb3e525f7c2195768613a50677a7a068d00eddcb37d060e04a92a4057a527b8a7da3a83b1bcf838dafe76c861705b53e67f272e0a2f2971a8e17671fe732ea5c5e69606dd5035ce5385cde6f444fcafb533fb53bfa10426ee7ca966eeae6c3090;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20db2d2f4841c93cf509413ec1194e983abb569345d16d517a2e6602c5b6a067a2030ca0a6ce1682fdb5632e5bc85cf927cc59b042822f7a5567e69d066cf1b1441bdca4ae9803bae1cfcee36cf8e63838797803739d3dc946e0722d4bcf07c154c73028e654eabb10c3555e643e8dacb4c6e0863ed115b01a8ff7f1b59f59a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea68cdee693d2269d4a4065a900e7d35c4610bee50b6f7ddeb006283eaeae793bea043280f66d9b1c5428887a6edba67249f50bf77d2c82f89d090069a4c4ecef2ffc61617c2344e0c365a2caa40eabd13eccc62b831659129ad7dd14167f396c405147df2b0e6e775ca5a64f65d2c832de5b9bf55c75b45383163c8fad83bb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3425330f7e9931dc331dd9452368fddd07e6238698de2cd9ab880978403141ac86e3b0c382213d9549e7fc0c9518f5b8c81fc831b3aea7e5fcda8d66ff1614f53f99046581c55d0408876c0a2a35ebf2a98e92d8095b636292a73013cd8f337f3cf738ac2cfcf46208bfb99d7acae1d16b00465a0277a3347884718104175904;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56fba216406c6a7c32271b389c1f23ab5905438bfb6cb6c7d76024b4292aa5e5df19874a80911539170ca2e2ee1c25b9bc4eb63ef056afcbfefc2e68613d62a6c5bc815618d2c297f9b4c29c21caa57d92464ecaded2d8dc8918a7c044ebb452e750d569886cb946c85e6b62c39e20d1805a4d64d2a718ce370e733e93e6d9fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1d907240fd54046822ff0ac9637175b047430e9e39dcc1f4596aab78d383051bb2b287bb2e3eb9e2251bbfb4fa2d2847ffa65f2db8ad85cd944387528c7d650604ad8f79f82d1e9a2bb138f93ee5b7f11803d29a4f1a1205ed00b2786fae9d56f3a559f06bed6d2df727a03b13a7f48e0a5e95b20e344e18aa8ed3171acd7c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe6fae3fdcb3df5594183615269cf5cbcd3b2df561490c3f283da769f81e57551136c3b99ff0b394681cf122d3639550817a02f0551f4c435b9b85bf0e0abda551536b30419e212821d31345621f3e344b54397454b3c1f3dccab2437cf5901266545cad314276312dfd7ca55f8956fc2965a648323deb09bb348d18ff2ecb86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4aaad3a0017f2aa205bac00a2c1522001edf2998b21bdc6a97b11f048b9c28ab9c4ebed2b7581609b5657a6baaa4655545df836ed2622e94c7b043ecfc71bce2abf5698bdc9b6ace61590a462d11116c0b8148b1044bf5e06943618ba18ed0e638a256be6ff928b32102661266041539f3a718dae1b882e37a4d63f720c279e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca45e13f7262367c2a3fb3d24f2437bbd99bab32c81789c0f68744519e8ce12293134570d9497d868c9f7a221a0dffc0f2d8a0d8c945336a6e2cc477127274729d7397bc31ee635d21d76d82db0e597acb854d1f21607fdfd90b351bb53d589cc75b20333f165d1d36f9f255e010630374156b223e9bc2b193f412fcc371d031;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9860905e863244c9300879c8e0c34c64f60b5976559d57c49ecee42012e3274f89af8163c6a6705e54bd8417e16ec3fb1a106c8f0d9c8b56a4864e9b3d9b39a92c958be70b4a934d531612930526254660ad949fd2eda71d930feef9fc7d42bea76f9d19f34a31f173f0fbf8f419e0d2dcbb781ef204131b5bc191b3c0fe4c5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc01518f414d699d1f792de99d7aad96d09814680612508ca64929745b81f7106f0f2b2b19839666d8615ab7307890ac2cc70b8a0f90d50caf23d7abc8bd247b15fde31b8cb22a7a9418025c7644adac062870c3ac7d7fb9cadfb30823fae897adab8c4d7b68b2f28e356dc64cb0e71790b3df855566321a6410d8df8801f01d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h871fe2aedafa4455f005da9a945d79ee14ea8abac40d3de5d08b1f1e68d9a65879e7acdb94bb5dab6bc50636c23e9bf575d9c2ad1bf0726322dfbb7b5f7ca0731eaebda06d2fcfb55c911bb01d11b32de28061210245f4e06a3af17793047f970f343821c3286f9dab5b601dc7369a70cd4056f952de75bf493c0330dabed0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf652a67b622367274d786e1054dc977c535edddebf02d5fbb2bb9b6b13b470bb8c6dd3ca0ef932c695597a2759cfe6a1d7b3ece9582cb189125ccfdcc59e5a0ecc792a9334ac12ba6fc459459b428076dba21379337094f5f835840e876540829429d7e4a1763c9602972485501e7e4a8bea8bb2ed5807d14619587db6ac23ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61755c2096ac79e2d3a8fc3a5a56295cabf69e135b5603590cac55d08b7b4451be0cebd2350d8033233474e01b79019d466567e316dbe5f98c14c726caecb9b898a2ddc8f6d90f8ca97c5cf187b8d9630929a6e49b8e4a2a90cd7f9d6f6374db5a553595e2dbea429d34053814fcfa5ce57cf140b7d60435e2fed956588dc62a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc36d7b842fae114e97a873e9fb3ee097197f92fabfd8126a8b6838cc551d9d52c326d54e993e2da277cce820bf6de2b727dd8c36cdd78ff92f46cc3a6678b72c7664d0d1dcaee565dca925e3731ea3f89fbc495995c0a5c87beac7169d961316a5c0f2917c43ec78ac9de25119f733d4e2512e3462efa8784e3c0a16d2268634;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b46e9941ea66f12e9d597e040bf2e5287d7c8ee88225b1f2d3cbf736b22907a9a86745389669e211b5b1b5c12069b21eb91c2a854bb356b32e86ef8eaebdd7ec04778916bee4d0c8309248a5508b123c58769dfc7cd01901433242bc7ea634340c1c24ae81594fc9ec59cee294d50268822ecc5c36ad546211765e15b85f20c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe1453a0967db96f1419ea7ffbef0110584a079972bb070f730c54d433dce4aedf954bc5c67d7658f7d89b8e3f71a73f719cb8f53f6348b62d70cd29716d9aeeffd280bd3d02ccf64368039bd06cd3b4f572962e50cc50f451c50f3ae162a9796d5bbdb516cdc7cfae119276c07feb515fc190aaccc529dc1cb9187c462f3182;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda15ab45ee7424f8f5417e660d18e440fe37604f35f47de847a1d1ef3a0790d168daf28af8bb2fbd766110571871d51f01262786834e55286d18b95b71fb344ec7819078a0e48e41f093989785b05882351f7abcbceffcae6c415875741fcc38cd04f652829a9316290e7332d3bf2e220072bd7c898bd28fc4951d9f6eeec25a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf25c043975e3f194371db4a9449c952d0dc3f4c0b9d79cae7b6b3e1e67abac402325edc823a377c8f01356559a3ece9d8728326c611fc2d82e88e56043f064ddd3c0728bdac1dbddba7432e9425bef519d2441e0d14acf5da43d99015a157ec11e0b0a7ca602d43bd7c638e0ec3f0438a1bd664cf98a6cf550602c3414164858;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4ba7f36983febdcc1fdab804dcf260f315b146ff8af109f3a04423278f5196a4ce5150b21bcdc2bf3e6742d94e72812563f3b85742b387c152361b8e77cf3edbd85f5d0f7e61a16a311b7e2f32ff4913e1bfcd0158d7621e2f7a32409694bffa5073ec110874f07c6b1db647993aa0a04726b2f3cb4a20115a7e9a3c064a4f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53460d704f127211be916cde06b4d6467481f5c9b76989ec584395338024f0fb1d624d5c0458ecb4bcd93b24ee4ae64dc89c99960a475d9f61b4adffa0218fec8ea45d9e8a962dffe8fd34163cfeac034423ccb3c291919f0913537c0ff6d090ba5afcdfa934da0ca204210effc20e4d02bd19bc72a757b478bbf8132faaaabe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ec4f2b6599ad1529564af989bb746043e187cb7dd9c569ba5f24b3c2b265a650251280b7ad446246c8312cf00610b0d61a3b925077d8950cdaac58b5a2662667139ec3da3b77b686610f4bd346c70169af6b4f8e78571f27b8f6c5ea260db3eb33ff914f125dc1e2f50b1939cf11217c8db1398b14d52604e4418bbc03c3536;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h484553557bedcfbce817fee93c5a58ee66e82dd795d29df738cbfa6b16bb53da66d1850a00139ad57f53f3ae01fbb1ba7a2de40480e766d155177dee7f9f48c7f8a44cad17805c06fa66a11954a6640ad6c41767c920c51efb536fbf1902b46bce9c45b5dc16b3e47e572805b699bd57aa06f85da059eeac301c4773e901e352;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc04c31b99a7202d837d6be6353b5068f566aa82e37ad3ec0696bcffd9002353a5fdb3bfaab5ad241894846ab42768f75fa239328d5b00f98aab4d29810580072702905632e83f425a4a2b7ef9c7d3e904bae9e49f75eb2dd782912bb69b656e9205616809b126df84eb4490e914c370ce578396768647d864f7d81565970dfcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b18404a2b914ff07e19a399fa9ede2974c6eed4a1a8028acb812bab7e77dd0aec820d15e44a01a5fb490b8c4b612badbe61c7b729c910df7b432c33bdf003b9bccfb611d12ec8efe811380d5ddae17b7b27bfb3112af4bd6c9464382447cb25bfd23c6e533bfc2ce5d067d36ab6195e66b4ec82eabec48dafdaec97bac75ea9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37d1b82444d2b62c804f03208e517fabcb4464c7c252c6e2503d5b1fa647b95c55babc4f21b2a0365502e0d230eccf6aef9ec40062c3a50ba90c5c4c9d015a35652840454e107a124b822431febb73dd8b60aaf1d353b42027caef92ba56b0e81d9b2c8944a0009416747cda990bb4b90666697363dab560da09a16bbf550303;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6276dc8d2ed8f705ba9127686c011351b86b53828b4222ed8cca5b74d383c596e976d21aa86420e1759fd9c9a168a6d4604ea13a532ee70908e8560055b26f5626beb4f80df71178635b41ab0e1a0db9b2b5b0ce8d0041ec48947ad7d4f26beea3fe375133538eee2db405f59290aaef459993254a25075d0dc177b98faf72c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadea346e14e67885f32278600d57d29cd87481de18fb3e42363665f7681dd10dd264cf047d55bd15abcfef1ff8dcb96405d4684522a7695e2b6de1d83efcda3debccd9359cc598cede7d44c37387a532b60b08d86e2d64a91a1026550b6f3ce5f4cd6c99e812c8fde5a1e19d58d567ce957d59c93ce59fa26344b7ca586f4f77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd215c84f4964eaf332d76d972a9da8ae4107585d78d649b16f5606875429d22e9042032bd0c36df6ea59a526860e23a76b22bf48389abfb9bbc95620e385e2566df16a678b1ed1dbd445c991a6757bc7266cc35941c75905cd2f0254265ddc861c447e8bcfa4b62b6ac5edc2d25b2a7f1b15e26652aeb1bf97bf61e0d030ab04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a6a312725bda3afca591664066f1aff894a02131c195fbd1559d3c5638c977ea5b002e672c327c5b048c06566b52be084571da76bb7ba183ba2c57d606728f18d4bf3326637fda162b59dc6b3f95df40f01d2da2c7cd72a67c105c10cfe584b0e86bdb5072b8886441f224465de79eb2d49cf9f33baaf3452f8ca08f50563ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fd0847a804d2c19bdec14b96bb73256dc0bb7d7def28292b26c01ff44f733c7dd9f5d5ae63f7b4886b507cda96b3a8994595fe01ed248208b25f8a1c16b1800b37fd3440c6ce292e07277d809d49de690e92b5201bbbd3ede2a01e2a5eadcefa9c6b2bd1ecf100d4a61b37555a2c7458b15a8b59d17f1dcaca632b1b76b58ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b3440066132acc5f8d7ed545ae9d21e65bf9b269c17c2671275db7eadf81ee73e91db986476e514a0bb05a30a2789446c407b69e162a3f0838be5e98a87b437d6a8b2438f26ba94ef8deaf6196f3008b0a52e52a694426a6992ae18711d4b8d991421bce2aab0e47af8887fd0ebc57eae148accbd2f9e8331347bbd8c8371a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9275a0f504d8d80b6476fe530bbf7ef029d4ef8b676095e3cfb0285a9a32eef68026e0349d3a7063d1a0483e4de39922bb7e86baf170cd45d12d595d4e877b79764f23e2c5e20d44a6c8c96da53fc4044dd91ecf741bb6cec1eebd8c5638b9658f35b41d5b5201229289130ee288a35e5ead0f645132f5d299974eebe1c8776d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85de3ce73c0eaa1bdc0e3a48f3c96ff8e4f5e8daa9c20f215f592a180af03cec3479bece7305ab0fb507a07c49799272b6d03d26b17a6c961460eac2c7308303bd5b24126366f97ba22bfb4e08001fbcbd1cdba650eb503720b14621d0cd453412434ab19ec23f7ec1ebb1d72b40e8a15fe902df53f2e16018c6e2acb746bd10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfa7d3d387e9470f7ca37fc4a2f47175ee0f52358eb6854fa79a150c156ec227d78a4ed1da66d78a1adc8acc4fbb3033673d03e5e4290deb47ee7213c4bb7e3a7a85b4cd6dd6d0d2ecce8491c5785ee2a7b3934dc9d91fa5d26dd1fae98a83f3b3a9ea77e037c27311eabd32ca8db27051458e40205a61137273f8c7282b0ee0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd4f88e6cc5e9bafded9904985359a4817c0253fce774d0e9897e80156a18d7b400f9f530ace9ac3f5d23db39fc3a0311758ff4101acae99862c19750113a319a553b23fec12a8b8b09a059a8ff3ef72c6d7e5455d0e5e8887c76a820c06b64dc5c1c8e976856deeba06101028e2310d65553287ac15246fcf8db1421090a1ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65cabb984d972d08dc81e06f8c048bc344747a18cfe2dbcef7a91d1744022ec8a71f11f19bd1390126f965bbe1cf30a5f0bd5f5180c960e3e1d51611c251b5ebccd586ddafda6781bab5739314364681059c86c3d3bdf857ffae5e0c41abe9170b27a068fe48263ccbd6ccc1035e0769b6f338a635220c9c72e3004e1c12b7d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1700e7d6bb479cc287e36bf404bb27c9125028ee87ab3be98d3c6430011a82692d8c15ba42802bc800340614b264927768689e094c1ec2aa09dd40d10a02f23b153f727eee0d8f1b76942307ebf6652d9f02218f26ce9db8532740280cdbe5e63cecc832b3e9f6e6d15973945ab98a24176da6d587796e5564af3dfd951bcc31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e36f99239e57f10520a36f322badd9b30a455523a5a6c80a6b4c6ca05990990a1c60c2e28e94eb23b3f9007924d6e5259e86f3dcef8db9098360cb12be608ce933b3ed264b774907bf5ffcc209fa47dbe220c33b85a234f2bf818c8068d84a77197df7c81a07511e0aef29039e54962040864b696b755dd4db9710e4d43e58f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae2b8f960722a1a569a8c807f901723634ccb15c32f857833908faed8ac63ca9991e20181766e703bd1f40e630a7d6d318363bf39aeef98bd466d9ce3413d0266050812b5c493f753995d5b47b8c1670232744df104bbc181370350daa9ea6b312910c1905b883a34409cafb3b06915a2f10d7a2330557296ec221446528739a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1143a8203f793c821f549698f681515ae904506b73d961f3f31e0424bfcba982259c217e90014449c6667f906031455c7b4980ed0233316002a046a6c0897010a04f8c6aa3adb5fd18f40abcdc3568ce95e2d43ad0815935309b46aa4b08062bec90037bdf8a19600c1201d3ee26063f8398ec26dae2f9a904b13fa597611a21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h862f2c564890e2f50dfb5d222fad5cc548abf7b8a1d25a0838e46298c27cf29920c62edba4dab7b093fcb60e872fb784b1d7cc71822192f560a147dded5460a2be68b8c38f4737393295cc377af1ce03925afbfeb2c3a080ac0d78368c8a19fb1d91d718b58ff5cbb55dd0f4b2bb3f0f71fb2c25dbd8c9ea3383a56c5a8eb989;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2571132456cca8b4c381d6982e9db3b1cb2932e450a8b1e2a76f20bf648167f96f5c33cf590dd514d5b2c0cad3c5f13a9b50d508abf593e42b2e7404a22a33da1b73311730c363b2c6717f8c4d6fd1045213993782a74fa82de64f55c32b6a13bbcaa0355944168abffe2934f9fcecfbc071eecb24245950178a0369a67967bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c05270b4273417a567d54e305e857926c032d86500419791b168fde15a8f5dec0d258b58935c2f95d67d8adc64722696f285b740aafb0493588a629695186470ccd46460c66b7d08607eca9e9b096e97494e426e74ae0225f67b5d692213e95dbc0ac9e2fa1128e86ca1c534a3c953d4c67a328d62cebe87f330a74ae7f1197;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h691b5e63ce671fa3a8ecc1398a194485928940d3fb3d2deb08b600519f445cb56f5204a4d03cb39d64a931336f3248927360d87896308db7cb81fde184e277b7d91dce26c3ca2616a08f9d03a24a3e95c53fa8b1aa059398ec9c0eac4ffdd739e0f261ee24d64b81020a44f919bbea42c0377e6d4c581f263adeebccf6ab6e5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd51b3625d14584b0259f8ca03ce446b4402fbd63ad0f22851fb702ad9bcd894ca810765064b861074a5b3c2ed97158d6a2d48095996a0b9a8a4888b2ce2ea0301fe7398e794d7be07d126b0de14f68e420aaefe6300b8556c6123f8451d6b7f4cfa260f0df749ab3cecd4fa98a7064963ed2e8a7bf3e1ad2abc095a356eb3262;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8acfcf703e1b473df7c298bdfe6cdde17f008d9a7089619e464adabde82d7509bd8e76be12d2ec1bb31c6280f43f203107316d4dde4526ebad5b12016f73a97201a499515ea9a91cc7c5906563ac74157303d4a264119311abc584bb3581d0ea3c02e8789ba6af96e2cf7c8ac544a291e39032d715f5aded888232c1e487b31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h681dcc6d2ee0e8befadd7d08fba0a775ff123b2cb87f7ef391f641a7cdd1a80f100d2d02e89348cbeb5cc68e987d94436f2e08fe06de9b698c2fa770ec197f263c7337beafd39d61fdfbf0a532a56c76399254d5721dee5ea3e043744724da8ebb93a23b2bccc80e16b671ff05cc67190a926fb173491458a75d50b7c13e3e6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h509fbc2f081a4e4dfb4856c2d9d539eb4c35862d55d537d2564055bc1bcec0b9f3d6fd2eed8db14969d2fe1ec8626a49086f5e54d044d0ae88867cdbffe2f5ddcaaf65ed19cd289ffa7efdbfd92bb081209a89441f763271ab382f6f244f7979d195bc89bc989559467833c81f62db42005b26e36187101ac6e99dfa99501aba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffd5acc30e4c9fa57656927c2f1085ded97f5fe801b4df7239b769c75e852b7afcb0ed990700e1aeff2056a266aef2da0f80ebade2d06a3b6fffbd3fd3c9d55910ba85c90f0308f499d590ace3d1f3f7abed6279f9763d6c96ae33aabe1572530a4c8958374b67ba1606a684b9a4a41b2c7c1149a6bcd1910857a43c87394fe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc45055b09ba65ccf9b92619790739eb4c17a117072696a3164edffdaa23f558b029b661482e3802144001f27a6f93ebfb640b2f2bf5066b02906ef7f662adf07877ed55a54fd9c988ec4adbf611086a90a28e53c72c908b718a6d11f98ceef214fc3af8408acd0a4cbc5b811004078091c540ac102038a7d868849096a656c3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5ffa20292c9c48f69fa67b5307668b286031216abc47c550872460c4c418d77e318750e94912ed2e973d0262a74bc015b60c8012bec10f9410dcde4fcff034108e8fad4e87884739cfac98b9cee85201c26087f28066439c03ab3fcd77adccecd686db2723f539c147c1319fb1d01084fbf055697c358db2bde1b157081899f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h701dfcb81b81343aca0e6b525c6b3dfd21c2d55395e06e38e16b8ee04ae95fee072878764e43375b3b1cbc90a67e965a1150a7eb8527d737793dfd9dcde1719ef9f4a5034254b860631fdb2c3937c965cdaa2b3540af253063707750105074eeae364fcb286e0850dbfc46a5c2fb09044304b2c146f1daa9aa1ae1efa8e81db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47807fea45de7f31b4686783c8f8cfc8d4b89bc168463a72332adef43852e39dba33f8acb83efddf90005a3cc31e4347e54dd37dc4ac008b17b761f6399b7999a3a250ec2cf6deb52d7e7256773fa7d1eeaf530196d6b92ddaefe41b0999b47bc7058717d7b9ca5af2a4289b0e33af8304607cca25d5775ea684bde63497102f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed67e6791765ed65524aa3592e5354eb2a2ba23b824f8b05dbdc2b3c41d51ca78ca5af7a766b48eb6c9d44dd98ddf11d28e0551fe4e9060fca360729526cfb5db98a52541208a7d6196f6bac84c88b5b5f6e1d0ceb77efe81e4da2146e94b06b0a974f57a5ab5af92bcf93520d799aedfd583ff28cb79b03cbe4bc24a8ca60e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb28a6f7a1aa56d8706c52c0971160b330ee6a4be7189db9317c2de73883aaadb01e78fb302f8981c7dfa1edaf9752e0cda7bb3003dec5ccb5bd42f84acd3f107d1bc5dfd18b8dff3d6f349b16dc4e04f4a1741c587e79aece27113a4444e51c91f02b8997a4863ff262b701ede3df268a853c6745dc8221a2a4d464671e2c28d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h313c465ae8c63c30d5ed1165b64d74c0c8eec7a3f224aca5ef6e939433c5ba9ba1af80d253ba95e88fd118a7eade39d6a8335cb2a997cbde788fd61e0dd47318ceeda037a90b0ea387f53f2da62663e5d3b0de058be1a957aeea06bc0b4a48d02870b2facf18f003365324fd4d7ab62919e5ecaed4f52656a04d641fadbf1b34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6df117aa1348c58f0665323e389c053cbcc743dfd946b54a9d6ee4e80b51bf3dd4cd7250a65913e5c3905683af375c1fe67a8612f5da95117e461bff7843f33560654b04886a7d05a398817280f3424f06c6e16267b585fe67c92d9e9bfde48525a06ec91ac156abfb8dad3db0edb56f1c0c2dfa629435ecd95812285779e6f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc437a77774df11aa2663997a690b9afe300c159339e3bc47618a885fb5cb51db44f358638ce7e4caf8f5cd29e59366ad05622314fc9966d69b2bb8085180b7fdc5dccfd71fc49de1fabdd05c58fe9b9b57eed612381fd413198f85342dd43ea8787533c43973b6a443d8349214256b7c1f742fc0f47fefcc89eeaa7da33f80da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd255ab7ab0449ee4bf2316d17a16a2bd51fefe83933ec67efbedbde01b63b4a0fe3d1bff7fefc5839a37a8dabdcfe11df97c30b076f35c3639f99652d88c4c419e928541f1f50b461fb30a2670c791369682c6e04387ddc7a2ba344a1dec9633e1e40889a82b347f32a5f55d3e93fef7126a9ab1d9ee7e66438061414c9c2fbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h407d7539ad482c59f9e938b0dd3f1096ca405d708d905d33abc3946bda5f4467f1c4c08b5dfd25edb19925456e9b096cf26f5d326aa6965f6cf6748cb7387f13153bdcc0e87cda0687d24595ff00e0ee720f02a325f5fbf0416db37bb601a66c475c953848d2edc2fe6dc6ea3fb28bff4d4fc186e6914bfe4a13d19d24c23a1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ab06a69eb3ba90697279fb8bfaca7f318651e625ce91ef7245c3723efcae33bce9a7ca56d7955165e00d916a29707fe67c9418c4dcbecf8914ad273233472cc2bbac534a8209cf8c1ea72cdbb6589a13e14f80089341199125ade4300e232f3a55bf67ca67ef7692d973011b1da0a98a5c5af6c34a53a2e132f6b434dd21ed4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffed473b2d1a8fe6e4ed27e7ee820a5077a3e381ab1e52a6d5b5116660391b1c29ec172c0774ae5985ba385b81922f5239d39948cffeac626ded1fa16bc8c3156ecada87990caecad0bf8f444135975673f51c73e3002420e93521ccf0c2f03b3e59b9eaa90380746dabd6193eb7b468ab237e7a7a855cbe389329f929e23abd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe3c98900b2884992fa4d0bc0183874a5a3fc757ef09e197fdee5794e162f15fcb23742a495b6e5313f949245b9347aeea6a9084eecaf15b45d6f1ebf3bc506bc7c92b77ab1aabb1d0bc29c41880d7423993475430e45f1f52380af5298ba0812a449bc396f739656133535cf4028664415d568585031dff5f8d315809c89d0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a06890670ff6af4e2be7d5db50f46fd3081c9effabf8f8c4e8266719bb7a93a4ca5e6427546edefcaf990e9217f9a44b5faafd930e705d1f36acb2914d69a10b45ea71df7c4d66deec3c469cf72717d123933ed78cb56ebf0290ba7a63ed751efdb25c5468efbe345fa3c74c828fb4b85da98fbd0801153956581cd18f653b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac34e9460c58b73ac986ed87cbbe5ade0bb0971ab6d31eb6563842e5b673a28275e2fb7243d231e222aa65b24f6ad3a0f90f10c1e0a6c204476141eacee6f17794e0ae0076ad4e8fd66999700791400f7f7673e0181457140813cd5e818243a58a61f5c664e24e72d384285ad2f20c76638b2199e322d32d7fea7041f04319ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7294947b3957fa44f347180198543044c1562453f754de636a6f72e8cc949a61972f6869395c0c0a87106c27c66ebf56a417ff729dc1671fe0d808d24ff6fcba0fa0e9e49863745942b4a02cfe7c7a9af06a3b57abef80b5659e8839f7ebdace3fd36e85d69194583e0c1413d629c3c0da228aca03733cfce5d50c7795ad1275;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d63e3528bf640040033b9b45e1f91419c2ce17b302e499d80e8a30b4fae3781cc94de19ff6bae382dfed9e382fc4f65e4c82233fc815b1a054b060baf45bd6801f449dde6487522dbf11f434ca69a1aa3a4257974b8e2e25c914297a43726e5332d69f010d22edb2a3c5adc3f29cccecbc8a86bb9b4a338b6ea48931dfc8809;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d4e68f751dff35169de8701775df79d78537fe92371fd79479a3765a2f91340aceaa56b7b743d3cc7943d0b2d3ec5597dde1c4da29fd18c2ce795a2a714e791263850898f20e379d27f7539e1cdf92abbccbd90c341708dfd14e5d4ffe0ba869f808f7a4e2decd17dccdacb380472098e3b42565fea497d197ec839bba77043;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32d2d19a1035e2448320f9376f55dcabb123b64f2f426591e68481f75cae46305089e4dbd9a1352921d8df788b4dcdbe229da8961d564db4428601a9706806f035dcae89b9866282912b44c02b42b65b774b3226f4edacac4b00af80c8d00098e402df722cf169d647015ef13e2260a8f8ba789393eef3e3ab4bfb9ab5ef532e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10b879c5567eedc3a10801b560d85643dcdf7b7c2bbd1305cb8e99291b719febcd83301b0fa7b1a47b9debe4f071aad55bc749be67280119c9ca224b46325a4a6e8791ef08e7a0df68388f5739b7fe1c35d73e604123ec3875b844c951e332f9a4d264a9a3ce1fc2c91c2ef66c42b9117f8c1020b3d6c5f11d48a3ba90855769;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce49c803fe27702800c4741bfcbc4f891371d1fbd758a069f849b3b03c8e3520d92b0445946788bbddfbfc00bf56a4de0abe1666204ab3c32e7d231e27427688101a9a5c3d1882e82411c80f9371f0396629bce3f490f08db949e16a56f6354c2da038d79efdd09ade7c3af5bca7466e5c7662a0b24363fc8f35bab51c022aa1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a78f5d6efb30f44f9cc4acfc92ed66e4559bd1f471ff7a297dd60ba38560e631d981f1d61bdf897c0a7d1536d25c388780f612adf103179e8dfa393b7bce79cedc4d0702509be1794912b9eac20b074c04f222f4871a93dff5b3e1d4cd5f400125fde3144cc5f23ab04d059529cd8ddd5600622f9c177f59c96287387e7c104;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h315484ebee43a14e4bef01b5f9e26d229b4ca8e4ac858f7c167092d01b909f716215687d44446b7f5bcfad8636e1b660bd6469ed9c1b6aa0296a763fd627e065af878dee9779804b47d3c95c0e97a1c8ca1a094a737ccc0e1eb827dbaa103b44a48ec44c9f15246554647c6a5437e6959b1a773c6b5cbe318edb3236509a448d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d242c799ac5f69f623723e4e633edaef3448f5a03ab4f6d26d7768825ec0561d35a2bf556a955a27e46ec065d2dd2b0150ac7eabcf2a3e51cac63a4b8499d4a005510dfbd174b3b6dd19155e2d529160e31659e467e3f35056bfd7a4a513ca0e4069cc2aabab0b640ef2db66ef5741c88ed2c774092b34d1bd7e26c7aea9f94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e70d2e0f800a8307891ed8a9b0cadc37a74747790ce25519ea524ba732526b2211a979b7be0a94f434098191c0b380f291ac852f7fd17c678ea60c02cb7240453c5725e567a780de9688ce7d4a556c5d66168a7e8b40a6b7bf2be1502da3dc87775b1312cb42319cf80b9274d4163eec347567f6c710ab1ee1f96252950510f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha552bb29cfa2f315a63c52da9825fe8bac54a16baf28ba23fadbecf4698255ae5e8c1c4ed1bfbd8b7527cd5b4478fbf67256e0cb14d49cf90f9663e3d3eae9d73dcf1808e1eb1a5c98282ff99acd8ac1f56e024efba92a249e43be9b0f4e94f4e58deeec768414afa56bfb4db921656a16c5faf67e3f901d334c6871c2c3b252;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h714a4c514eded57f7c76bee7f4366b3b89f5feb67bfe9f322b474df74a68eae50124ed7440c5893e822bc9c490cc0184629e264ae24c7cc8e79f085fc2831bb9640ae423eb0583bddbefb99ee4581e7f3201cd6fd784977177f2f9ee36507e7a0c85e758187e94b24cee4b29d683d4e57e6c0783b10af62e8d03c6be0d6555fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffe27a5f4c9b1a127d6049ec3c3eeea47fdff0b160ac0cc3f0556393fa2a9d6a7295e369eb62ad47d782e94dcdb669e960b9ba5f49b4bd0a1ca837cd9d9ba9a03ba8816ea8e0bd0f7d055f6bccebc9af9c6a854da4f3ef7d4f5560e574d506eedbf47d7e342d87056fedc705de1b3523e37212f8108a14750082f4f6ae8c8b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72778c1ee92284050a7399893eeb04cfc3dc7be56ef4802234f170d5c76a06f8e338ef5ddaf9d230b76d50409c50ccd3d1a30bbfaf269e1c164225f78d43e48c3dfaedc97cac39f34ea188251a914d06e91b7525a865fac3e24155bc6a5553edb6fb28b9838c7326c608837869153beec43c9e4d4822e18e4c2d0e0bf5c603da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ad4efb643e6d857242c622e03cebe066f67ce6c7515351e9cb0ac996c7ae8966266d42a44ceccb6109756c086f3271336b8fc5a07ccf18a7a3ca15693aa7735e8eb401b5fee25bf679d8a845370b5d1881aab55638aa38d684e492d647820e42dd50faf18212644c95f286e27f8d83e3943a087a030bea33022f8254758def5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c1e48f2a7f373d180256b834d44a8ce07c11216b42382af6e3473e320f1351b5b57a45cfc1ec83547f6d03ea61e537fabd08738f1b22971cd96dc80788f430944ea75303a7103055c2bbc81e0c8427c1b985cde626f56a500fec09f820f181d53f01a98d504b4e11e4822d8774440807013bb46987351762981d6ab84a68146;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd7ae95a87915690cf9ce4e88bce808532640fd49664bf27f28ed5bee68b8cce589714127abe09c8b6b7e8b71da63853ce79a05e60e931eaf272f21882c12aa7f6eeaa8d248242e6e209db0851087812ff099b450220da03ca3a1f0067add4c71b4baf44bdeb7f5c6cc8a3e8be1c5a6ccf4a20d3e65a50c30470030b03fd0e0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1422f864854ae84b3b7fd9bd1bb3a8d722c62b4e05aad609570712a6bb1fea815cee1f8584584efc66e44135033243fc96bada09e50ce0e2495420c6d1ffd1d529143ebcb9435665e7333df703b193533dcdec2a3f06c1ea6b166aed6f71414fca6d813225d5eede8179fd28b0932315122d62022ff72fe0883747a6c78c6108;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b14e6cce89e66e21f99ff96e1cc723c20165fcfa383809a8b0bed263b09bd674c2ad04706f19c0e3b08af7365c0d696731d408b2343bf9a4bd201e37ab14f0417a053f7f49f8a4068a57cfe82498ab67ac0d048e0279ecf6413525e8dc35e02afa5d75ccfbce90a2a739808a79a3ac63c120ac15cf0c29611d21fdd7f9b9ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11bd8ae07064083556dd43790012ee07aa985bbd88704cffcc8b2af1753219bed008b4cbf9e8a28dcae4c7fe958f93c4fac8e3a570f76c090185aef824fc6de0362c2b6ed4f3717432bde8ffe935c1b5249f534436bf3044e20f534419b37a16d5bfc65b026bc8e1228a207072d5530a5dddaac88b0282ac0d02a6c04a050c1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a068c9261db3b1dfc404af1543b7c46168cbb161426f5a69ebbcb17419cc7e3fa0897b9e19f59d6dee5f94d5b4d1660f01575b020980dcf5ee664682f5f5284f50e4d416b384b184fd2ad6dba6e6b083e806418d26950bfd7f60251eda1e3e468e27e9ab2113017f5a2a1e6d60733603afd6564c7144d8d6bed8c4a18f75453;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c2b5ef8016a4c7b50448630dc44ad4b2a0287f7cea49fe5503975286433f231745df4584dc9f0359addc99fe79a60c5bef48a259c29a17c350753f99b3ccef0fdb15ff00530f2537a51ec293f44f2f9be8b606634ffaba8907cbd2443df73c3514f0be97de2df7693214e0d9340e8ec7ed3ba579f6b96eb889b8dad707e53c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8894df670fa7dd0b866e1594a00292b55d2352bd67b3d326c48b96fd6aa16a325a5352b5ef65ffbc355e458ce1921a80a3063de46b52a115925648d5ec463cbdbc9d04d25ed2f0266a74393b411904d753298aa30ad590a05c474494fce46c5e10f0d7e412e3d3e38e894d368dedc3e04c58338a2cb9ee9158d819aabdb46de2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb13755896fad3b0a5112c905e7f6e516cb1d0bedd413d73a1e432c33ba5299975e4be9fd9996c6e6e03d1bc2e674617f046dedc981c5c8e3cbf21e6d1816283698868d5d615735e83857577eb0a9fd5bef72f77ea3fd811380044ccf443c6b63db0c8be05b0694baa4135c5eae3760e1c62d7ca1a7909be1d8e305feb669151;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc72cf3540688f7f17a17882d3423ba74def0d660d5808722f8e08c6cdf7edf563a3cc2c27b88fd4ade3e101cf7f00f8390f825b05557347f830e7dbda933fe6d9354efb147f013523218a9ef0bffa9608cd7629292c419e654ef6dc5725dfbb5440407489b0226f35e9084e969d4cba1afe88ea4333dc594f7fedb2a31b1ae49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h737fbe86e397d8b6887bbc8df182e6700b0d83db6416ff1f6431baa86b2592779e568d4573357863e74877b32820621ce2e2f1016be0b3d5fded155ec353dd9bcec2b92c758ae2a30632416aaeed6b38ed369cb80bc6eb27dd8c0a96bd6ca19452dbc55198c634ce8ca9ff92873d8b1e5302b613e740a6024b86724afc1ad85d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb9003765120eb89c366b05e1c947e31db1cc47008a258126a0ec0f8e01585f07e07bebc86fabe9fba93d8b1979e4ffd8a719c7a4acc9e69bec95b6917e01f18c4ef9ea7c06c784ceaf0ac1b7a141a590f3a78e1a6e8d8b34dee7232538a6793e334b61a54f2f5335f25078202f361ae538bdaaa70f9a0fddd8da2cb854dc2f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f14bea98ca3306147b7bf882c506573634984f93b7d9e924c4c7856510fe9a4c3368286ccc6fb783111092dfe1d42008008e4700529c64b336dec84b4c93229399d8ca0d945db2aa216ac1d6fca011aa2b071a93d9493858c2fc79294c49d38fe9eb2792bd8799c6240c20fe4e5387542ea6d0e70ca897701d55b7cc42a88c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3e16ddb2f1d0dc2a25d6378ea98b44f2df30e959a6db6927b2299b604645043cba7ca48bb87141bf4387998638b79ce692b6e63855c1949c7b36ef7d952635ad13a005b994d8c1c41aa30e87979cdb3c1ee95fc1d2b292244645e9c502b37617855e594c3cf60513de10a2d7e91093486ca41d2abafcf3dbad9a2e1234fb051;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e4e21925aa048b054332e6610e204a55dc3606636b49a0a6de43f9df0435efd9a43fc6d95de888ad8809edabe3ce31a0df6e7175e532d4d51bc9dc442eea79b64e14426bf8a1cb7bd7f918007f9c244641b7034fd76f90be3bb0cafff6c01b140b6686fdf650226b4ac94357010b4c0282fd62a6923968a72f232bf5717634b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8865fdcd242499fd09ce6462e1436f8add9f5124762a5a09afd44a71fee0f59ca4602e3c7e8188f7267452e2d7a8e359970a720e70a3de39b0201e6bcf8c24ac0fc28ba6e1528ecb0940fdf82213ef913bc4b59f68372b372d43a8a442c729061c666d43d9d22042d5e58a106b4d1b2be431884bd2e3debfaada48a4892b188a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca25747cc4bff13fdff940ba4c2692185c674117575c98ba3927cc18a1c9aad12495dbb1921f2d1bd513313e4efd317bd02118b9446e6b7ef98fa7ee36c878eed79e2e3baca2ed8ec3c2ff413ec0bdcb8f4a5bbbfd0f7c19d3a23db60a04f8198d72ad8c250fb5be4c36edf7aa4356392c530c959d1f342325406cc70cb4cf31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a3556d2556d3c4914ee1f94f9875225b6599150d8f966362496b4b87fa067f3f5616c7c78c75a7e77ed1b106852cb28aed554eaad76eb58e3b0333a991abd97edc0cc993e88d8b5ce809ef762a56daa9373bde491d3ba5b603ad8e6e6626cea096188187d62d30f704bb6761a7fa77c29723a4d5e6c9293e132957a876afda3;
        #1
        $finish();
    end
endmodule
