module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [25:0] src27;
    reg [24:0] src28;
    reg [23:0] src29;
    reg [22:0] src30;
    reg [21:0] src31;
    reg [20:0] src32;
    reg [19:0] src33;
    reg [18:0] src34;
    reg [17:0] src35;
    reg [16:0] src36;
    reg [15:0] src37;
    reg [14:0] src38;
    reg [13:0] src39;
    reg [12:0] src40;
    reg [11:0] src41;
    reg [10:0] src42;
    reg [9:0] src43;
    reg [8:0] src44;
    reg [7:0] src45;
    reg [6:0] src46;
    reg [5:0] src47;
    reg [4:0] src48;
    reg [3:0] src49;
    reg [2:0] src50;
    reg [1:0] src51;
    reg [0:0] src52;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [53:0] srcsum;
    wire [53:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3])<<49) + ((src50[0] + src50[1] + src50[2])<<50) + ((src51[0] + src51[1])<<51) + ((src52[0])<<52);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1075875221783c3b94a082934fd8c318eedaef768325dd3947074404ac4fec536e19745737808a977df253f12aa6ba398888eb5b294e72fe72c4d248320e95a96dddfc5ed90d054097c52361eea1bb8e43fae1dac6227105b3433f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14673507e557ba74c5f29585d9ad693e5120639a94c73201ea6251f408843c1910ebc6d0c8c891c8ad71f2b8dc2302e069c870494100669507a9ca4b7b8cedd6459749357020627df0747e9da18ef2376b8efda4c427c1a35336c79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58bbfd9ec750f1ec12f70f62f1986ac7c0738b8d477b8093d428564a1d20875a42d2515c752c72dbfc0e4567bf84a1a000cf97be6ee7054ea2f15c2f34c7945caedd88b7d6d81b279ad6c01db5d4ff1dd9526643d1e77213be8c19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf60818176bbcaf98c847421def9d7679ca653a5cb82dd3c5497341105276d3b7ca957c85e60ff775c2440d682e0ea253f538f3497f92d926dfff6d05c1bb85cd411be92d0a288eedb31b27adc8361f6df1fa6a8178e6516099c35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d93a471efdcfabf2aa92837c4229556436cdddcae4118d79eccda93fe2f293cf768ee739ca9357bb7433a845a396465248bb384046c7117fcee70d101187b6227b139d4b5487d03ca78c19aa97a5cd1dee77b692a45581a0854da4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1971c4485564b9e24073e11a9680fd8cada4096e637bd92598376577edd37b68778f3c0d693d16ee9176196e7b323a251ff6ed63a779d167d1437acf44c4e918ce4d2042dd91aeeb2f535b965a5b201a2e496a4c6cddbe542067655;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd7628ec2b43121b2fdf05994118d9ec3085dd4b69b0ef94b01352c8190d1943936047cb0709117637b9b8a423ffc9121aef5d859ea6be60c838fd3619238c7674305551eb78c59bb72db4eced162fa853977253141c492d7ca63d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h857cfb7bd0ce6420428c335bc8f48de604ec33938f1a4938db67b79ae86f3f70b2c843d78763d9ccf9dec05a2a7d59415dd98684917f643af78992d27063955687ecae8dc8579b9e46d6959add473ecc6ddba9b25d10de722c4c3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ead515a9134e055dfaa8f7de863e6aea1a8b8a55dc38dfef53e8fe9b28c5815cfac46faabcf6eeeae8c8bc1b1c036bb0f7d33e6f78441651c123e2ad3a820f20bbeb8a051368db987b943bbcc6c6326073afb15b7fd7cebca2a04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1457f75ee6e3759614ba766f82dd5bdc1f51d693c7ad5193c42a87dfb6f6298e86bc43f6ef9520e37e66bb0ba5c3999f1cbea493e5fa263f71ba0f7f2b7d92afd8e58211d09b67cb4387e63bb47e854c819235aef375b9fca4ea7f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha35ebe6b370748e61e7495131cbe510fdcbea2dedf3fc15aab2fe13e2798128848cd22db8c9c4b384da444c286995542765e0e85cacc1464295ce9719c655451a3a3180f8b92fef528cdc805b7ad409b3d2c11491759efc41d375d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd7fe526171462bf17cbc46bff222e166be84041647f844a8668043011f02e85f59f654465d340e91fabf6bf6bffbc693ae0219d049af27dcf2b13454b4ea9377f3d0353ed4223d69d846fceca63e8bb7b9bdf1cecec4bb662d72e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3c86571b5f7acb5a60b437ca3cbd23f289f602bd41dd16f0ca9b8e473a4b83a5e49789980d792274468393abd1cc4538bb7df9b743bf654994456777e7f576a6d33a181cb7d7c65503fa66c95b5bade9757fb6a948abc34ed6164;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18937802702ba81dfb3d8c33b2ea87913b6ce79f464cf0cb7ed883ae20bdc355b610805fbd20666c68e5f4837539637a6aa91eb203df4a73e77cf16c2923fbb5a4bd979085b1fe69c6e6f248a862056035f6f0488e767e4de0e329e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b5468267c6183bbed4c8f81610ee49975cf088947888f211bebc216136de06d85106180a898966a9868bf7902fa3216a8f198bffdddb87b602723e0228a92bbf723dcb5d9960d5c6d2f3f9851600b55342900a219b9da4ffc90f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h811b1062a42453d681068edf379cf2e957c4fea62da3de1609e7349f2983ae4603100d8f36993fc31318f7f5b24ecba0781793832d82077f6d83f22287fcb2e5897345231fd83271dee15462c832de65de2a2454fc201115166b06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa28f094e083fbfb3ec3772c58d3fb69bbc4de52030705d197a49f232dc673120c757a9dca832160856cbe280509cc98127eef3d36284bcaedaa314670b042d7400dd926d0250189c36c7c926d5ef30bf7bfc690c2ef9dc05e004a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115f6fa541d297c2c2378450c12dd4ed7a0bd38616643f2f31e8a31fd3f4959687437d38a7a179825acb2d96ea89d310126afa0649cd0b2583518ff18c7e7ed8a9063de74e2903a36a17f0f6eed521753722a91b19a76784f0b0abd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de58fc4a41c82f74e213233391168920521fc030d9fa76819a05d25bfaf4525988764a154fe4c2c88d986ac9e6b9b691fb1ea5ce1e4045d98d936cd831143ef6b9b2e24d348d6c7a897b3ee3b3380ae643b0b26344a4449d86206;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18161ff96736b40842f26cf7787037fd568717369d70cfd3ecefb189c756ce4ffc73a12ad053bbd9a47ec995e3db3ba8ec005452af3db8bda270fe03765560164fd5e46b85ae55a56f3a97e1a62d40a5b66bd4e4715f897d6f95cdf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f9549c890ef87e52d69505a84df2f66bb410fd046c22615fb1bb7386df3dff9819eeafd716c029d1f163119d0223294370704707e571fae0d0b2f6e495ca23c04dc3523e1e992f7be08158939c04ac115ab0f93fdb7552bd284bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f6a95344c6c69979d1ba254f4158bd3cbf802c9a30d55e8edfc91fa13ee95860e3a7f43c28e5107c9e32f2fcb42a032a48dc972db3d2f3194e1b71ec53370792090d98fbe045b6c8e83c0c32bb9861ab2c2dc3a56171657940720;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h984048a7dceef5678b45b600825e89f6222c09d018fa8f5500b12c370f2d9fbd9326fdf7db0d97046b0f1d8ea8350f2cd21f6460b241adbb53d661db3c9c7c297a0c7c565957261abae201430d0d14dd0d0400ac7ebceba36f0c94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67cc5a3ae223c1bae964a7e0fa32e84af198f69af5893dfb1b6d66ec3b8e2f8c642fd26390931c6e8a8a06229d7e794c0d7591da89659bcc2fa878473314748311b75236ab31bd9f1883df785defc492e47754a77e9141ec6a6242;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51db832248d4d850ce3bb6d572c6cf0d93d910d731257da57b81df6b968aaf7ffb51444d551c9e89bb19d7a6ea4f8a896a0ff9ef22aeaf82f92ab6833d9b7ae86ce3233148283951dafbeceb1eff7b4a0a5a08046d41c974cc8e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f169f3da8ed0c2af06e93fbb6cf562de6c05497896becadd57f4a89e867d04cd4dce24211ecc6bd0fb5f7c43b66cebfe5441b4f00f5e5680dd2cc09eb12d7cbc33e6730690c017c0ef44ebdbc2535ff75afbe29df494884ea2788;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13087d34ab5f100ede0a8af521396667e1ee1f4940e27a265af5717164fcc9ea00871d7e1d471c7c7d5451941fb8c963bf88177858b28b70be09855d05d7ed69e44b0a48528e96cda142d0c5cdd3bacc5fd308674462a845e71c4b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192c60d0c718227e61717ee4cc2d2f175529a124b0a63bb8e61f5e63bc9a0da5159b17c38a784d5cdb5f2f7bd91abd25741c4b601ae22d207dc77650a80b4361b9dcc5c5481661ebd229c4db419185d204c1bcd6ee3de9ecad724df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16668b0c2ad5aaeab6eed4c7fcefef10da7af0bfdf658f5c99596ec5f343ed045b11e38165badac6f24854ae7211875e9edb4f877770e3a189a6bb68c01a5f8fdc42a9e9e6245b1caccc0fb69ab2eda6b4c21199a300d4460563d10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb226cee6904aa1d845bd1ef9eca9d89ffbab5aa45ab1514e003bdf155d01ce0b280b9dae9e57f475df41f5b981285f69ce7586d9ea87d16aedb7a5f710666e0cdd4e7944966e613febcb8c0bb6cd6e080f7fef67a510bc32e04a2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fb784bf026865664ee1251d762408b2c086a4e52f1ba92b652a14f9e34b502adb2078db7aa91d81da5ec270a76dabc33116860fcd9e38da71c2f52807de1cff23cee6e856533d2954da22da13f99b261bc97d2aadac87303c046a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb76fdc7e710d01617fa85c1931d8ab010e5047e5fbdbd91e85c2f3fef4b68206cc4af017756fae08ddab282ba01d368f9f4acd9fcc5b70016bb96869bbce6bd9dfd3778f55758d7685954519971a64d4fde8d7081fa6d29e5db48;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bce3fd16170b011c95f2f1cc08e7ba55079dc6fd05b956c0e16ea90273d7f63f582b71ca68ed8144186cd0de5a4e17cb3dd6858291bd9df018173bb3aafdc5e0e7ae849cbcd25ebc7cad8653063c51d50588f3cade3fd9e6648c9d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8ec9518ae3b522ef848023cd823658179762d9a5048214c58b3bb57be5dd9aa653e7e97501f6f341e79c43a54bb3daad27364d655c83d14a533d1db7e9477d951ac930fcda2c64c37adaa9002fa544f8e8dbddb39776d28d96e64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a87cdbbdcf0ae79fb01e61dcae1c91685b5231ccafb473cbeb0b40330d42ab70d1ed00f34925356f550a3f8751b1b5e09a0aac68c8d03cb9bde1bdb214cc7afcbbf441a0e2dd25c146a1602a2ebf2759b11428472d930de2a7f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4ae9e1f4b8bf05f6a0acf5fb11dd0c86383ace247bda30ad2744ab3ae544606a33d9d6d1779e980645a5d4a84e587fa4cba16a7752870285c44565a6b042422ce0220c1b962dcb96fc6870b78260be07972c16578946bfa248b73;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1500b56280777ae29aa3a66775e076db2e4aee25f24677fe61e0a36110597c71fcfe7a1e30a229ac90d2c28ab33f67b060476885015aa406cbda9ae18427dd64fb1295d57eea15bb84e2be40dfad4e1707b513d5d8d83e39ba729;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3e04354bbe18f2687d3ed65eed7b3b751d9bce93a7e37b1d8f4c965bc345fa82b8cb8b62881e984add2666a7a8a21916a47cc746bb94ad1b2e3ea5dea359be0191ef3c918a5a159668bc51e2871737d6908e2b70addac4e8a67f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9d602b29be9dc4d19620895939779c26d7023ca61a51e0f519a6c5237d0f10e3564bbf7ddfc2093557d915985e7650229e2d2801bc320baf6225cafc5de10606ea450cf78f4cdf610e645420d6fb25e5e8d3406f2a63661fbb7b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd30700b63cd92f7f139e0143a6696b9a1d41832f7e755ed02d5356d485bd80b4cb290d1b698d7875c14eead5b42653ece26c4f13dd815fb56c3ad64c2f6a6e01034aee1bd1b5c30d27cdcceb5f39b417f4660a2903a046eaee6344;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa12d8cbf85a834082be2244315c622377233ce31ac0f1d694842dc4ab96bfea8b03ad3d76253af28fe66cc3bdcea46510029550ec665f9393fccab1518272b3a9734dae4ffa4dd7f9b672c7def158c812b3734a35ec73d78cf216;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2edb8c307607c28d77f31ccb780c339d87fd73ee53db42518e959b0ea4fbec9c8ee328704141e43c530a1e99ad8e02163a828d00ddcbaa61ffc87406b826b91eb4535a10006466e700f36101d8c56042e753440be073911c973ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ded91259ec94896a31486452d05806387bdce0192c36c531c3fecf735d16d11a76e1f83ab5546377afcd3fc8e2943aa1d0dff223bba98cac82170acbf7ed62a8fdac74aeeaa5100b5dd6aaa081448bca9c447b9bb0fdb0a58575b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114f83bdbd9c4be10113fb3638dea7d1d9f9672e2e76e2abc92ec97021a5f1fadbc7bfa227d9c2f32e74b606091e137dbc53552e964791a9fe567ea9998b8aa5fdca12ae110b6eab7142499f91158191b75fcbc2cee5ea7890b6198;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee8e41add475c0b65ad2f4527421e2b94b2bd61a7b9a4cba0fc9bf0c1d90e1413fa54f68ee81bb5cc41f484cee825f22e9d6a46159d146cc8615d6102bcd83043cc95266e9c35248de7170034ddaf165f0ae3e88fe4f2685a3accb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he84f1f0c6705199368f3eeebb0d425187bc081a421cdbfa7b67c092558894a52905fcc4a641e2a9c934685c893ae136bc06d2ee9e8fb7729b7082b3bb0e6714d873c4f5a70a9d3ede2d5f608871bd86e36f816cc6c7206b0e78918;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6a5f972bb903f6a0130597cd4226618625c7663eb19b77e842acf2900b7f6dc453fa84989fc4a2728d23e80a90e2e79bc94976227ddab604986a81c1baaaf0a5b80b1beb85374f71a1fe225df23ef813261843b10383f5112d52c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha68c5384fe7f7344451db4360f5c739b304971c6d08fa543de2eab2ba9620fd0bd4cf4ecf8290d64f04943515de9ec2367ac3d75ad328eee0f62673da66ceb2586528bd666a033d5696ee697d6b8a9eeeb6761a8d873cb9697602e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139fc510c262f9fbd54f97b3cde2e910269a8b315d23f0296dac23fd51553e4efde5bf1147fd699515dd5f44d156932b3aa43146d7a2a38980f6359cf7cb0fa41e6cd8c2ea69b1fd61b8cb94a9de8c457db86b150ea8621b9e90670;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e521c13c6249f7929fcdb9dc93bdeddc2ff41df828a17b54bdfd7c358e8d91b72d19eed07ef22369293464c1f3eabeffdefb804e70641d90639a8ecd9cbe17d2bac22b5c93e9eb1a6cdeaec32839aa2a7027848f5b1ae687c97dc4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h543735589f5372480e6485adc8ddd36ee436b232bfacdada8a5fb2d6399acffb3b88dd1564e5e93ec93ac8d026ef53a30260a688ada1603e9d269a848d390af1c9a5666ea90d039b2bbe40a46ae4f6af494ae3052df9c89bebf0b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49ded4d2fb0580e0266ca5d51e1a511e3b55d21019eb50631be82978950a8618c0caf05334165b3fcc56d0d53cdfe802fcc3934ede098659cc271379ff7c1ee58e3a1610e4ba1a073da078d446648b958f7d5d30d5872d13ee3a5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96d2cdc70821f459ee090cbc2dfa9348452dc2220a8bf6c6594af681562119ca38d13049b9bce41ff93b5000bb6b94d877fb243432810a377c7e5e7da2a9bf461ec0e5a42757d1e22ebcd5a9fa10231d7948566be3d74c777a3659;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110cf38e6ae41427fbe8a0e13b128fe555b1241bda48eea5f974af07bb58d3edea113e206ff63c9c6239f312223d036762a44b673cc4a6128d35893a64ee9153aeef290f0a4a82021d15fa492eb3850bc8376b4dfcb9760d5c154ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h56ae01133e439c995c3668729853ae40e6f4b78e01a70ef503801aae64d942140861119a6e1d534aea04dc6694b88cb3c90eee9b6b152b873c9ea26b930a5a5530fe5b5f7b701283e342b6ec91e5c00b8a73b85f034ead1b777fe7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h501f240f68bb375b0809959e00d08afe136976cad95d692470506238955b367d3372745615388a4e8dea9996c53976956c5a242e55fb1d924c731e949fd91af03a8c0e36e2ddf4049da07c12349c53e2215f1e3aa65c2659feea93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17071db87f69977eb39b49053141d2da78d985bc2fa34d03cc05e06a9dc37045868a82de3884d8746171c57c547d0c4f18b9474834d8c88ba080542e5a0398e389e36c31dfcc6775dbab799621c55f96b2d6a06f961e22a8f4d7418;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1686e78253d3378306403bd2b5184664f157de2608077a0d40084f20db7975d6126ded6b8ba68e714860698e3e580fe8e5c23ef5bbe559ad9211466f229bf486d2858112457a75d3f3d8117e67d741040018ddf0f9d40a7b7799a3c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1131514b999d9f9ef4009851e2ba277583b43fe669a3282c65a308e4171f113e0f4bb5b12b9c1f20ba88d61835355ffce41d52f96f4f562755f5e8e14f932d5fdd6ed00f9c13ff09541f5efda348568a352bcf9c74241df6e5a9be2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23d3db2fbdc5ac1214a04a355836d689aa084bf6ab6f417a7fa475258c8cc096b9cc3a52c5f1624a05be070eff754c682c12949802f13db0f1e067f95a8d38eed1bca345bdf25559bf5d8ab9a6f4bbd9700137dfa5e0b883fe8ef1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97c3469dc1ff6bd2e4086135064bc4f717c697c895a39e988de02b26abb7d0ebc15cb43d071337b3d2f8089a8620ded1d44f1196427a7b4a058f2e521f82a44a1825841e8b5f593687f798ed6fab929937dbf5c99f31f0d8227866;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14da394a514f2359f40b1307d7e0a5dee02c271d289a41666e13e8075b3f47915c014978ac313a6113cafc69c9598b2027e9d6e657e673762ef0e68595317af6c7d99c2b6fcc3047213c5042c7aefa8403a20673c491f09de04e1d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d4bcb7ad7d612ef2f0e7d90d5bf0f5a8ebcba3d81775e9684baa5324d6c402d398a700feb7a1fced6d6cf3f0ce3a6841a9a56ad38d8c42efaff3aa644f64b72a7a1392ee8f5c828685c1b03fbcf0709f1b6f9411ce6b22b4634f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf1538ea15db8e9f7b9af30da50f2f45dff2ad45051ac2381c0afe349911ef3b785dec4363e12da95a9c4858eacd7256116a8fa59c68c26827116d2c661c190efb033a8f2f05c34bab95f09f4f954afcad53e4dd76d7eb58340b04f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc85ba63512df4742567eefd6eabe8609bde020630735aefc6727ebe5461438bcce25a1d2beaabb8e689ebba0c482a86b004fc48bbc0a7f0edfcdedba19c48f440c229a8ef6a12afcab8517094585d12293863826f5e38873525729;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18565a9281fd07d5b682b582c7d3798b10c93948a6c60a52aed4e353c15f2406be10077308a21be16a33a69e7c6e061ec3d0d524a60b9e64be9c1de3288e469d71ec636b2ce3f9f79941a5bf388d06ede7be1abf6976bafd96e8955;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he077198bf5139e59e7049f0a1a43d187d3b511edff160c8c189976bf0f9a33b5de597fa460f18ae3f20a19aa089b3758db13cb49247698dea7af4234fc3e85e3ff3b2225c02e752fa89000fe6c57427e08022d13f2814e3875c09a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9dc16fda3de26f1c261173a43c820d6c76dd0381a59111b0c8a568dcd0bf48c88b579cceef167c3fa8f5be33a811c4b70fa94ec8e016e4d729572b3fb15f85b24672d04cb094d41c87d9b7f52a1a9e7f8a4baf04459d9130232a53;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32a0a829ad7e636884d94f24106835ab641bde2b7a7250d98cca34276ead66656b634b0366f39d2dbf42b40f157e62b860e252de00bc39a988dbfa922c147bcb59cb1a0e7fc0a8d90c4e961126f3db86ab48c3acd8d27d04f9515f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f85d4a2aee38e49aea39f9dceeb122d70ff79c49edf067cf005bfd062f54b0a7d2fd6aadfb279ad4a531d443cc9d873c6f6a82f8642b2bf3d839e3b694987612699c21c64d993d2ccc4e1de031865b547cf46cdbdbaf50399f1ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6c1c2e21a227c92751feb6c4f15321257cd9b1f81d5666afe7c888a8686169f4cf308f2a81c4acaf61a7c5a35570531604854bcdee552f27617d384b1d72a8c7096910ca662dcb5bf173219672af323b1e202b689868878c02553;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17aa36f0cad62f923ac8693cdd1b39df073874becd6c19bc7bfc78cb44615f8f3cb11599601dab61a496566ce9a1637992aa0d446ca11f3442443e3bd5bb6e86db573a1e0673f2fd640be07e2b0cebca45cf16b0e551df6e1713f39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf502f55ba567a071c9e7f2a5b4de51f4b209b3b003f79a1d96b7641f9d29f92e8465d58f28d8e6849e27a3c43f0b8e2dd7cd543f6fd33026764503494cfbf1622c2e746dd2ed9609c56bb5e455ad5c094ff4a6833bedd9ed72b68b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc10831209a0463d1a15bbac28efb37853b62af092651f5e159a69b106f3ec07243cf2416e59281ee250a02d67314cebf070cc49bfed313086eec9ebc6adaf9617f68a201c3596419bc43389d608fde46c4af4b997757cb0f3a09d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad6745503232ef468436bc41601ddaca0b4583a1bcbdc3fc6c1bb19ee46c54c4f7e084ec0c49da0d20f26aafe8fc492f80a74a7f287b5c8f599e1a5830ca02a92d50e1eaca3ba240ef4ffecdbc3694b00d77f2d1f9c5f1f91c4bb6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h665520743cead8773869eb694a9240ee3e59ef0b9cff9284e370da468c26faccd29460056f067f15991bfa5dc51b698b6d5a94f8f34db52bd7e2de0bf057034be89be1e648588117d27c38046a5f0a81f6e01da83f5ddd4ef0d986;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7043e3c219d4d7884573773afa6ac8a1ae352b1932a048c9dbb03f211c8aaa8d1960c3187553727a63f1cf73dc79067e331d19a4df117d36f76f8baba6d08b24f5a48e73df6f7065c8c1c1a58527b9e58d151c119d1081db0e17e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc85abefc6077b4269690dd79f49c28e8036d83bcd630ee0b28dbcb564abe15befd3d30381038907661ca97db74773401fe0142293ba661fc893de75bedd9f45067f5d3f0dd227a20b48d098277959bff0d14448be5020b3306fe2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2400282f432b5d154b33631e72d8f292f2c7486bdacf014a4ddee0d0c7f1b6fb709e8b814f587c99d2c09efb1ec5b9da5a1e9a63519de4c42b91e90e470e33584a45cc1eb5ce78919018ce6e99b99004a3356919ea60c54a23557;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185cfeed6de979d729fa79c0210f675c26efe99c70bf377b102200f5a58f48b38241f0caf5f7af1cc5153eeeaaf92fcd304f70b690d65b2e9d2cb09e43fba58fbf7778860b5fa6e7837205355e293bb07dc62bca615f09cea0eb6f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11044f5afd5818532f539b5992075d5cba276b66ba593dd07bda78d6ac3554e0f4fbed4a12e8361677e0d25988f3fece9e9f4feacdd41a910a73e18f8180128e9e122734787b4c82ee1946a446e345fec0557d69bd3d234dfce706d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc32ddb5c624e7c2f57723531cb63f6c9e5c15c901f09e237a3de827263bf91166270c2e59e625c51ae265766175afb28112f0bd24edbe4beb0324b17b5dc4c62f7a2eef19f00d1deee9e69babf4bd0542c2457d5e15bdcd660fbc5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be16ee02e2618e2a6312dd4b63569cfa46ac44424a52fe82fc8e1df7fb8637cf4ad7da12c6adb48d6c1f370f15861087be116124298f8a769d9cf5481aea14b5a968104d557e550f956a36b1e1686f13641c22e008fff4317c8cd6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dad735fee4e47af8484f909e7b32586040967222f71a93d0ce49b964424cb8d73f421bd6eddb1de4fc63ecc9a1740ad3a2a436cd77fbf5a687d384ee1702c087fd12221d94416acf484fad85eb4fdf68f7e8a7e70f539e72bf5afe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdb4de72a3a107cd183714b09654695fc1aa2b49b001a87c1f169bbdb8efb3495e33bb221c784d9c4b4b13c5acb3f73657dfa3f2973454bfef56a3edc40f78136d99d44fe97146897b499f3120ca40ef0ce96780ebd288b41ea716;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2175439c777fa678df662b5b85acf9f106a3017dd0f1f58b6f3b3f3ca40eb82dbe14812b2c3f2ccf2b0fb9727f369687eaf6abb4dc0ddbce0b584f040bab0a2566d112e13ebd6ccada88918db8e32c39d3dbd688a3c9b296c8632;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he442ab1bb33c3f1ebd7d28111fb32bf06406db7b313c99c70268fbbb8d9b61449313989fa965c76236004f05090537316d13588eacf6d56df9dc61a236652dfa1dd41fc752dbaddb9f8e5ddbc24e54217527b10ff0a51245cb53d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a341d8c4c3a22646330efeeed1df60caae23c88092f36b00b48111072a752581f34384df99ca469d031099e5192c28bc5b6f82008e81f925df72028d40b2a15b333667a35ba9560b8059aa8cf75a0c02e10bc4af15ea71e355e4a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8784e7c47fa010f99c1dc71f71a2abbca0067467250b6566d576e9e1ce5b72a488b0be3bebfb6a7816a59ca5e0d1f4b06fa25d68e70386fa44d722b0bd98a9ea8e9c44d68f9385419167ca81f597a46175e73c5abfee022863e23b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b29f02c43f0c4fc4d87490256b1533df6e2c6c99063fea2f28ee4ae959956dab202dc4cce4fade13b9c2b3d44b647c9fe74e44e1c7e13b50e1c2ef606f4f03df9bfc66e71efbe27fdd4bddfa09bd3e1d893b42f26671eba19ae31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha98600c83644ed613a23e94ae3e63350f9f5931ab6a2d82ed7290b8ccf14d542766a44e79644529815d9c1c52a6ce0b76bdd79c4b5f16a94abef92585355ab038a2a31be95393480aa7d39961258fa25902e22ac62086bf2279860;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha631417bbbab1f6babcededa2691037495c81974e4d5d7dcdf58fa110d73a7125e2924d42c261958275e48af5d728d7789e51dc901db2f25516b484b3f669e7d125ad5f7c23f45cc7fed9a1c649025fec6995be8e03b07d4767bc8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1271b3c8639cc9e7e59faafa8728d2008272314f76bcc42670a1c4723a461cdc0d777ae3d275eff1e194ca5c9a669d8ec1b4f147b894d23dcd4294abafce0f0089458b768ee284df933976c510fd5b5f203fc5193d52ef00f7a61ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c2abc69bd20e1790ba46230ca9ec5116400c55443df077e2766c3bb4591bfa2a0f3fb71c99ba58bbb5bc18e79451eb98327ce665080b731db2de2157b2f98f5ec125fa61f52d0974c8b5a16dec303b21ef1537685f0034b0c93aea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ba77865e24de114c71f8abf5e677208078a6e5f9c5583ea51a7fd43d36344b324df8d696228885c4667cd4948d1a1b984bc484795c857d9c9c7d3a43ee538b00d44b6495ec930d6c01b4040f4c98a9c6cb32d4143474aa8f8c693;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a584336fd6614938ed7b9dfedd9517fe71f2741a17b79190d0d65ee9a31fd8bc2bb426d20355936f4bbc6e11684f38118537291697f0f72b859685a3ec3e1f3e6bc90a434591b4855a7df2d0e841dbaec1bd47948ca88c869f59c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46b52c3fd54aedfc1e128de48cc0c1814dc15e3a61aa0b8c2efe1e0c1632ef1d3f109d43ea8dfa80e18c03b85c51081f19d06ad3fbd32e0b8a4481a2c84deb43cfb8b97a6f762e52e8027cd6f024acb7c5dbd1f2a086df9f54bb5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81ae35ca91f7f7dffa1a0b980a9e2313b5030169fa4f595227ffdffca3256307a69a0acc1cc309a0d7ce37f491454a39d32f522130b264706f25428443ab044ecf5d354db776bd16794a21e53ed28ab5c28731ace1e9bed4c21751;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec9fa0b5a709e34a57a5c24ce996aba7dbc313d94e9b5bb6095f8620e437d3f01a1814d6fa770171d30d62bcd2ec877e6117f1418de9c6c3161b0999cf9830750caa23027c1cd0e5a5d26e3120211e56e68bf0ceb0cbc1b0de03bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d7931936672b50cb63c0393f39e7430a518ed8ac65702723d2d3dec45ee61347573981857f14f51a85dd20807c67a3efbbb21aff715f1b9403cef601416193784248e9714147f6920edc034a40f6b419cb7595eedb010e7ed1c49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f1bafc53c4aab62a1121db07db3d1ceb88dbe1c9c4180c3025fd4c355955aa03f43728ccbb02366739859f81f1327a935a3b52c1e66cae91d8c1f64995913ec2b21b62e63439b226d0f7b6c0a5af47ffd4b2e351e1b09cba6e157;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8606387ab3ceb4a221662c647bb3ce2b7b8a09516dd9d10f228f5ea754e7b9db30cdfe4ae6149a5553ffb47c94fd341bf55ce5d6beb4160225000edbd505b579c8777105d87204ec34a9732eb0f8227353343c5dbeb51088ac46c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc28202b86d58b2b0f5690f169f92d241be9be0b11624e710ba11a1e12c6c6e512b93e7742b211a1bb8509154377cb47b901a96ed75af4f6d0201972ba819a01d163e33b92ca238200c7cd8f15f06c873339d1d533d4de401dfe1c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b78c7a6c45cb6d3c2da7d088afc11fa628bdf066f6be9b086cbb782307b1bc691ec3c8cf91f58a537595f457e5aff5d99a835aec3d6fe549f1da5e57c332bb35e70ec9f550c52cc51bcc4666d8936a35405e029f306285286b4e35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fc88f8570c4d94b530c1487bc8b44a388586f714991942a0762628b1e0c0c505e75768dbe7843ec1d1f5663cac9f5150d9d14e64bbaa28f1108c8a5de943cf123aa086ec899a679961e2ff999e093810d95da26a633867c07a967;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e703001e325c420865b75bbf403d14d7fc69e916554a918f5d474dc1f33a1b1a08dfcbbd70c1bec743c6df2f0629c6446479990b0ef96129ac7900139e4478dcf9e6b704df1267d97cbd6e241b573f9372e957ccee96540390f8ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158ef6932ea48c980dbe345546065851ce09a7ab79130ea13b4c13ac7eac2e3ac05f9c67ffa88c7465180ed72d4fabfefe1c9ae6affc05ba02a63a2a8e67a92debab4616b957f6ad92a1d8a6d0e6ca09eef5d924bd02d09b726ba06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9cec5b403682f195cee44bca41d0c717c2236ee3ac1d6f97766da3db9b2f1a40aa19646fe031bf43268efecb1ecfcda8886d383de73825742c9097ed413eed5c15335c8d26835f9579c2a98e0ae57d601fbcbd977241146957b431;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6daa17b670572083fb3147cf990cafcd9f5f305f77b7262b34bbd0c00a11dd559d254097508f9f4988816a7dab9564c576588479a1ec3a2676cb62b23cc351c17c8936c9029f14a1dd26002b6f72bc5fb14e34d0da8b4431e25126;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1dc4ffbf38947a603abfb79c1b7194c97c08a253003e1f42d09a57694dfa964296a169c6a7eb7a7f48575e51110daffe3e470ef46f4091152e2b464f2bef3df1733a64d0d9ec1fabfc642698d694b66005e94f3ffe004caeca0f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1220098e9b22d5177f7566cee5d6149b99ea63fa8a2e78c2f21b7d138055651dfef2e39814e233a3e74d7286b673d3c0953daeafba994452a15267b49f5bf8e12f080c54a934028b6a73b32f7e311e9c4aedf189f0e5f8946237d88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5ea0a74da61c173efeff5902bf9afea826aa44009107c34bc35cb47ab437c70c47ca142a3fb3493e1790083797e7f9ae206e2b72b9c291d0be1e0a3e4f963ee03fac1484ff8b9ffdb5930e6de88c5f6b0957041a0eab7c21f93ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd305791381f192032963f3bf37ab492f08038e7c8098722cc8c5ccaeee6dfdbc05ddaa8df2cb2e409536a694286a3ebe2f577492805afbbdb432b40fe91a4cc104c0b7c8e4e3fe73c7c5325b6497c46693d92c902ead17a734e349;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aaaf3a451d65ac908029e9f05c2e194d7a9fddae100f6418c2415d4c79117214d5e8a0e48eb7310fc10f84a1d43d48f7464b23d2470c7c260b0b61c32c38be5ca1b5375738120735a32ae1a7b08e426f4d629670e3e58df8ea37ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9485c7040b4bb87989c118d5ee322930b2b1c3370a0800a17fdb473e8092abc7ba92d3fb8ce0d5cbd3aaab7b89d94e666ae771c065403b2b0f5283e9675ddc4ea2977cced002fc7f06e0b4345697b35fb895a907d343e92e35a31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6ea211f4c8281ddb77cf648808574d74f03fe147e2d7fee5cdf4b6bdee8cba258adeecd5984fb962a771c939fa323e41cebb8f3ee330957fe5f6d42326926deae53897907231e435ea33beb51f0f15619b953c9e1c25c4b5f594a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a163bece5aa26710fa2953e77ef3eaa0442021c1e23bf37fbc35f367f348eb51e77fbfb1067823378af6db3364540d72f1c8a82d5109166bd0d6684c789f90c7fddd69a6f608fc401fdebaf2770f6ff36701a53de5f657e97e158d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13abd9009f2c87b24beb92374eef2f8acc4449543625398332dfcc314578c2d1d708c434cb42c3cd66cc2792c3cb202ed2ad3c9cf4fe23ee04c6dc9103ccee7732127a6c6e01d9cf532df45776cc86a197d32b4beffae8e2fbf958b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f73959878ee58a2f648ab7f49b908f82b834c45e0f8f0d65c212f8f8bb6e3a1dc827729cd50198e0fc8f3f8c6398f780646c3a413a7baf190526e0b263763a56943eb3a3ca7fd20721f3ff3794c32f73fec918802abbe6852bdca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1faa6ce25900a06666101f85af15b2178d4fa4cf6fd4febf9c0d5caaac7d157a1e8aa8dfac3a3c6a12eb9c46e06b2f91edcc148a030bf583ae4f2d3b0d94ffb00ec0da2aa88b433670008b2a8845fc1bb8853f903b0f6e77b6a9e9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ec77bd9b273b66babb241a17c661929c4c976381023c21bdf9225f7ef53e8df4b8bef335849cbb887ed7fa78b53ae8f636ccbd2af33dd3f765893f1427c9b416fc4cccf5724a429c9e7bca903a12ac70dc639e0933df4861047ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1975efabaeada0cad0947df47599b8eca01327556e8762fee80a2cd89ec6a028e4a67f18cdda5c552d8c031dc6ac17dcd89946a35ef00c52f79fbd09b0a467b69a085cda7360993ca36f62ea233ff36c65abac63c3d40f775495b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1383fa32d741ce3aa1f24a4ae9cd5d5f916cfc9e90d14a747c29964cab15052e2036d71b1cba2f68a20a5e1a87265d6fe3fc43ea4cb1f33cd0121a72cb444e0b4cd7439d4964e2ebaf5358a119cd94e941aff8d81e7a0e1cb162f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f9283ec65dfef932b68999625d025ff8d692c5937c41abe2b066c0d394a8367f83ed674035a326f06c837df01269c95c5f52932f7770e52b04e145bd5f804174776c8029a613761baa8a13ac4cbcdc4c374ebf10648f2b6a0f8062;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e951b47bc70bf7bf8f36db4c63fd208357594e567d6c33cc68510a29811aafca27c4faab3971e3a4326d47a75ef1d0de2d6980bda5e4bcb26213900a2dac1260742caa387f8853142c63045d22778065691975ea55c56337b992e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc296a99136448ad73941cf0955227541df833b95917c25c07a59377fd3077c8a9dc1780d2939c6fa15f0dcc811911951771b76bb1fdd109f0406b7b744e83c9173e180984bd1b66694d5ebb71f98bb79a1c02ec17f5f5735de702;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb16005e163ffd0e58cf05b65621324b0656409370a9f97b70ac91b5b480b7170993de43a875d7c5951704a6b2c7a40b9f957da5c94b933e368d83ef6dbec39d2bfe45c87ab8344da06853c2ddc0337ccfc644623c5fb39a52fa658;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbd35223acf60779d6f786388bd890614fe61bdd090cdaf72e0f7be26c6ae092bb5566e6c69c4ea2d35e3d4dd9e33c7709bb62a5d20c0024310c7ca06d1a83bc2579ac6d7a9aa7e188a4af4e88adb664a862ee629b7541469688c65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0cf6b94ccf43296021787f0160e023a5211b86a09ff569501d88ca5f27cbba2f79e413928fd465ba07f0277cb24f93cbdd383d706cfe5b83975c49fdf3b40b1d6f8872968b20a18785e7e468174adde8d7178abf8db3772f738b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha237e848bb89890b9f81cb3faa77b411f57eb1b65725dd386b572394e14e2dfb4c005b15ee3b3d26bd9e5bf5d0c12cbd7def177180027f1a5b2f05e2188acf6baba18e7707070e050182f2447171e1e6cbdff746be1978e5cb975;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b6c83e630d8d0068f2cf8e4f72522617e905f317b283df2c2ed8d4becf9d4e41b85f02a71335b61c7e03d521d4830c5bb56c5f997d556429d7ffb81038eabec4960dca310da5bb9cb970726215c4ebdbed6fec0195d9a55d657bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3cc63a4608b7f7153ac97369f006e84cd613f5aa5b49770e8f14be3c316b1289cd98469ec98f5b7b038adddb815f6aa75ebd5df43cd789ece2dae85b1c61f855a22ee7d0880989618bbd2be5b2dcee87e55a59d67823e51af26588;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa25073ae9779ddc0b22a12e6cdc037f41796ddfb3a22dc853d48401e1a3f9e62f26197d39abef1ac09a63cf9dcb3c7f9957c4eecc970427056d15caeadd6bfaaae9f711ee9b04d05cb612c4de88ec72e64697fbd0bc22b3e9250f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b1cec4f8481994d54823d17c464d69accff556465d46091b9538feeb164c432379cdc5a5211671016babade7ed183c67e678b61a5eca8125db376ddee8db197d3e5713ed59ebd8b983ed098a1704d2ca5221752a74c0be566193c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a5e32963bb8a4ba79dfd52512120f3f6035b9b74430eadad8f734128b268b4cfc6e76950e272637a7a79833e5aff29fe4b17383227d0dfe8bd668080684f41e8e46a65258404e05c0aee1ea06105f1986e24039f255f931eed98d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h690c797e095e8dd69c4665df7a15cfe73717c37fc2b9feab9eaec8d8839179971e097e266cc024d6b135f96324f47461a7bc0a225a91e06fbeefa53a7907158f0d4bffe8a2e25c93df07b624ea53acc06964d3b5051700a1edeb35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26da93482828604fc05d46d48300f0b7a98f1b9ce41c1419fc59ce1fb98a7ad5d120b214d0051792fba99c9bbc1f3b0ca54cf415a40920d985e9667a3ecc15244b26220139a6b1c8b2c5f76a2b6eb7618992bcf766e6d6d5e7b8ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176e4b4566f23df0bda579628fe71b9dca4656082708e2e5bfe9424488f9fa0b0ab581c35f4b23216bb4b5dcffdf905c210ab4fbb3fde1919b8984ef6cfa5aebce96e701a1e4fbfe5d546fe7feea0f804e35cccb22d6faaaf3f82d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2e52692ed49147e94dc9c885ce5873bee4b07f4402321041cde41597fa9175a1f09d11e49df119eb5c188b4a2ad9d85ec63e150092218e39aafb6f15e6fb042205d87e6b6fd3b849c2950288f0957bc9445c2911d9b960216bbaf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18046a348e3e1930349bfa788e082c36cc2fa3c99bd37c6e91faa883c308f55c25ec48c45f1ae435c86e37a4d8a3ccf5bccfb9f86584ccd379a0cbbcd8f4f9e0428919edc11a1094e67af138b54177428c59ab30b32c63c60481c22;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf96626ed387ca8ebb517f295a3e5fb3eb0b15ee33df4d2508da4ecf744b1faadfad6006888b5298a48de76487600246dc42a07cdafae97d806a04e9e54b433a566ec6c5e896ac55d4e38cd51250bd4dd8457cb42b4ac25a2d86ad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed9be85b95a2ef6c3e36d1a3245c0dce08b2913edca62c6098863a03ee752e1f8ce2611c4d867e81c9d4bfdb43fd352ad3fcc90651fee35eeb65449ac57487745f39eefad5449fe6a06504c0eea274c24ba1e77acddf5f893c5738;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1510088901eea6e0cf9dbe6be29cbc4237e65841c13f163f5f75ec1897382a0cecdc109c240ce36af368a1e8e626a9d6a6eb090ce31d2e566d0085c4743959668c7d196077d1afc00b194cb62bae716730ca8e858e597f4de4eaa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ef994dc8debed7ce92a4e900c4e00f350ae0202657bc8696bebd4494a1be79fe9ce528a6416b194d96606567e4981e7a63929dbe8a23647c5212ffef216fe29e75144d173f6c187678ef24ce5ac922af4c8d6909f914385ab9b9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c5632252878f8ab230998a3db23a578dfddcfe526bdf4b5ae95b6e5a39486cacc3619c20a54f3d107816126b163d5e92e6026c2209735e2c2457ca6ceb492f334c793c08277fc7ddfda6371dbcad4d6d470517412333f5509f6a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180ce0b56a69e46e6fba26125ac2a16924175b924d6f21b1cc3fa7f945a1cea0500065182d0afa303c92aa6301c7bf311e08bd4b6bad781ce59c373144ee3a7d6eb06f3030135f09c668cb68ba50803795853be40ead1caf3578541;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b905130fd82fa0c7b74d639a2f3f67450424294cf64a1a627c28e9c1340b83883b2c71c14814c127b6099630ecb55536bd827b3eb8f5f772da39a8eb3a4f9d54b0f9e7761b69ef0dc985cf4a7066c6cbd249476171309e6e85da6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd68c8e122ac5020c7cf02f1d44a7368bf375f5e8fc4defadd34ea17579a07300e3885088411c97a40b87b7e2e72c2968a47b5aa65e62ab601554bd18f2875cd6c64f2f60dbf418012fd520a8f06b4afb54eaf0a3fe2452d02c5b5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102fdcc2a3c3c8a38f4fbc6b2bfecb517b1d895fe3dea13dc3ec7e5cce4a718d3b1be3126f60f454a52f14f1133634d4403a8d8f671a9bc96588e34753129000e17af1ae073c210795941c16c06284cde176b65443f5e06b72197f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdc07bdbc362249e3744710ba235d54285c9d7a9bb1bdf3f04f2635513ab06b7f0e9cccdba05cd898021849dc2171b05482686d305d5dc24c4951200d4e2c43380aa6b94f4f7dd887c7012f9ac53f16890e60270908faa8c69d9a1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14190fdcb2d38906fa1e88032d666f8e824370a32ea27a3d38114284428602bf9709496defc260cd8b397bbb9910b8ab2968bf047fd72e166b566d447639bba5d5a22a210b6944cf5acf4399395efc460d2824851a34d91ddf394ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abe55256734f5486dce7668764e552ade827a942f3bc06fe4b133c25c2f7b53d8719df55fb4b13152de35e729492dd3eec58110487c77b8fd9ae477177dc177254f023dcc096ec5a2c04573594333ef6b6a2591c01f2d5679b0af4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7970deafd50fd7cd065f483fe30bd226ad71ce028ae0461ef2dd49c3d3f5af53bcdeb88ea75c1fcfce2e2b6ba95061ad71a0646dff89c0e064dafb95cce10e3996168ff90a650238c62cc1b3be973c2add8d2614406f3a2e446c7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f3d28870f5c1a1b10388ed966786b6804d2b21a3dca042ebc16470b9b00a1ec909805bc5a5bc83e07a5b56bedc05534efa137d2c2c4cd6bb0d7e1703bb87df2c8af6c4ae94d48949f9c24415f8d01de604cc880fbba3640dc18c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ab92ff03a24abf80fa58d8d1a4062edec198edbd2fee4c676a1210f6f44b58049a17fb20d2b749bc147f23873c3f373b9dae7025403b0e60d66fbe18372c6d28eb81f6fa7bb80309fcb191a696073cf88ba3dd65549a413fa4ecf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4957428517407d5f868ef963efc47368a63ff8449c9afc439f61192d0237aae4e35a7cc5c646a2dc2019e051fe72c9d709be74e8c37a7882d017881c08c57c03bdab9cc79af51be1b3b44961e0c5be7213510b01796c2a0a26eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b58fdc05d55e7dfb33f9d8166b3bee21422536bd7d6e22efa13377192755e473ae99519239e6b4667e778b94aa6851529b9667d4fc1d7f69c5b0e49bdd11176ae6f2dc6a87b2ca1e3fe7c67075707fca1939f3c134ae0c16a4bf4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc6db5ce61d5ae007082d5c415409d6da8d156132ddfec77d6ca92729d4e993f92a6d5cb5b771e013bc76123ac5d85e229cdf611b067eb824014b972c5f4952c9e5d31792eafbcbe452956acda395eeff0cc49658a6669aa4dd9a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48556471749c97b2b5e6574014ff434f141837fc4934a4688de43af4dbbd0c114d9f30f7d7a78b7a1a78ad551828104e1af4f1c0232e0677531709611ce71b1839493013177072dece4b0ef50cbb8ccfbcebcdb493c1d2e5b63c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6292fa611622b4c94bfcbb2353333cb0d3e2cd6c4f54fe7505ae19fb458aeb7a09222143007bfbbeafe739efb570cf2a1c71fd9961a43d651988997778a8fbc0cc1a4d8bdf3fd311bc9ca861a92092b31cdc2ebc304533b09911c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed81a267660a560da4e6df3ee6a0068677314434218d06a5b192b6a0e98bf4abb120d3842e11a0ab66376379e26907a8822d3a35c1480a49e6d2ab3a997e62cd00cf6ecfe22bbc8739ef6e9e9ade790b6451c85aa51737e29760fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e556a2fa75d70b4fe6e18f44a3afb1bb9c836b106bc60f6baf53720ead64fccfbfab704cd5fa43145537b56f091266c752a9c9f12c6c21c108fa18a4bbc2ab381228955994def9579e8a0ae801fe899170df171cbcf69941d3c8b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1384d3efd3ee4afbe132194e46fef17cc06a01aa6f32eec4660d0ac1d2d5c2745b95f42e2f0d1e5b6fc8c228aa6aade8f0fa5f7396014c6e9bc08fb9d5d7712ed87bd8639a0b7911c0bbf18106677fa3b0a036e0c639900999eab65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109df7492011fb19af7ab7ecfac7f858c65fcac9826cd43ac3e876531c80372249c9c9b08c1fe528e05b48d9e96720e35bd407d0b8a1f2f737bbc9d5a7592b959044f41bf1291585eb62b71d9a696884fcf4aa2544327bb28c59281;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16507e53457ac000383c9b567e5af28d642f540e77cd350a744ff45df64b72e2a4c988392258d5858311669b26224e0e5f2053b7c6ac2df0216204d862108fd855c4018445eab3808dc411db899503aa8d8cc05a1362a9c13facf97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha168d98cb0ec758eb7ef18d27fa07ff4e8b591c06d08d950e624cbaa406d58fb97da19934531d2c5738aa667a802c59a8420f7fb0b10650fb86ed4295277f071bb99957bf8259ffc200dddb0ac37274b39940168961ec867aca66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d168c35909ff09b7a1051002a9034f36f94e05c508aba692ba36dcf9f0aefc90a811e76bd8548e368efa099eed030dd8e7d19403d3c0aedbb03e8e009921310cb96b35d9773bc06ff01e7b9e8bd6bfaa2a523fe4502c7c0f435de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12fb175eeaeb4c5d57ef1819698ebe0b43790a6542fad77fd551493d2df77a46de1eaa175f6e330837ed6c49291c40c61bafff8bb93f75a08494e5d1a0381bd54b35b631f67158ab56fb9809139724d48167f964d38c2e29d2efeb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfcbbd4f9e3036183f4961fbbf14bafb27839b01070087f0e1cfab206ad055a258cd618ba8ebc10852522e5a8d6e5e0d7eb1a114823a848316b78a839c61d54f815f9dec06bf96321d290834a82d7662025fe4c3168ef8fc3cc4ba2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c1134bdcfe6fed71eb6f9e88d7c7003c861d84867655e28857ee631069ab1f6ba1611fa5cf75222a23eaca7994a538502474f2adc545cb62aec5a40b5e0ae6bf144441c880ea36b8e217a65cb2b70debb886e9095e4b54334a64c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1a17aaafa4779923a4f921968396ff86e9f39b6f9f0c86eb08ea94aa3c6032dd9bb118cd19d44af59be686d94a1d744732d85ace267b43047bdf97a06b3da4ff3fb6f638f2d97e9eaa4959dca6656f93fc8454f50ffe2fed8bfff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb129f89ad71349aaa43523ad5ec2549ad227767e48f2fa2a89eec95d768b530625a282e1e12904e68bfc194a7758cc9e40f037e9a6e51004d437b0f1158fd8f9fc52aa2aa31c1c12636623f0c5501010ac6e4b3365c6bc346b3168;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1166efafb9bb04d56df1fa6ec81e314c3279611cff8421d8e92d852991d2021426b004430eec90e1226007dc8bbb2989854063e8a7b5da71a42dfc416367f4e50103c89bf4b0067c661dd3e1bc260a02fb087aa1dadb750ce93a6e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58e32fa7fa931e10a05dea297a1c0c9fcf5e512d9a02b1cc684ac101ea384f222b683f13686211ce271c30d9128454d1ee2af2e9e19fb2d300a1f01813b838d3f574c967c20bf0cc30c974a151c29384c7fcf341e477f1254751d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h28f764f72df9eb96b62e193cf099e1400c4801dab64e9317ef26083a7b0687b5e3415e280f72d4072a69664f1793170ab418392c00ff756b31b776ebbe473846399efd815f73bbee434ee752773c1cd8b4fff8313d30d12f1b2303;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ac8c2a01b796a313f2b57e2d92ac9e03acaf2c52350c19231e8b0b452976c6dfc85778ac0034f9a005864cbd6cda53f6000344ebab19881a26f3b3548e54e5c02e74c1af574f5b4fce51dc1a866c6733b552850526cca4d2f3b68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1764974c3c7fee5fe1493fcc2fd4b09c7c97005e9c2f21b2974b38ee37a9d11b6541be259caeebfa502f54f0453e3a9357b22d3431e994a39f610d890729c632b4a89c93fdd7c0b759ba1c44a4338c73bb42e1051ee4f250ac56706;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd56688cc7fc0b067cf69ed85cef1d02f636a4c64a50ddb2e967df5c81b7911eef15990e7b301e15fc86c7594d5059cfafaaec17daf538f5ebaef39e7163b9ef635dcbbc50382ba77c64f3c4d990d8045b389dc7162a6bfa761e6c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a90d7e3b26fecda0e0fb1b4df4af04acc870ec6f4bded0ea70fe4682fe03d8d1bd45bbd0a48989ee33af1f3d5e2f0c94190df56a505078fbab8e3aa0868309662e77778675f1fbb1b792124ebb9b64f5c983fb243ac34f79b6060;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188cdd7f2ca6842d8646419d23de94f3b0087045b944e4031bf686fb6a1e291f1487260e9bfe9e490bc961e2e640ef06e089efde284e01ce5a16925ad12f508690d2407e8ba09a474627c8777526426fbe5df27397952a287e6822e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf32370d021c80a72570ecb689f6b2432f92a80d0eb89715da14cc103da6f453f16a02a4715ba33fd98e85a1299bacdda249ffff33c2e1e5d2bf478f2d368d6cdefcccc94c7e9179b42245943c611c4e6eef6780f36b2c8b5fc485;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ffbabc9ff74b2a771e2049292062d8381c2918ca4e884e94576be5e7a4750b70d5dcd9eb93fa7892aad1673f7fff16d780444a47078e857c438ed2fa7638849845975dfa3c8bd66e65cf7e6a99c1edc663adccab1ad396fd9041c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158f0df06cee699f230c3a9a15ece5bf081c083278692e2cffad96f09f9a2619d2cb1193356fc024df02ec4830fe06b3404ab7ab5e1c8b06a9492b54eb820e8a253b4ff9b00f10574cff06123bbdb0006fd1bb95a8df535da1ba98f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3df19d5bc68a993fe849a28017156bc833b96ca5f5042c9db1a51098c2b8c1b00169159271265d7bd3fb59fa6a8c76f9fd8760c3f479ced7e9b0702dd3987297cea8ae010e12c3f3a00eb8626c0e43f5ca2b9f96437ab72e301c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fcae4ed0720ad718eab0269c7fb976f640386bb7b300f469132bd9c1b0f55e156865f8a87ff14acc19672eaa60e8afd15fd5684d0e75077fed28a85c1330add4d4adf9569b4b9688ca9c8ecb9e654b9e5549a428e7d1624e84d14f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe18e5f16175bd0235c3e628454eccf04d4a699b47dd2fbe92a2dc8967d34df88d6a62d84a33f1058eadddd48ae3dba85a459b637e24b1c8a803b9b4a9be63601dd62e076fe85164e5814ca514c3b8b422d67bfcbdf90c29eaeafd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79c4e2900a5e2f1e658fdfa9b61c4f4a25b3d63e1c5e8a7a64a8623c4decaedaa6fe3842d2e74e17f23a43abba99e11108e9ae5899609e0a63ee1b05f65e4a5180c8f52528f0cde078579a1fe983e6eb72a99e6203b1f4e04c2218;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a4b7046be12879fb6664af1d41a6b1625efdf80ef54e0510670c18137185436976a341e4fcac3b840fdb06f0ddcad88f13083e3e035feef93bf29e0d132c32039256d6e4022ba4ac318744c2aff48b6d856109f294242e9d2ce5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1871d78ae6b02ec11899a739a434aeb9db5098d048c2ee849328ddf67da0d6ba88eef5b4d6002bf3327530366adcbc0911d3ad6b51ba54da587b23eb686eef22ec9ee33d637fc32ad99082f95563d85e43d9f577a23f02d8e965f3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1208f2675bca56708f48bcf4e301a07f75898382e081b6be7911aef40ce3ad64f007dcfeedab03f744eeb6a1b128abb7e3f66dc2d24b6acc494fcae46a984ede5c5a4201a7a97e8910b4d82773496819aad5d4362fda685c94b5185;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53b9a758a4950c208c9110cb811c69d17d78bf09809b14e8c818f0889daa123985bd12ce29d00c560ca5f8d1ce7772161c2b24772c27c0357335bdf4e9c659e3899e64db899d49b2ccd0036b8fb887e32a8a92c30e6606ecc28e96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h363bf6c82860e8d6261376f39f6dabb68f9ad3a72a3d28c09d17fa87c0dcdf17e66deb36c9f7ae5aaf5c90db6ed5e36b1ce8ee81e8aa0e4b12c24ec8f9157575d1bd4c0bbed58b1095a5f244aa71a7e70d5019cb114cb30683ac5a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d184f89c9c0d21f72021fbf598bebe98dac2a4abc236fcd93403caf62d4a66f86b443ebd0d22a245baf6b25749e4bbae59ddb68eea224a6cb9f9f26994f396cf75539453cf71404436e0446544867719527f4bfac21b83cf63b41a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcaaf1c2c67578936939eb7a5e14752cd7e041e0f12a93344f343b91821a27502b027fb396700a54bdf54a7c6315735ca6893fb40c0604f43775790d66c5e80027fe77d6844c32ac247735976aab0413de79d187e3f61b04f540612;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c719b6bf46e96e8bc840cdb451d0d76fb17b627820bceb1c20e62275f053cd5fd85878abb7b512220c85b87c2fba8bd94e8c302eb5dacd500e2540905d71ed27f293c3644552a4d1e036f1bc9dd9404d3412048f101925fca77d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4c19dc88e6ee5a301644c05a5b7e30fe2002c3cea65e466fafcae059f755ab4bac6315e6fe7ece74df60d237242ad92efe7b15b85305180bb698df4e28ab9ae938991c7ede6c926e884deb1ac1beffe7d97da041fe325cb547fb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102beea40d23eec644283f850a01d7c9a460d71300be310a2df588a2ec8a0c1c4c04387dcd204e88b166b636fb71262c42a686058add2f3d940cbfe30d29d763853c77853c08c6ca65b4a50b94878cd03a4031583639f6c5528aac8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6c3280bb3ec8cf1758d55a2d5e0338bbdc27f937aa5993e3b15e3c7ad13eaa2b6e739b5e9031f839933f810162a9dce4bcfb584773bb8c29ad0d486845acda6e2d2d61ffa68a27495efc3445a17f62c5b2f29880bef38a1f876f7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb8e4c68718795b9f31a8a26f0637d85aaa02273a57e7c5379ba858be56c8e89feeab537afa42047d5f89745acd85652c50bafb2e438f33894ec7b96ab90f169e09bdf3d42d16c0951fbc4a999c47754714f9068b80cb47d630e91;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5baac7702d13378786a1cba52100723573d3dda988783fdc06bd69c34851249929891f0dc6b0742faf19f29d12f0929ed2395694a470446271c4e4a0de2c0b6549a9a42256daa810a756693dd25d80448811ad9fd6c6d69c25af66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137ce02d1234f2ed89b9eb4bb9791f67430ac3fa3274745c19d065e4c48a912c720f7844b3ea70f0d3716f4f33ada97b1069678c3ae5be10fae31c63ba1f69315ac6ca8894363fd3b97d5a6426b632b49989b142bbb62d95da1c1ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2d6cc1c95d4feab960a355456aa8fa4498e1e42a9122c77cf4afa3a40e8731249805331b79dccdbff4944d7572d14682d82cd6931c15c85db740307da330b695eb5d4004116a22f905c1f369c71ae55e9d8120ee39006fb733ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ab4acba1832a5ad42dadd7601b00abd045a6d27fbed2f787e4a22db6c42d6f6c963f7cfdca21952e22744ff866c115debeda59f4bd190bf13efd2b03b2cbdf799bc86eac14e93bd44441817cd94219009c70ee26b8625b5ee23a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130cc6795bd81d5065fcf0edf66b862985f9ec179b42c1cb2d62f9c3cb69a2dc9e913d3a0d5fa4e7008c4ca7dffea8ad2f7f5496f7fc8cbe2e6676974ef9695d31c3f0bde11f80bc5012206dff6f2e331141b432c1a81d6f526e755;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a7045a197f23e0c7588b17c84feb1026ce744bf33feb7d72601b46c243376517fe98813f41e90a716e4c42beabcbae28d279a09234968f6d6153c95c5d1148f9e5b249969d4053ae7b25c15bf07dbe571971fc2ec82ac180e2c6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c60098f9e5e34b2cecb4061104bad6446d083d2927690e00421b224282f85d711ee44219a6adb9679c07506faf6d191100acdfc83ce5c0441df93a4bc057f6fa3cbae0f95ee9b3236c8dc938616ec91c15c303d8b710f002b1611;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc55a9fd2fcbc2d4900921efc9440ae2382379f123723f46b6adb356253b509dfaa91fbe0b49c3fe6a8d5aa52e36becab0e836fd7ed9e4691665c67b02d88c5c795500d7965e61033c17b1f50c85488b4cc1cfd9e9c8ecf87c16d82;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191f317fc44b1bf78905dc5212206525f7c11f26f21896da20d24b25fabc9eef5c3309defb9b2cb9d44b5a1200dcbb0060c66a535d09cc903c56dd95cd57818de258d677aaef7faf8e23733777ce6c3fb1ff10039b328f73cf1bd47;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168994c07ea02c5ca26d1a133151fcf94e8cf86da831e7215104f15f21624ca360298125066823e4d41faf04b9f3a96f9211f4b977b921000727e64935a12f1027ece4e589f3b0d87fc1d56c6bbaaf1f0e04bcaf04e2584e700bce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd4e2e911da0a4560287aaf95c96b9b23f28181b3cf214e30834078b2d03576849388a640d15447fd34ea3cac0c766361a04b984efced2b8914cc03ce8375787a8728800a5d39477743b4d46720ff3b790f55212a58c314bf61a1e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8464e0bae5c565cd3d3acdb0bc3679871ed6968c9592b45209c686b85258c30835a82e154eb99f90a9607027ca729999fd68cd27a90d4bd4a1cffd6154ff59ad4ba1a359b26fa0278bf2ffe21e02be1c1b33a5bac9c5aa03b633d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfa78e496ba394c6cf01a6e2943d545d2ab406b81fc2e6489e8d12b3ad9c21fd02148da38b3c4ac505e6891ac5a482dccbc43c97b108a04015102682e4ae78dd2bd92d8dc7c6b55ab45808faf35b5a8a2742a1663bbbf016944890;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1431298e5123437f9189b415977a245188be5c368904bd7795ce9c5adf64f8fa0728d25d8c067786d367f2c184cd89fef91cd520dfad759e3c6bbb9de5e6b8dceec326a3700ba170e9ebba7dc7641b2475407da4b77bdf325a3a555;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110b460554adb29cbd1d1887c7112986d9cef8071d01fa1e2cb060418460f0b4ba565e22a22793821844abec9d50b8f4e4182ce1e64606ec6cf31f6f892b0792244614ef85b5cd4f34ca25a61a53bf9dd847e5c2d4a9a1b78d757f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecee090e72dc149d0252fb0985e265ff37167e2d858a77f83e6a26879d6ac88479f4dd9fba4ad96da25d4be491a52332b5acac6a81d26145c96a7e74932a991a9c25787a826690905865112c86d8be70b6f971f550ad166f063433;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106ad691aef279c64d544608774ebb34365e8d11d0886b4a7e61770553ebe9c589c132da812510abadd25034b710f75c732b388284ded8bc8773be6da339332911d3322c2bdf5fe3e152f2751521d636ea6bb837ffcc63d9af41816;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72d88c4f80a81b5a2bf89dc0f28a34751455b6192e519e703fdbbc19632bad2d0ed6d1921368fec5c8075b32017049db58c3791bee745159cc7f3cb2f6ddb7e484069a7fe6e444e5f0d6c15a8e70ae570e6dd55afe7f404f043c27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he76bf13b300c38e9029403dc45dc5e34d470afbbc3178dc441e080d86176cb48466c068a78380c766b6129c978bccfaebf81068e2932694b23b4599bc32f0bd748299742ff22e01e05b5b1bd80382ffb9ab557b0527398638d211e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c55ea198d7c7048c7a060e54a41fe80aafd188111cd21cdb59fb13531965b4b18ceb0347031a66e826e62162e71e672c0829decdd18b6e4217b2aa679d66d6dce330c8848938ad21f38841a48a9ae90eb8d7e56d18acbb513cb208;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4a919dacd67ca610fb77236d009131e813dda56c2a502034b27c5b68f530a46e4a7781d98020a3870ae32aa4c432aef00174fedf39bfd3213f47cc8f578401df9ea9b594f2f2934cc273ed93b2551d70c1c9b70550e93db019a1b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78c5f66937c57d84044c8291560281a952946b0fa1758e549cbb7bca358625d9cddee4bc76a59ec635c817fa68e79c379a95d4572a236b2d3995aa5dde827533b8e4aafa727ec0c4296c438ffae72e9ff5cbd070d9bf90a1820857;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h346a5e27c216dd622493d59755aaba582fd5e0fb632664a011b32a324da8ad270991344f4f23cfee1a27bae0c0edbfdac6408fe156b35ddd91ff49df6a96e4982f654a4d8f7a3f381ec9226c1bd0493fcc5da6c38fa86f9f3394ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e016902524183de295b3e7da9914f399df5b2b2983c53e35655cce52111d274a2606d2e2aea7500044d142c35900a040f68a73ec726d1372f9c16e076d742d5817030717431a39bf1f8c3a35256a5f603b46c4a4712b9f006e03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96fe72d145a57cd41d7683b67cc90199d270f97154ca49673e79a9d9c0d8a5b0034ef43f4fa1efca716307a8d1d3764237f32bfeee8fca846adb253b23492e61d6735a40e5e9aa097af8e1d60f1d2cecc9e7cb83dafec402966a2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199342dac79b65c4a28d4428fd0ffcf0ce556766f2d691298abef0875589f2635c2f695ba5bbd55e61a91419b59ea599d1d5e27c2fc0e8dd7f36f27fd774c26a183e14d521988a7c5571b186be03f50522ecd3037f554f7f26d40d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3d1ecb8a2a6dfcdfd706d0d2bd606b5d7206fa90ef85f1a0fdc0398dcf1efd97f389598297a67bb897967454d4f1f73a3020ac097b9e93bc90a3d110f392b22ab60eeb1a0894ee4a906895ca15198441821272a7bd48db1357be2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14044fe2834a994709a3e0c7c8657d42781766501e16817f37b26943e8cd0ab5433ce766c210b245defac6eb19a29c5a382c639467bb3b77b43a72cf366f0cb2a0a361053e6e88ad4402bdd2e2008fd5b6b38723d8b144376ccc60e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184e58ca128706d22aec21eb58df61c7086976074f442d2b8a8142d92af8b4e679b3fb026f97927f3e6357d9705111e56f6bf59eb734da01c09ed85c889eb44bf98925630ef3ac29d582ec4db5bf934ae79528c58f28f3366d09921;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13daf2fc76452c978467211195595f898e1933c18482360d990cea2e1d625262c13d756adc67d7e23dc91f891f4e4c07e23458cb3c2c9c7fee246ab3a217ab948a20c7ab1031fde7c1b2ce0e8523f6f0d2aeac611a4a63000554014;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h329db1cd1d331c94e39dd5794db18240dfcd5052d42c19615c738353363e8bdc4c4607ddd732a18cd317065db2ea0b3803d9e5503a53a0191fbed9142251458c3aeafaffd5d74fc776fe33d20a0aaba9cdf1ea5eff737d074ad80e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc276b75d9c75168d5eadc6cc6ded3456b3c151a34f8adcb36471500d046552c55ce485596c18ceb2363bb48dba65c05ef1a3688a9cbaaabdf03768895ced27861cb086ddb7bb6eedcf9d7c5547f35fd94b4dbccd865f6cdc252a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3abffd0a8b73d7d56a50a85674d2ff7ba0fb5a33625bfff99e99467ad235092d165397d06ad0e593a726022d5e285cb6131352b0e4f48e8e270e31d714ea2881326a85eaa8a7eb6b0b2157f0bbfd0c7e8c3a80c7b432807d78717;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a000e07056d02d7136d7565154bc5ea863e9e012622bb5b580c18cd0ac2d80bcd6276bbbdb7672c9ed4a2200bd6f9673492a89e86a8190d65b73e8001920d00b95cfaf0cf97d2e5d3d8cd32beff644bdea3261db1d35f33b89e2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18741090eda418ba8caaa1330c86eb65fd5772976d31540a1a14d83d23450416b56a9e803b64cdf60c40f51ea2f045cd0ffb01a9cc243a3ca47ecf64fa48c1d71a8a7560f74e37340f585341eed5ea3fa38fb808f9937e9cbefad56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa7670dbb2e344d25db43904840ebedc58997a4cccbbdb6f685ecc1743d5274932c17d52b05637c7db5cdd677d3ac0797eaebaa0046cb2ace2b0558b97483c9499b355add6f8f4f89e72a404c31443f1b61d70837b66079a88f23a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h433a7db18ff8d361bbd8367af9cf2e57ef24b964237bcfd152014d60e88f8b6451f92389ed9192eb6f71768e7609f61a885e12155944be0ecbdd7b347ffb6463d2c9bb90264038788cec4833decc32ca7f284b19d91339a045ebc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h671532dab2b29f709cfbb02f9cf1ef6ff8293e388dae6b363b6e94efa5dc7dd29ce2eca62d218bc5715de29339edce0bdf52d4c192aa991075324f44d536ed5ba27a459358e7e080dbd11203d450e03bae9c7f371b4d6d23bf05d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1432b46f1659f92f9530db809e9fb9328c86c92369a0ad3ab19f5baa48291c5b95537b152450c347b52d4c98111da803e62ce01c991ec057a5015dbda3dfd53d9fcfeffeb4168307aaef9197c77fb533dbecbb317ba250de3121308;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a4859c5d74e444b283452dedceec9bb90a4f28330a5bf9e6844f7a6eb8448c9e561ecc7bee98c6cc18c1000fdc20496d9b2fedfd7a90a2e688356a8c201b9926a42991f65c4a202361931c429f56df23858b34def912faba4ba69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9615d7f44e133b8c594b10123ffbcc69612c047cd45b59fc45ea3618c4db6b56e721650bf17a86e8cdc07b745869a9d83fb4ba107ab5445d0bc7b6598126ea3ffdbb5d5ba9d1f750f46d4f46a28a1513194500dff5f5cac708db45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h305a10f0602b7c0270f2e996c6059f13c1f9f31a4ca4e198c2ae9313efefa74ef8483da640b0a850adce804e9a97e93da8391562805c372bc9a98746acf1120d3b323906b097bbde0d33c4e7c98b2498c75744b2def7a605033781;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b3df41fe072cd4b9659097b2b7b8106f0418671dc9423b586af731e1344df0daa893dc6139eb28a67d4f1ed03ebe537ef044e9fa7d30a6612e20850aa0efa16c90584e027d8887aa05dd8d2e96a91ab82b849d2a8e73cad7510b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e4e01891a489e50c504092ab2509717ab598319c0cb412f9848e45e7d46ab8e6c086d94e0ca0a16f523b18e9eab562088ef772ee160ad5adf87abf46dd664825f2c8a2cf3cbfb6b37a2f3113d76cb6262e571b7471439ab3dcbd8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd4c7888ee73a11af5c982e96d042b48a7ea05855b736f2a962a2b5969f2f4efc7edebd07f88e2ea7777033399bcafbf1105cb37ba20a6c27009475619b238dc06fbfb2885eb636215c4162b5a49eff450d4bf384c435ecd1f0266b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1098477c5d1c11355bf97a4aef7e63ccf13730a9b0692beee4373bff60331e72b4f6dbffa3645bb09b1ff8008f12ca8a6c5641ecbf39fd98995c9833ebe939e0ec2f4efe1b13732fc4b0b745c5e8a896f73594da0bf96372b71cf16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f48be21d9588fa2274c9efe0401eac56a9a9e02ae1f456f6b0f06c1424c746037ad7153277b12c6776d4f935b2cb47976fa772750f3f58effe0c97e6baea559b2a96ffc4cf92b9b02f2f609c13e8ad95e1d90da7034ef0c30e17c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed9756774e08a219797f37eae76576356a977043075cd6f51ba35b1fa9ba16ea6891dac596194caf456bf47d06f893b84f6fab0e70029f35b4f451f1d1dc824816958b5717c7d51d676afcac37ff1efa1a7129d1ed30816f863622;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97243bdbf25e88a37469a9a21aefb5e39a41a86dea90ab1b4d7fcc88e6c4e221cc133f417b4bd1108e9adc85ca0c49c8ba3b4f3c8153e30a687399465ea1c446cf3f89bae5ac0207f409bd8f144b2714dd7959bc8d60eed92c5eb9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h485e17f2d48b253df180fe068461f2c73091a554be90bdd831e14ebb4f92264245722d2ffb3db9e8d94e5583244f8a0ea2f1c22fa99669e1288247e0ff6f0bc10925e72cab73751940503a9aee641ca519a7be28a937748ae58a16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67530d034eb709457734fe4de453b805a4d66c4cd6ce83bd64676bbc35d24a5b0dbe9271388e9fe23e46f6c416355f7df706233e7506dbdfa42e24094690ff0b321a7d5a357210a26e214c13f2da6525e6e1aa54d2b72f6fbb9d7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f0e9564afa3c940279b5b641d9cb9eceb74bbd8ae4aa9290ad5ad189b43b2c4e8b41a24c511fbb7f7815c4534734f7f95cd9598d3b0dce1ab85fc40284836e59538ee6220a8c21b0ace50b21898d8e81a2c74bf3a60cc13a17406;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1b8c5d554876a55c7e6b9ab25c30f84b9ca0942686bc3cddc5b2a6434c0fe58b670d8828bbb6bb37c061e6082da08ddec6cc799a1d51bd56ceab1eadc605176ad21512129ac9e9b2492b02858e8f728a52958751d0d3339ee6008;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3f57e2559f6afe33745e4236cdd650fcbf9e685628ceafa156ecc7aa27c6a841d2ec3ed6384e7d7884f6826b4a8a42aa683d33fc2e8210ab097f562e68f743c7ac338a25d51ba423f0fa8c9d0c039ea45b93e80a4e41ffd4362e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18da20c4d40870d2ef42120abdebbc2f794c454a3d57424495d74621a4e03fdec5135fe999fa963b4774af3f06a0ca8b192d1ca73e0911b37765bc95529073a11ad4644a4a914a26bf3db9def465a2b2ad9ee17ee093361101a301d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a09ad810226a86ea5628d74afa0c2c428ef2aa7ab31a489e3ca0bedb175828671a3a8000b91f85a503673adb4e3c0759fc39dd16dc8f55a03df70449f3337bdb34389a68a4e54802b4f22e32ffa05bcd4ce0bdad997cc628c3bd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3a8ed1e0c5c8495af62003dbcf0341510096992d6e208ad12c4b789c13802ebc10eb1f8697a698f016eb900df7716d40e3d1b0a9de1076caa6fa47298cf77eb0920a977102350a7889dde7d53192e1c86288d30f808caf769c9f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc88ffc5ba3bfb6ad5ac079b30adc54b980d10bce75b8eb2f37fe98589216f7a3ba62115f122939e5cbb57c4aeb752bb94f2a5f041494cca28a1272c61e13f75997fd357402f20a046118305013cc8d6a3e9b7e507267c1e8c95d9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125f9e0d5601e12e2743b28f0b3391ceb9aeedfcef9d3289fcd92fc7cd40dc516ef4e25b11a7a6b5b6da38800bf030ed98fe6d30c9f2c4441625b3dba6808f1a7aeb3c47d6b989ea80c2c09c870e08039ae8ec5bd244d222126ed5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ffc3dc9cde47fbd77283c4d9c391b9594f76392be3dc57452c688fba87d86cb2e192e4b9fc4a01c9f4eb9eb7030785c4bd9a7146214f5c34cad7ccd5a5fb403868ab746c12c5a3c56e25f819e65514724eb956f1b8410ca2095b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1baf325c733f4276814d1c27b37fa2770c8cf0ca573ea4770f348c867bfc9d16b8426f72a82ef8cfec235e09a5e45e1a7deeaf990b253db8aa5968669db65209d42d0f5ae44b9706b7f668df62330cfb34dc8050aa5f39236351f73;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185a501e7c7f813ef83104cb9303b2776d9256ac10ecc473b7a27586e0410b3c3b97309f35c27e9ce954005046c9408beb3a79e0f716a2a5c2776e1b0994d56fdbce526432d8edae09b9a6c7afd4cd6f902384d4dbc7d4a09fbf15f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3bdce2d6f46d83d60731813463721085e4ff0bd43ed957f4e0ee4a6adb71ec7ded8d81ebc76c03c690935e70d6d06c381e26e95805d247f60c8ea1cb1be7100cdcfaffaa630fa85d8e494001ce5f4b95743c0073192519bd2e17d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h108466301824e16d41f2f021e4bc4728a55b78375ed51ba9e4e055fd809d38e9cd998afcb4e9f86230468fc52a3eb861c5799d4a740c62c3bcc1f32c2fb59fd37643d102a766f456b8b7533a5f67332486d21698335c05053b1d42e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f90fbf08b058307e16d7fbed924a67761b7819070281898a3eb88ecbbc1cb58362a58bbd34ffb7e33f499df2e5a65e7ec2a84e8f9f52d9e0e0f5a7c05a634c7371c8d22f9f532cf25893bd651c7b06d9614b15dfd6a91d5e04f86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbec4f9362eaef77791746ff7820a07336b26ba2f955bfba5bac59792787e05495c35b7b5387bf3b0f48723b0c65d9e9cde5accae6dda41f9f42b6cbd3662a12bf7493463bb0bcccdbfe7301e0a5ca6519ea6454fc66f48c19cafb0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4356c888f63dba3f6982fa40d67d8c9182c41b5b4fd048e63ba4ecaa27d11738849fb63458cd85dbe449a00b14098197effe3a85dcc73021ada5fe506f928bb6be21f755d82b7c0c85fb37cba993392c9aec85c176027d741cf88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1372ec5ef9c6284eed741b32a30978d9b2881318c98c1dfbc1c4eab2392f17678aad8592c6af2631cb1ea9e4a8c30c71b629c941cab7907fd2e0f7b498affd9f3a06b0bdd4153f4cfeea59797ce414b9fbf31e73ab88d0c34eb5ca2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d0e61dc18ead41e5ce1f950e061bb741e897c7524401dc720196c511273f839d300a35cd58491d416b90cca69b75b18a642b55068e439abd0629d748febedc48a2b71cd5f4ab2be822d1dd9e01f2706132ab21a5649bead8f6ada;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha21b68c9406aa30f5718dc98f85aacb244797437135724cd9be112caee3f4033c7d6b7d44d7160fda5c5af67ef3a8e934ed550ce64377c130ba9609cac47fedbdb53a0889cab2db584950200e9f94d646d30f0c98a452f755e9356;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0ca23cfeac9b15033ab2017112efe72c42afbe993fc7b39ab322912a5d30c5d2a1dafab7ea0e01d9dd1f7b2df828fa65bb03a375f6a76a579d8ded49832f027202d4707579ee4472b71908360386598fd7a6083cb4bdcea5c3741;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127b40cbe76763f65903d4bd2193c4fd68e6548524d476d58c5de2db655dffd474c4be18246f13e912a05890143eb477cd9d378f911a903f5dbdca33a92c19ef0e42f61e8333d69a7ca097a7bce193e63f5679cbce48db64c11da81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101cc3480d14e2e550fb074ed0ffd6b78be8250e73bf1aa8ba6f5c90ba11345de1426a3427f70523310a967ee87ea47a5a0ba769466ad54310ac914e0f3f2bc9384e4a0f1088980693c6741f3394a607d619f24dcd3f8c538f332fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1179ddf3539c91736afd26d215b378d1438f78a0fa4bae7c8584165d838cc97fbd7dd46666779d65df1a46df32fa50fb6a32ed72c8305d85f7c85cb448603206cf97df20229de4584903dcf31fd65e23df1991c4df53a16c2f2701f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b17fd75e739e7b32f0174a3245b82b4d7f78e746903bede44a8e650fe577b27ccc3c7933c3f84f20b265b5a035bb6a99ff09b7473d95cacc73b2d3a15a33d31cc62043a130f4d9b6a4f8bde5120693250c4e32e8abf0bee0adee5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a77ff11bd4d13afe0a9439abe61a99e8e944b390d8d0735774b5bdc7b0185f097c8dcb624e2728e51d2ac59585f1cbae95e0516e082445f74e555622f9c9168aea2d8e907751f2f177dffe1e86f35ae961c719a28c1f3649d15b52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ff4e7ef766ddc36236b0ca9298d2d77e0643c9c0a45a232739fd93d01a908a155b3bcb7f086bef6f410f55a7c931a88177e436d0a2ba9264e3fe9df46bd7397f5845b167c2de4957ffa15bb63c88ef73c3f02ffaf1fa0ee9d7efe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16df7ff25aafff0e63d51d84278dbbadbe54dd5ade5dd32a0cd7c184f99c77cecb1922d165dd2bae3a9a04e1ead6875eb893465ecc9d7d560f3a515a5b6eb036e2e1fd5597d3590e7a97a7ad4a461f9e6372820cd72546348857a65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7e1455f3014a6f00b8eb59bdcaca96cf45221e5772261ff1e66ab3c30d4d33ab1f9a9dcce2e1f756bfed47cc727def4b46a24ea0a7902a59ea7f7638109ab86e05ca4f6094096231d04689f9a29e31a82e071debd2e18d7bb1736;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c14089a2977b7403dcc28d44170205b80c6bf590dcb32801fd9ddea6affa9255fe9cc35b375fb2e7f076400a9358f3c9a47862e2727046dfcbefaf5ab15386b30f1ce7b0da1cd935f67f021360b4e6713dec8486765973ea2b29f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed4b8d518826b1929060ba6ebf1f3ff1d585677586e9d246fcc8faf30537007dc27a1ea194a7471c570808be05308a7dba6f13bce11c0515186e3012956ce6f3537a5c08f62a18f08ae6d67553d3e2f1c3904cf8159e7b3457280a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef5f1ea8fa64b8caf48bc520e91f5bd912ef0d263d5986da02ad2c7a0621ece5a1f3b453e7a849626cf4e21ba0eb2189d09961a1e5df9e65c604aa9afd4aa3aa8f704f9eb9eafdd6d62cb7319c1973c1daab4585a386e93678a4b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e3eabbf50662b76557aeca62a6555af2f4fb7e9e456b6856eb1eea70e1cbc3948004725ccec031f8416ffb75be32e3ec993ddf08eb6a5e0390c1996c00b4a64ec8a3d064addc13d1f5dd236399822415d3c967069ddb95aac2085;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10190a707cdf555d0af410e6951d5d1d199f8a6dca77a9dee5dda886bf262032436627520131310cbe93002537af21da27f0f5827d6a73c546323cc43f69be5565912650160bd6f34500b3aea7a86f54b7ab3b4667a5751192006e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dd5ea623f919a1994658f231bfe92d16ac411c0e2dfca83f68e141d62f7ecfe69fbda6ef6d798ce036c7e46b1bcdb4c34c1cfbe6f278fe56f9121844850a30a1b1b97cafd38e83e8ca04a7467b1b6e41bb5a2c1e817bfc2b4bc552;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64fa0a11367f97ef17581e6c4b55a2423fbd0418401635127547b8502be080d22235b539df8c073719a6866639c052f67abc729dcd67dff63e16e7bb360f55d843d13de209b70cde2768646bde9bfcd1cfef45a2e2481fa44c17af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ea00ae120eccd819999424c55d2356fc9b032f8e8aff46000ab123b3f8f7d776132a6db25b328e6e363f27b0b6e715f62336bd0bd819b1ee87adeee29d0ef36cef6f55e09a12b1dcc8fe333168eb53aa63cdebfad68d8823f02ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h238db74d6fd504c4bbc066a17d3d614d7c45cc2717b5a9d3cdb9bcbd26f4d6236dfa314d46795f488854ebd5c18617d1f7dfc0b450cf98505d9ed95ae35b3ad3cdf7ef16095436500d03c249f77b72404f2adac86342f0a99aaa60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfe10fbed3364111b3ecfb053b490f178e3de14ab5fb988a97d2300fb3ee22a1bcefae56558715be239f4ab02503a6205f7757f4a29c0353590ecf30eb46c4bc5b516bc5bc97acff487e47a683234ba4fa27d05747ed7c8db42b51;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24e4a144d5e5f4852f0b366d4d70021c6e608d0e50b9fb216ad87b8efdb472cc206393e26a1261a1f6db80475a7d531a40b53b334768d48e7db8457d016fb6e74f808c2b966e289d8b8731320aa56fa1fd414e718ca8493ee62b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d7f96e1084d698849c5735417a2b920be3affc25edd1a03bbe4ead09adf1186c87e1e80c9a4e7005f86e33dc49c1a6126415f6be23dc8c23bf9049623a790cb56ad4c7d41cce99f4ef800bb4b823ba9e01c7c486abfa0c5ccb30f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1979e12808296b4d1b8abb915740bfe2f5a13bfda62e5650cc8b70ede62b415167c137aa1466d56dcc3bcc687aa4479c7a54e1e94d39e5a0cb65d19a22ea65d16961b4d1ff7505ae016c22e93197002c1778dbfc5b381257c3dad84;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b3039bdb6dd15054fd26aa494e82db34f0de7650847cf62fca8273c10c6b4bc134cb09009b374b8a0a70f1a76513f092c98048965dccb710078a574f544ab7a38336d51bfafc54ec46ecf7aa827e25b9007da78b902c4cd52b8ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8cbc2f8c0750963a8104a78f6b3c6750bb6c05a39974c5746f8f26d677acc7d4789468f84e634329da2583c0da5d5c927171db238f4a698a845b896b5c3e3f782b834029e776eb3899a7901b8b3f2ea75f0b913368cb006eff9e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca980bfd2b34175b9f023fdc67c62a4be509a9e371257a44c144c10cf041b814dd3a97f4bb9fdcdcae6fbab0f4f5b91c14ef4af4cbc0d7dcf13eaf1e88fbe71432c30192595dfe8c2722d96043c61a060266bf84879c938b42461c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce75684170bb351940d2c97a5cf1517d633d181ed5caf7d5b5aa2940911748c1b8fdfcc99d7edbcd427212d361c1fc536d377bb6c21c9893e7058a31fa6a031fae4c0ed11cc5960f894e1cd1f9f906384493484c010f53fdb896c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1edef69b54ded6d8cbf2e6eec0b73fcea2ccba696ca9f525068a34980e5349e3c3a32863e47bc63b1ce54dca3a29b21a586e2145e0cbb78ef968f17ef7d973e7a34c3105a497366847da4ba0bd469a7f7959b72e2dad884e8cdc0c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e3c336cd3d77b6933d459bc2c9a68630e9364d74a84c308e9ff28f394b0c783e488003903944a4100cc2f8b1aa04d2c7132a28b96625ea2b8cc79a920ae54fd26cc60b3bd53ca81f546f2a656c6476c94eb930af1366d28ffb00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114a2e63141db8358d621ac7d8dd9cebd36ec404a00881975b51862e2cc6fdffec961feed9bfa618860ec05bcce56fc26e4568f41bf456271ba07e261197454b0a1862e8b49138a56396bf2195194db7148e0ccb55fe208e707d78d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bdcc22d95bffc7a309c879a59178f637f145dc01429ad7957b9612d01d8028a0a7f38f601623271ce22a075d47dfaa333b5e88b5288c437192b00a82b5cef4980fd7785ff1f35a52fd990ecdfabb1c280b017b961ba7b77b0f0ad6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f73f71d12c70b409f403d0ad73e6c823394a204de903f9cd52efabe4fd23f5df952146b999c3e20cafc3110d73e53b250acb76b5a098d81b4866c9229847b64241185360f73fd52cfadf84bfd553d218e581737f5183562e752b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2228055ad8b15b7088134b2cf42395443e12c81653ce6c8e324ebc63cf11e8c2b0b8e71cce16a3b6caa9c3b22cc41eaf8d98e5b9968a85101ae880ff7d63735801616cc419d850966d2a3cd248e04646bf6fb5a5c245e5752e8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e7e34ae5a9054f8ae7f6171cf38b8823f1a1cf0a3c4c8ae41e99d850f6b00cef85743f3e1bec16ece13de974d74a427c1b6975457fd269d62e42f8010029700599a36a8bd487536d32ca6687b047159ad7bba3ef3be856ecf6f77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h871ca317cdd88b79711e9b5957a43f55086e14e22fd66b0ce9f0aa211915356e77488b0d362e7cfa410cdbe04df4466cb892958df657ae7005ced721b68db81d5bdca85eedf3d6603667d94f521308e0a3f853eee058ffb3a14f2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4f45fb04216b9e5e73ebed6aa0b090a75f559a9f7fce9a272dd960db606aa0faf7d22d00ad75de44101834c8d95a648a6fb14c9d11eb5689ff5b74efa04c89f64ff90cb3873338299254af3f4c0311709c44428cf5eebf333fa88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee55b9c2d4811b6ac28eefa27fa026daaa0d19a6ea91d1db8f50975469a0dbf4410650d1c51bb292a951d19104d3ef1cec329a4adfa22de3ec83336bdfbb09bb3828693a9214adfdc290c2591e8b72387721325c1269e27b0e9a9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cd51412524d01b9aa1d6fc169663c938a30a0ff7e20a2a26b83c37620a92f79292faf6c3fe27953894d136513621b76dc8180f48bc88e426681f32c2efed2b5bad0cdf957804012218effcdae0380730903580701772cf15a5ca3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fbaf9f19002de1b42bc2ebffaf7f59e7f840ea9f494ead869416900db7e7b05c73e8997aa7eccc01db9ce4ff158d6f0803c61c4edae69cb8ce4c037122cbea591d966f47f265e5c576c573022f89ef01d2d40adea97e73e99d855;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f86c16f1845556cdcf4a722796fca90f1b4cfd2f42030f4799027ff2865ccc0a0b776e34f784827b94f5922c4c4fd87a74218fba07d17ead9c19d0fc45aa204477e826e4bde6c3667de0b1dacf7cfe9f8283f9951c9d197784cc6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hff3e2b7355d32558a409e17700d1ddf0000c9c1c34ae9b9766143227815483d2d78793bda7b00887621f022aeed3fe98993ffed8a07cb46b36aef10d21669b66d73425064e2888c84b27688d9a6e7eef08a674806acc5a34e84e20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43815646d16747706592803a7737afdc681d59aa943389a5beb093b3c07c6f4a0969e03186fe319976c36a6402c74aaac8a97e30f04f9f2416d90edee027f6db54a0df3fc63c5cadae90963226cdb3a7ac2fde404cf0ca2d14fc6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98bffbad00821f43efd23189d850c44b708356a3bf9c47157ca97e6e776908a574b7e256e7fad4ffa92caec9fa41a663121d223b39dfeb877319a27306f4fa53041bfcf3c7b51a6b0e2ef80ce37f36e2770e00c57115a7089bfe7e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h577be4842f3f69268e31e807b96eb68c19a8b2f2e791b65b4a5efa42bea279ce717dd0ecd112be30703ecb8ed9d9859032c29ebca9a5a585edc87137e819fd19a23cbbf447155b069e6dce758d9814602c8cfa55bdf23e21b8a1cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133ef401b6b74a7fe87d49349478bd4a25af7c8d7b6ba0e3a2da8437b70c04a7fc59af640973a6995917ed0e1cb11c389e93d841e81f331bd4e038f09afd89d307afd1648104a04f4eb542ed5ed97f1846a5432fcc492ffb5bf3f73;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd1ffe86442f370e0a9b1847eb82e824746d49d57917d8a47f1d45c5751315b0628672d5e88332543e6f00c092d101868625065b004601243fcbb523ab621f1474d206ea1fa6030e363c3ca01f3e0089e4fa8176fe9c80f0e44412;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16dfd0f39e266b0fe65fd50d4e21b841a9423adee0f0c2ed2e242962a9f6d63bc3e2d12cbe3674411a3bf658e8e25b0773e3e993b158026015b00787046b98c2260f5044d448f4886f7fd618c3c7a3ef639a051aae6919c5754484e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ce59920e12f74a6b06dace1cb9ccfffbe8337252738dde2e5e9e7aa9bc0c44f39efd8b77b6a00f8ffb001ddbc8c67629e3d91290adff19aeff52f20a3ca0a2f52a333b040e7c4ef1f6ef8b815cfeaf541bbd44f342d1ac903a89d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e9ccb955ab4b0289a66f76641a24db8887e23598044d8cea1889b9cd9e67094013234377d0ec4dc7beb549be9725dfbaab0c0a99ba5d4424b0513c8af8673be62d27e044a62ecf127ee6059ad0497b42edc695c4508b056f8ab95;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41c82a522559036b99997ed3b20cd6d17800c9be351f3ea1a16398257de20d0dc71e3c97e28ffad4f29afd0ce466661937e08214f701d3410f26adcc45fd81eb8da12c6b6f17cb2024e986043d4e51ca2e5bc2c6673f9b70912950;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d41e7f181c02f41f5c155065093741f208fe889e3b8353a879e1731b1f42c4659d831e830f788399965072a9a778ebb7eff3ef816931505932d042bfe82549184b19f4eb1df573c0cde8bc956549ad495d53a70a0aeaf1ee6974c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fa020b3c263887c94b57e6b89950143eea7585892fc22c0dd9ff095353b7e044feb6e597fa41408e801a9ec1291bd16624a45ccf9372d5bc9c74312afecf6c1f6fa5f65d28bdcb8411ba4f26ef101104540a4ac82b2f5810f4825;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ea7f4252bceef2fc9d4468d53c9e5fa0413095c24cec6d82afd508c0e1cf8064ead5316beb3a6eff71ab7748eddd4258cb92bb4a6c5cb3c95f2c38d246f588cbf4c90c939bfd8b9c8ebe45ed61ce2d2c9064ae13883a3587ec066b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c2641f97895a07b2ee5dca375ac315ef9fc8f4a2543bd0a17522a06602e72e385bfa0e727ff30a6052eda73d345aace490c392dbcac998a935d4496cdef7026427c037e407fac7b2529c38fd23521c6c597f087c75782cf38b5db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f67b61a13d8ad7b43079444c6dcf7a0e639cc8027ad2ff94074080f4adcad9e086b7b1de9ae18df069484bea9c2477b7466cd31130b79e3048f2af905f9e31b8d59fd0e18c61a1a5041f9e60969d82a4b53d3e4012969966b9d9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8907170fc54e5a844d2ecc36029e56ba3d1290815ed240404e25871ee4d1ff3c0ca8dca1c340d705b72234b1de36a2a0c843e31abe90f9f4065fe7feca60c8b8fea3094ac205b2dadff18f68d076bb52df0725114d89a1ecc506a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fc1aa3d0c8074e0ace1a40f07fcc73cf24ced1e016c2761ce0b93210eff1d18ab1db4cc32282d3deb3b39138b582b1388446b6b3e67100678c73ab292597cde5f3c0e62913d87da73c74cd6e2b68306f05b852bfc24c71a33712c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114dd209f30ef5f5ea961e0de726400715606f265ac86168b7860a8f513333828e2a5a92f052db405c8b44484960d3d9c3dfe3f80fee948e7beb28bbb815d343b10bd2f84e73fee3b22e43aa84a9811f5d1ffd4ac465293503c1535;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6a4843153e465598810037157f583cc10ba96ee8360feb29f122790bc7dec0ac5b64ec42e91edaa6050e3a8dd3a9b4e0dcdc8b076fd2529e4155aa3c450a7f972b3b2771a91a93c8198f82a88ea5b6cd68064634d919e3e8f90ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b35e63c63b60215bcb006ffaa6c8ab22f8a995c5136fc2388778b962d50f90a565df0bc5f0b63fc8e3c799f918ee179dd31c95ac7c81a80bb93aa3e7d2453e7287ef81b105890dd75f176cb057a276c04ecf2999af13098ca2bc95;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b649899bcdc0fb307cdf8e0530f41d791ec4365e7ec0c0b00899fb552c6276a5367bb40cc7409c9efae5e661935a028dd5c045127ec3b814ae2faf63fd5b652bbc40daba429f0473ea6cf582bdb2ee51cac64a396873569ef343a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17692791d18003b49dad41113df533d4b0d750460984c46609d3455b492654957d0b3f4bc095f4a32aab1f1fe9f535f5ea50e1e707dc670d12b7f41f5f2a764b1d0f02ffb71e1c9b7b5eef0ea9fc0ad2adf6e5d8840423488113469;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1761b4850decedec33e55d9013c81a19db16a79daa01ed7bf0bb913eed263e50a8ec095e1889cec753a6d079a38cc609793c27c6da1449b56dd3885f624f11e8cb1ff3ddab9197756d4bef45d34beb57128d0ad6fd9b150093d938b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bb95bb6c8771d317198c3b2eaa7cbcf74f0a7090b1c68d63009d8d479e9d434904a6c39064332aff2471f6df813d0d00c41813c2f0f86095d7c199edfb9b4aa6796a75ed414c868aa2d10cbd05f1240e720e13572f0c8f8d7afba5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137cdc6b735be3acec1080e6d53a7bd1f02047896fa32d75050335085333013b33c5d97fd780eefdae1e2a4ed76b20730b2dbd08b554db02887c77e3b7f15cf4648195dc6a099122f3112019dc93ab31d63b678dd60d22dab4e0c9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9637e7a986233a05877a14de383a2c8e7af9377edb4b6f43b6778eca15c3e4508a9f5b1b0fecf8058cb6ccab3e07d2e6e6aecdf72aac597a50b626a1ed5e2fcd5507040518942c9e0792fddbc077de3b0f156b90d7a5a3387a3d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d655ed350ec2d44c00aade14eda3b8a78b9a339521af27c8eb378f15468f7e417c5d2d541b8c86d9d052ebdcfee8859d3c5f56cb9006f30e12518546ada4934a2f78fe0e4fa13cd8123636ee7eddde26b21bb3724785e03e590b09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128c1e693db3ab813be9a9f6027a11e373345bdd3ee93572a5bae4f6ed17759e580dbc93ec7ca5b6028e4344e7f41a4452716cd8660b971b5fd20e19fb3e4298b1c1acf95df6025081dbd7b768712e0856655885e5afb97bb86c225;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62e001e75f14a8fd83bb9de7100ee018561af00e25ee3a29fc929e322b6aa1fabc53f2e69c8cee61812c945faf7981d5dac211a817758657394d34a0576074218f9963a0c846ba6f8fe94291a85254c5cc9cec5e24513abb19eeeb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb15fef5f11c29be4257cfb9ba3187cddbe6c7f63594a0e84bf5ef9f353bb7d92a85378473c65103c9272b9fdde004902fce11116e7d303eb00e4f84c778d26f77c0936a354e44ca20cca03b7b1d7dc880736878077a27578459e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee05dad7e4a94ece153091f3dbc1fa398c4d312338978bd39ece70d6ebc08edbc76e8b1fcf9121f9a5b061a1d707960b1ecea8c158e5711af8aa0491e8ad3ef270404982fb4085d0c7adfddf0a99eb096d0004e43e1b22406aca8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bd19a378909cf1509f16d7c3f5746b739b8e6a1658410c1578abab66f042eede917624f52faf4d53a815d54e659a913972c2cafd1f5130fbef71c5d942dd4166aaf4368cc4e77208ae04915c13c1a7d364ec96bb8461892dd93623;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6fe0fcfc946944f1a06ff8f28fea57345055e4758e7774546233b0eaf1e35611ab8d06e0f79e34bde005735ea6a1d44029b63aae8870600444069276098efbc13ff36300a6b9bee7170935f9851c2aa2c6ddf4c163613367b520;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd8743fb00e57a41eaa79f9b4d1ae17a7960da2394f636cf7c390747e41af70a7a49347db1ad22d5c6fcd108125c386776f397d3258662d6468d6850a332d19888a2e1f0d9af1070df07562be896891ecc78e3ac2d8bd714e31b8a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2aeefd3d30384a51497e41597ca05115150a79280dd9ebe3bb83f599d8135aa2f0a625234f7136f9fe3a328794a10d8712a67a9e3df71a11645fa4100d5b992d1e0425e3d7ed773c3617749fc30e5ec4098bb0f6e53a21bd61081d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154f69747b3606048a13b92194a953ce9627c9f5a97b0fbe2eb393fb2ad61d94782be10ca638f0974417935996246f4f680bcf39b01c49e132d028f5a12c7939d48b736eec7562a488dd35978796a9db5957af39a06fa0f13a602e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189024ef996131a62878e5d03633727aec5efb7a6b6677828cc00e47069ffac84aa78f1030f56427e7aae341dc5c97b7f7cc8d9bd3afe3094f84bb9a31f40526a2ca3f6eb9f25da9dbf993e8f21094574ffb34446846d6f6cf5a0be;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb82dfb6999fc94eb8699d02415a4cb999739bd4effaea11472c5ca2991ca407d298435c2ff509382217dfb9a04998a407611e147ab2e3dd137404da97ecd6d8d8a8e8e4635eda1212456fa682eda6cfdc9b1fa0558f173071ecbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h21c2635040ea329d7c3767116a18dcbeb9b25edff1853f568a6b958878ffbc7255816cfaf4964f93ac739937a579dd4d43a27dc0e09fc23b7e955eb9892c3ca873cb2ef2b586a5c0ee67385de48faa8d138995458b8e6d4b3f1a87;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105ff42a211f455a0d814142fe0224fdbc80aaca0633cd37b77784e0fa70f2288264f5c3616e54d704339d44122c6dfa1177bcb6e3e7b5fd89b6a1cfa50f56bdc8edd016fee39f77c9380d971b01f9ad7bc91202bfc5be112e2966e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1597a198d4422019c288de707398d34a4d482e3c0093df2e356c1e3d4316fd2ed5df71771ddd86d45c540c7179df517abe8e9623cc9a47866c6919f14048d596435be1ef99aa34ce969b35015d491fd1b48613b2ec0be75a06f7d33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8238b65878d547fa521e70bdd85fd170621a2f412f82160acd731b0beb966baf15b82c0400ed6f46d3fbc29cad0dfa65166771eb6b342f58774c45eb6b373418b970082b58cb0bd958b9e730690aaba97bc45dcac94c79f0cf92f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b667005878f7dd72624fb1af4bc6eadbf0a4148c98477521e9593a2f6ad3a8e8ff8bd6c296cf2f7a33064c28f90c282056382104de961fd1cf2f4244bb6a831c8aa97f550e9585c0c29644ebcdea5eb730aa352aa8d3f48d92b04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcc4be6bb2f9f5255cd921cdf4090d212dccff54fdb971546cf91e968529c1b95f9bb544d372a8d5484ffc5da3a065cf8501ac8459108ac0798887274f05fdf25c6b3c21a31e3403ea6266f72ce95099534b088e91f17f829e6a12;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59d9357ea1ac012411322cf9e756486023b13b078601a08474d9794332c723e228300767a2d3ccec168a9e2c0e011e25ce86fcdf90dc45e3bf1ac9fa2f264b3f04fb3fd933199f4af6534a2010a6b5b9484ec6cd9a04a30aee6683;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba7c338bfc66bcb7a5542e794f0a00e1a87b8c13102bd25731ed3fcff9eaea284806cb83dae5305da32ffc4619e5f760e20b49992cc6b326f7d468f54d6edf58c1f9fca0278ababbea409d9f9062e39361fe13c1d2c47547cc0d24;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h214de0567368499cfea1e7b3867e31e9a9ab686da219ed73e52b0ba0bc1f4fa2b0dfb1f8a87375f18373fcfa436a3336bbdb6f522914109bb0f12d38d549a5f974fffc866c386d4cca8e127540024fb004a19024f7a8e96b3ca2b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h61710697427e41105e4fb13ab8ffbbbc6f69ab6610deb124bd454cdfc74aeca5ae8925c1722a09ed7e225569995deff5c1cf381b258744d3f8d137c0345d923bc1c14a0c31f4911ece630f652cc80ac9c4f6165e85b6efee01951a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81c79ce7463a17571ba78c145f37ba6aac8241615ed6f382413d693434cc3ae362d7b13d5da6396ed2d97e1d6cdd8c7552bfc23a4d5148a3f6516bb62af7c6593f33c90f4521ee9f6c71e99ce78a679b2771419390e79b749f4ae2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186f05b58ecb6bbf69e9fa61066c2ced49035fcbabf3c9397c102f4b0d116b2e8613d8c31a7761790af9d38cb0dac67cc5cb928bc46fef861f468449781f1f637bb3059843fbccfcabe92d6375decf133c0f8a07629e98ad18dfa11;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7097c290350df1e30a44c95298b71f1cde21044e9fa8c2af13ab0e7221cd4aab0ff357a69705262c08f1d5ffb46b1a865dccdf255fa848cf3a73682ba65af5066c944d5698a1fb4daf937015956a7d7d1aa7000c207c343f92aa33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f13b984e4584639d6da53e6b03a11fcbd6a67b7d10e200d30b19fbbd441daf960e826df7d667c46e3ed379bdfef19ae864c9a421a165ab8b7e88b3bf39ad9a06c10f6471bef37a5967b7f023c1b8dc80da84944ae464059073a75;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec0a20e04901e716d5e0888fe146fa3ebb1f76fb61afe0253537739b570ab008d9bf8f294e23fdde8a4602acb43147e4ca688eb9c10061fd305abdbb2824c6f1ade8d0a2802a23a61dd28f7cef7c23077f3cd548a0b718da6bcd20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d01e76feb15079b271d996438936a3e8510526f0026e837cbf603b5fb63fd30f5b93375ac2c0e47a094860d32a9f64926f385662567a92122dc62af2c85d54a6867cee0ae04e36e5fcfff0036d88f7c8bc42d38407520d9bf6ea8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc73fd8131093c0956583a5383c4da23535e107cee52975cd4f3b40d54f827bb7f6139d1bf777dd883f397b7fb69dd9748677753be1f5ac320355d463968ff72c803e6d7853b2d6dc5eb5e576bd5d240b2db9ab18b45fcb0644cde;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180aff6f491b0eb0d65b50f647814d25c973b536d27b1085cb7c9d2757929d845fd4ddc757ba0ad3cf4caf7415f63fa84d0f2e7ec64a7da5dcedcff455b42510d0284ac6189ab88cdcac6912621409d0bb266a8a31139f81e745a96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188bf8d9cf8195cb546aeb79c057669e8983b5ea0f6b3c6e772c61cf964ee10001f399a8486255ddca6c3539a0f03e701e744469a0355fae0ee25e25ce5328fbc5920e217f2d13a6e550811e8277a4097248af7fd3cb7d3cc7678ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h371648d999a74f26444cc376ef8b641d832e2dfeed284be1ccf9bde41da486445ac7ba70c5a9d0a41341e7cb721f8cbdde17f95501424d8de42e14e0ee5e6359e8455c0dacdb21d9fe6da54cf00b2b09e930073d9e413823a06db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1e1b2b77dce0d7101ab19400aa4bf17fdf7274f0ebf9be8e3faa02ef0b937f96faa0cbb363639d4815af1c5d9e1e6cff6dec029fff064d848f389f95586d1ee909fb8bff70251404e2fd3109a8f641a51fd5b45b5847af0c2ed33;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25444509e9db674ec8c6b85164e7d3dbb7f8e4fa08275d01691be727400c7be280b7c20b9291bd9e9927f4fd880100f27f442d37cd0f8c42c6a94b0296e63202790dbb7740a74352aaba1a432eaa75632d767b150f2bd659d5c49c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1442429432f0a981e215607bd09caaa81ec9bbe912fc5ff68ff5a14146798670945000f864502dc9af1a115aeb0bbd26773b35ee0518dc4dc14d58959ef408f2ffb42f769d8a819f6d152471d653b27a7e62e2f1c5c2b7a249dc6c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50b83fa4c185da646f56799255fca0477209bd5587c4d85b8f7bf5c57e4b7e68057e14e17c96e717c8edbaeddbbc7e12592c8129409013903ba0132f66fdb3f083573453a189d523cc3ebcbf162d4ff0ad34ea2cd3515f9348a155;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30aa1a18cf9c8bb4bda2cbf26ce9dc038d55c847ad9c68fca51e66d7bbb771f646be51698cbed91e26d9eb7f4bce7b57a945af950b66ce775bdb8616f82676bee1329e9321f851431ce5c287277fe0249859afe40a2da7d904f0ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164816c1e9779375d45ded1c86379f8d4bffee808561fd7ca736c7e6ae801489d0c5209df6e90be1430c849646a031e5d2ecbfc94319a919f7dc58de5fffe43ebbfcd02241f465e3a6662fc239f791cbdbcad7d3d8d3f7c27477cf3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc177ac229838c7e8bfa44a150ff530fc8c3651006de8472fd27a4962e695c1f5d75ef0736b83a6700702fdce929c748b6f28198318b7ac51929f698d7eac7f2e99de79c3232cc9b1517fae2208a08a003abf3d1a29b34e335be53;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1996f507dc6874a9463643173493e53948521813f27ff2c686b310162bf19048daa0e5d7c326dbb840e8a65b29001a050ac9b3c200be02e28f546ba61fbf04e7654798fc649a462fa1a626915a402ec55a851fe2167e7f1dbd21415;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17dff613488ade3e33951026e66710996a3ae5d2a9e115988939afad7caef488e0bd382f12493ba6330aff64f09e682a201b3095405f9e612c55e6ec76c118535bfee62402242d974d617a49d81fee7b2bcde86cad6180bf2d4fb0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h943389241008003cfc6e5fe172fd05212199f45ffd06e042c5c6b959ec4dab1774bb19fa5ea7e15141be6958a0d6cdde3c764b479d8151ba0224bd2f03daa46b7f120d76881068f0c65902780e47096742f5b6d431f2166be8f3f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e622a6d7d1ffcd1083a70e9df58727d08dcaf2b7e83d1f7e9cb69d4f4144dee3c546c5ddf727d24878a631a919675496891753c64451eb79c676b1e2ad94c7c5be973b27ee27b9e8af24d205b6939eae639cfa45e930e3fb313ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc354c738f26e9ed18cac4aba7fc8e663e18e75f4553403dcd17e5f161a1381bd2e8a716556d74b276266a61d9ba9ec46f7afb9fce52cec5f68e885307a248d9a7d3421697f8ec5c43eb59d2461f7787627b19d6b17c3a9c703e408;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9b9af8d94f48d2aabb9a4289de1c913f715c1f231e67324477bfd0d10e873a32615a9fce3c44b1a6d5657f9588d94ae595f2ef14996feb871907e6a81b302d165e0c46bcc568d1592c295352eb89871ed81e027be8ffde0653603;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6feb04c19ebb0b39a69ba3fed58dcd7ea0360474d3d6b0e122dd20a504339d52cf6e30ee2a6cc0f0a9b237cf3a0d1af6f75ecdacc0e22969840c2583039259440d4db0b145714d78b4004b63113b34890e68892f0ced9c337b5030;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a30924de85fade43b7241c7b911b949840e05f998b3ead460a0ecf4a6c7ccbd3e28f473ce030d2ad88975a3cd5851dca6313398635c4b84b223dadd973eae49094cd10799d7879858f003b31a196a3ab3d1a7f0465f7472c3aae4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha47419dd8df94a8768a0336e080b53d0b6cd29fd6d0f8839ecce893b40386018d621ba9371ae9e39ae36b036bd00c1e0f7f1c899b67766cb7b473ac2987d42bdaf3fc4a8d16ce1ba30a54af45ab19b59bcd2404c98da35f4f60a67;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100b467a979ac3d8183bff8f5ae43a96b0c8ad535e36789b02e9fc431140d4945c2abcd2c6b5db67d076d38d81d731ec3c9aa382e13ba2f7117796355f5ae04570e1fdee07897d0f21cba0f98df5325c145e558e661630d795792a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h282c0ddb9a3bf4bcb755841307698bf2cbdf5ef031460efb65bbdb15003b0691b874f70a41b95b71e56c0609d3eae874c9ff260de5667cdd24b19ea6b964fd15c9225d50f42e7a87eed9b6d82d120941b99b054c3302a7f1eb8c75;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86e01164ee95a31fa6ba1570befd424048e0762b270781593ebdb5117eec603764111f9fa59e2985e0936394d232290ae7a0a59696acccb16b4494e1c187e0c8113d56f839f2a6b6c20fe760cbaf90f3164f96e1101108fc16f3a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15fce5a5a44c273e73b7afc38f49c7f20f6850ad3ebf566590a38aa1faa9fe43c15cf61392a51fabb6884b53d4bb7a44b65862a2e9003b03df8a200188ff8337879c2d01ce527a977c7c8b6fdf694eaab9f041426461b300a0806a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fd58f204941ce6a885b1b7bd343979c311203cff69585ad4ee36c9ad8f1fb3fbe5e4c0277747dbf0377d2db529f2a2215e66f80aaf3b9a6d4333f9c66dcf425e40b6fe0961ebc4916b23a282b50341becbb89abc06a19d21be836;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f2fd38d870e03d8eabd2c654cd7766d00251967c5a82617168f03a7a25e095d4a22ddf651948fe93fe283123a6a790dc07c8274803fa5f265baaeefc047325a27cea186e212c2ca5f63f3fa6911a2bc8c12f8b69d34a9c368d672;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68fbed5c6e6828f218650dc9f51e72abfb2ceb7a64995aba28c3b14c04d72724fcfaa8a8d2b09a3f1c98970fea9058a539b853b315e2ed5e2d68d53d70ae290c468d02584c7d1cca4d03e785356cd9430c3c8018b760191af68743;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0594c287aab8b8335033938edf0ff89a6a06943ab826c3c5593e6ba4164bad5e70f214e7cd834616528b81673d9f768b96ac9f4280fe5fac33e229ee864f7fb92504c37a992c4e72a8d7863528aad08a4f29bb65b9e4c5bf073eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be2a1eb6c11489f9758f26fb7e6e9dd8bb1188730a5e05229ad86d780686c8cc5aab5acb4f9dbbf1783ae91b6983c67582bc8969e8b709153c9a030d7c0ac587638727e20f86e56dd443c368bdaea6ad3553b4d8ba2b2583bb8775;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6f1be8543095425118e4fca3d4b6acb7b2f0d536173e64f6c3eb0d7a275003848663b2bfdf11b33ae45a73a64dd28522c0bdc5a1239076708696203acc908be1aafcded4e04806a0f8919148c8efe15fd8a29495b60903a946107;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13bcea1a359ef60862995c5a944119b6bdf2dcd0fa06179bced6247dca4b01aab8b0bcfa00e2d286fd6c1613b1615f5007d1a0d3bab41ed6f37abe9468649c426e91e855ad104d2ea53a068d93c0fbfd02b10336835e5a9e25909c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191cb37b53ef00655e527cb7937699567e548fc1f0eb98f26cfe21fa09331120366c258bd2f6401980248d15db348c33097319f0155afd3391a21b2ae1eea277763824eb02f6ad1d7787f9818cea95809ffd6404f2ca32ec15bfd52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e97c684a6eb803bb88a2aeb9949f2cc4847773c5a8eafb0ee27f88eb05b2c86037ea8b65af0721d11de687b83de3c82ba8e26c12f335ac72b974c774f59f5b4b726db6e641a375185062b11f1d8ef7b96435920c5032d56c3201;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1621cad5f73b82ef787b03d1de11c5f870abb0bef4d96e9219662b5886918375d31a602ba98ee0e0b8f1a747a0a9cf4e33534efa09e079111828d2e219876da519c20c6fb4027cff006cec2ea15cd95d940f25292d292fe1d7a566b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164922f2c7f950ab4c4444ed4aacae1cb617154eadaf75112e801e72e1d74f4c621b2d54baa25681195ab1cc29ca3ee7ecef9c6b9112c0262b6352bc324bc79270ac368067706022b91e8de3fc4b1632b918bbfc971dd3698b67b00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h94f651ee3a42acb5b5c4b1a2eccdb9754e5fd15f8e3037d477ba472fc3aef0273c278b728ce8f1f23bc9f5cdd1e91e93f9e23e367d7dcd2820f966d096bf8c994f71ff7db93459a65de3e88be03cc0ac60824da87860e5c530af7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb76a10a08236775eafee6781bc32b48b87ed703ea2fa61852a4a9eaa4b9ffe193834ea9e707965cb859d7ec14a816a2354f6edc88d9c02d50e0e3de885d31daa2ad380b613b6e0800cf2a200e6bf0c6afcd2e1a8480e1757f4e6ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hedcdb89436bff7436d68cb85ca7d12a178a0c7297135dfd0bd1e48230387e16c5f81ca87c269cfcfedaeecbd8f3bc24a7685e32acef0a557348c901723898ee62ab8a1dd72537c9f91ae57522b0536b4b10e97c215efc10d181f20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f569d7f182c13803cc9591a0138228432a7830a4803d836bffc223ac23899f0c9ecc59a6a2284a92011223dc082ca0a59929068ee6c2d4fdb97e01b2bc4bc6d2a10174b3728d29340c24c7f88bbacb8478d51caab10cd9c814770;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8636dc6c478725aeea684cead325efd5fb320a0638e80c48df2d1aaa14914803fd1bd6fa3cdf17d208fed929c5bbb8f95996e22fa7c1c771e2966b7a3edc52bc91fc40e44ab5c9b96970b7dca2290033cc049ca8c4e26cc0b4ad4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1776aec12456fa52ea3839695bc7d6f2dd4d4a166eb3ff08a0946a7089c006bbb7e319c05aa98e4b56fb69511d4871287aecb8ff68b53c67af240b579e5c4fceb09715f22c700846faf6e24ec276a660f754177a5bab90d3f250ccc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16db5e31774018ce31b9f583a42c849ad1a6741fedd61a62618bcf47db6e678f3847f649219852041a5addb1583a0c43e9ec46879436021d5cf9a1f3a5f9ffb71e58ca36ffaf4ad9fb4ba33b19bf12696ac15daac7abe7d206989c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1394e94733650b30250a36bcc72a2d739d0b080468a0de7ab7d642a1b82a3dc13ba98fab8c53706b8140b43b72f6a5a7efe82a1060489b506fdd16517e5e3a2ba256719e00cc4bad1d0c5158dd9e0525f7dbad06f6a0fa6d576dea2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7dd02d96e61d3aac0327bb3fcdc3eb3ad9e966b5750facc6e1e71371f3eacbd9014ff051f5664bcd1c501ea210d799591226f86e8a46d34bd946c402bef7b23db59632bb65eb46ebdb09733d88f12f2b28c076f34cc0e66e0b158;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8ec39f7e1413bb3e0810714d8a5f068f75086cdef17635ae7ef368957e4fa762958aad67ea1c2a990977a921d9e9437ea23871b74af2ba86d50ebebb92566d8aedd8d9b69bdc99ce928c537f7921b4a1fec80a3b0a18104268f1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fd821b2a5e1b2c44cb09cb6ce49897923e0dc27bd40070b733595d38a56cedf404bc651cfc0acdb25bdb2a5a79b50d101fab87128764961d07a5b280b591090081cbc8727eed5719b4e342603814addde4da7a0a8b50218d15fc0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ca78ea08e895a9ebdacc7d93641afe03dc0e26f1d26beed274c78642b4e06d2dea9b35e309123db2576608d331aff836f0fb7bba2e8b808a23a046c48312e7aa6e9712711f84827da1ff3422ceff015650440c733442f35379326;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcfe50fd1681c536bf1881dd647b55fd9e717a5eaac69bffbdc17d12138c2e25d3f4802511fcf7eeaf13deb9974ba325b4e1343ecd68a5b35408c7ac4b4b1f395b4cdaaf08f468c82fdf8e127729f2a3a3b6a2a41add99d624139c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ead94923870da3e706c2c3599745732e35c6bd5b5fb2afd956c94d6853cf2a97507bce95f3d9c90e96a2c4eec072e42bf395488bc951a8e80b2ea306e961578972fa8bb44e36ab9978e2b7580e7fb8f107874bd8ff908b7b897c9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27afa8cf4221adf7579f866860cbcb53307d0932d86181d2c63179610e064a9dcffd3ec806e25073746e0bbfee3999fbb10d9eaa3b40d4dc09edfd4cbbc5e22799e7f7a4c2e483f6eca44e6009683ad6bcd3ac08f3576254cce20f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e4b45badd800ed194f6d67023d19eaf8adbd16dcf9a0d1be5e5d2dfd94ea0b0ba9e9c7e42d18d981333d830beaea8753d8f598296139ed15e8952318a3014169e1c08c2da75475a8211b47630d277292bb25db04ff848f3350a37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe2da87bebccff9b33a4464599210aae129d87bc5e0374479b1f7588b719d7d2ac9324daf7629529a638c172cc1922d00311e2a35565a4ace8ed4d12d7a3ca6b430ac559ec00b7c4399f432f397b90deab63850267134e3ad66e68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf47b497ab2576def74da7824ef7ff3d10d813baa44403d4ce53e71cb7b7d06844150de1129a5eae238d84a5c182ffa0b65ef464f1a22e2de76a47cf1d3517f6413abdb04934aa98bbd1b4b63a7086cf489c3e4d1ec822688a9467;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8177ff6d9bc8bb1ac699913255307a3030cbb52f2a3f7b6384c5413c5bfaae9f44da4deae93851e5f22e964c281429e4622b637ac789e0a812cd92015fb88a40aa89e2516f200034a3bc5ff591ca48691788cb0cead578453499ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d4fc6aff902b7ba52c868a121ee107872d0a8b0d7b774c13291060d88a42c784c02b55cd570ade0c59c85364e8e20e364a0b0192e82b83a345a2fabb236c85bec8a8cf0cd921821ff6616f45cab31d37e03717399e4b25f5471134;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5dbacabfcf1a788f477f08977f949522cb1045f47b88b74d395eb8ef9fd76f63c70e4a5a80b6efb214b9dc1973502de354ed27e21d02a0ba2e68683eaa495bf7c0b46e9baaf8fb1cbdd4a3218ee21dbf53a0597bc20ce7d0c866a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cae0e5d2c0cce315dd5ca2d4cf5a2315418d6b1f8f153c4ce62e6bf20ebe91484c77ce5ce3dd09749578b09082ca3e7782b2ed585e7508b8240af32ba39edca5e015c8d14e39b5bd8488e8239fb569dbe4aa198aace35932e5eee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9783073aac0d2e9b2112559e4f793ef168bf6c4ad037260008fd133acc2045ae717ea30984306df2fcfd7944864e6735388132066d1322fa20b2c81a9fb5d8e23492821ccd58d67cc32168fc2c418d1e6145b23992cb4257df6b07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f18a06e842108152c8693fb6f1863a94b4550f3d681a14a9dc85bdf98fe8b3e6eedbe80e3d7627b4ada1f41d64bc8607018056c48c67e72500556d0566df7874eb69d215fad1a2b3b737214a828c999085245e9f143ccacb4af34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce8935dc429838a9d71c8225490a5e242b0b07597b86c29f8aff0cc141ad90550ed7fdd32e574f688b6469ef2143fc175f67920608bf908281518a22a832fc238599b13d976d26b7bbcff23120e954e720d68588f0bd66dc0ee846;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd21cce9e64933cfb09f749661e82c52c3e85c1ce59e0e0e141da59ed197d23a40febd988d25d2af440ae60235121363db6d0dae7628e94783ea9c62d4978f734c663cff176ad30ee7ccd59ce3b333d69dc3fc977125dda51314b22;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ed5350febfd26131bdc51b1d1665efffbb4206385b5f225c6462097ec3e7199a4b4bb22e395173ea89403e8da758ee2533d95e899529920933ebe0857a7303a6a749ff45b16ccefdf87449cf150d54228a5a5bf3b4e0de0027acae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18890bda6e15d7c33e26356162cf24c105fa71e0749aac4b19da3e94f89133a6ad4471ba7ccb0e8fb45197de8164ec4af4ba7b1bb55ca346b1b9b442aed577ff264a1948ca6d46d0c5a6e76141bfd3b773c1a7f8070ab5a21e46e6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b111c06765ec2311e27bc974536bc1fbf508eef1fade54598e26dab53c23901f893177f067adb2472ba35f302211f116726146c0cd413c78124b5fb3b5af4fc8451ae3b9a56aaeb54020fe2a1e0502aca0dda871ba325ccce7617d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95bce7a53c8de20002e14b7e7fe328f2bbec870004e20b4b0428f2bf852812220b21bd3a650191967882c89bd80d427b7d9487706da5364ec699a6525372c8bcc863e77ced481eab83619b5326576befef67fc18894eb7241ea43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166bd6196f0e4a9d6ac306f8850234c8b8276666ca4b4d13e8c615549f8f774bb8e402299638e9f241ca9de9d071a18c66b2c6f17cbab2ed1ac530141fa88b1e28d2ed7184ac49de1a6d9a6f83bed36dbbfced1cac867d0ae17d3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e77133523e6c157010e2fa444e0daf6bcb6a18499beb14f53e0678a56a27f3f78035dedc78c24429924796498810eb750a912b34b44b48aa977267354b8f456385daa9b5fea961cca364c795bf837ac6c078f0b287b6a7089d0106;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1279cfa71651fcbb6fa2b29313552eb71db054453dce6a82447f0b560df0492392f918b490ec35e1741b84f1c8e2800b8d944a7443befde6d1f3d8e08e40c0939c5e4e2ca57efd945ae5fd5aa8eccba540916eb2c05796147cee69c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d01285444a5c440f5aa909ddacba53b3026d9660d17870a91ea0eb095aaeb0de4646d094206da6d310a80f341547f70259fb57639bcf98a3295699012bfffb452c05910b0ae1fb6140489b5d1d9dd4b4be10867c3cf61c6671b80d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5d81ff0833ec1345a21670f290bbe09734a3b0887b6fb551567cb5efccf926566dced9adf4a77114c0f36b2697f49d2c891d10a31c2dd7cbc7c60e780c59d88850b8fbce204f63ae454b8e55a0f66ea73a29467d1783d9af24c87;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb8cd3728307750936039f8d184e997e3892f534a612f0cf733a54f3223941e1627e6b92f4db3a2c69780232fd74dfa8a2c5bd6a0a431b6976fa1662bec7cdb375e0ceec3ef70409f67022eefdd66e3a5e47770b29cc82e2dadc70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100aa91039e947ea5f223f1a52d8b0821bd945521b8faa166c1aa39658aee470fbb269bc319e1dc67146f23eb04cd11f72ed657b7eadfecd9246e4612e1e15db9089fc1078aa87b8e75dc0d9e4d925becaf1f862073fb36c3f1ad1b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1586cd0295f6527493a6340529b73c1f286a0b91e9b2aaa5b542cff3d468c1ab10426ce507b5cae4eb5415bc413f82f864b63bc08093e72558bcd3f6bec737a4a5ca93e07d5bba6df208101d24df9cd803f44cea37312407b00a467;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c501bb8d779955ce0ab20acc1200d86fbeb231e00289c5601a041ec77d3b3ab3081541fd7b3d51a7f9d0050d07d490d0efcac57b9076cd3c9bd2193508b0ddd2c33836df66e3826bd0e7bccfd1d4335baab18a1b3484a74d1dbc4d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6093d1ca5a31b25213a27bb1d5a0422cc0be5b5bbc8e4ac0fc212c227574ef43f59f0390d2944076d7ce3f5a88b63a430aa15ba635254f7e52032d0fcf197a5c5ca4f13f367c24da65c98454dab52bfae5cf8d8712d5b1922a44c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c25969886f7b3d8f59ced3611b67aa9b22f4adb8f042c59538b8a8566295fcc4e4ee570a5635a720c05acf9149a4c1be45f49496268cc1b18ceb4b4229213a3dc20ee26e4749dea990def27c486f41e6e178a3f96b83e0191c2a3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a71138a179dd0dbeef2679b615acefb2e85ba3d41d5daadf65cb095de0ae77edef705561d331ccf8cdb1b998fd07589496d95122d4248b05c7f3808c7b311698ea5abc00c39602d56455f6c161a321fec8f278a66e0fd7e144f2a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36c1095b68828428fc4e8527d26cea2efd9f26afc2c48f0960f96cf533fd6a4d75adc751329d53d8a906f8705e2b03a1810ccbf2c24a2bfcf478427f1e617bacd45c02f26109697089baf5c79852dcd1fc5892abc23e599102560f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187f7e5455aedeab04b0f3f4c53a0a2b64db655d3caeefb6a5b688b53b02887c3a6c20e4d1837f674f701b8af06d302f44a8f770824d0a7c7e10507becf9a9c7918f075fd988f05d2746706713cf735fb4fd583bf737d6b7d980c07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49002c698b23f06300d1fadd2bc6d16243740fdf1d0c08253b0bc8320dee4506511de6d72eb6b4c835224c039e4c4b4ab62b229a63923a66af40e55d4433e63b71fc9b8d944da5a104c7764b75e47134c874ba9078b3b39eac4587;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80df4de8e94aa61e9d85079ef12836192a46aa881b249f305a420d137b3481c64c57ab2a37660b84af03203cb53d9760cd546bee642d2bbb17b6df74670c91bc1534019715580860795740d08b959020b9cff60a88b9c75814339f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfd09e486234781fd51465b092c0b5c574c6d5841881aae89ae64203cf28a74cd940db8dd85b3fcab6c29090a1c8f9ee01ffbfb1cc11fb7f14e114007b2df63e38f6f33d98bcafa7bb53af996ee8bf0740fb41ec3539202dfee1ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c70d791c371eeb55feb8745d2cf0b6a8e5ffaaaacd869c6efc0c4244828b6f7e004c89b97a7232a7e3bd50c799b604c6c6c9ab9500847ffc1859c66a3e99190847944223d5a28473ba1c3f14095ba2b21c1db6b79826b8540b97d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a8348fd787733ac1321c6060c042c8e61fe4a11ae87d14c3a888b042c17bc4b0ceeb077dba80faa2a7d769f1b64f75a191634afe0c5cb540eba86e76612a6150b162ed0eabad5c9429c55d5feb582db75f50771425f621db9b4ea5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b622d19ce5ea924ef33ce0254f213adaceb24518d8703bbb09b97005c525d54219edbd7e4efdb7d7eba797b4b2badb8095d95a5e35fde07cf35b0d4929160f570bcc2ac25f04fefefa774a13bfe87f7577a3cd7875f1f5ee940a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a69d43f01acc5f18b499af470b4a163a5a898c2b0d41a978cace624b53ee6dbbe3b5cc04298ac81a80ccfec39602bf6c114c775097f3c8bcac230759e6ac78d8fbf4ca8dfb42c10392a377e4695fe752b3a1ab66dec9d2f80e1f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7d6c2a99b8e395a6eac448d192e229d630b5fc15bc809aa5d0ac22747385f09b57810b1d0a2a74a6e8d833dc44472e34462c007f9653fc9ba6b5627b50cc2e6fbc638e6fed3de1aeb802d58e8897a13c8ebe87f3243ca9c369fad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1579463d973907b2658b3ceb6b697911b484cfb4cb9a207c6a0b20f65277eb2c9bb1b87a25555f419c632a943b9f5e2305f76428cf35e055ddedbd5d12a91c18b4650de08cc89aca8ab6711d58b5e2c625d8bffbdb5b077407703fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4db25984a3356ddb31d94e987807d6895adb6259fc9cd2bbfef997957d6ff4ba201d5a509a52f7391e9310b6a0593dc7ddee34e1f38265b4eb71c6edc50c2eed7d7fecada22b2e8e17b05b60acc39131d88317b1f6f3123d0fa587;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec371a27df8ea0ce5471ba76870d20a26f23e97b8cf88c3bd1f40c6f759139b42026cd1f2effb6e6f7a1b6c245b0ab0134fce8472640fe1538e35bc46b2120a4ef2be4be9a4bda51e62beeb71f8d4ae536e303482039f23bba1141;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24129cb47d8ab7e53472b2b5c52e60f8366f9cc10a2da1e7832e5ce49fd04f1293daf93e9e1c2f138940b9f3dc957e7dae318b5ac0fde6d4da541017a4b0b6a7040065b0512c51f875ad7530d7a2c9acf765907a5001c03a9665cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1088de70b6d8e5b16992d2fdb7fe7d1d924c4942a8c5d266ae99882dd92d520ae19a0c03bb5fb434b5a107c35c9f4662f35dbde3baf5c32d99c7ebe83dcdb326bcb519eec8b0f615cba8e993545d851a9dd761db3fb722db7aa0b70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h675870c2ebbcc0aba5392186f8e306a969605c38e2ec917746062e41c08be7860ff3b986eafe06511594d7069332584898dd4b314231e8be68867c690e31dc9abff14ff3d6b2930f3e1c746150ef4400fd5be3066d489cde50caf2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a9529e428de06406659adad40c9fe6d93b766e826d119660febfc7e6aa67498a4f229a58c02de182967f018e565e4c424522a809d7639d2e43e801df467e37d3b552a03dffed5cffadae6854a1db7985d8b75db592d6e18661022;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h288d352dc45c3cbfd3385f93088cc82d29b1291262b938345e431014997b6d0156b86bbf5f3e89e4ebb63f0f2838f3fab1c66c9e7004efd472e8bf428e258c0974a4f8e8ade7b1990e0fdf8cff88fede44352aeaf33d3986118657;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbee1e1d2b50ff72ceccf4928c1356a73c41915a7206906eee9d991a7431041e5925a1973a5f1fad16717b35189698282c5325d8279ca8e4b058d8b54d383c298cb0e18add7f60c075a667b96d32e260772023b8600b3cd7183805;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14588b63cebe45db8f206f7158fcd87e3510548de31832b5f088ead07a516e17bc59a792803bcb739e425eb89241396a97273ef23456c2b112169cb8f4170fa62ebd4022ef2e0ad12f279393cfbf9b2fe0e63c4349061aed7abf2cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7d5d9a2b48befea762489737198a0e56fc1a45d6ef51d212cf696d843b0156ca3d5a248c3f7276def4d0cc5ba83ccb783954ab594dba0dee3bec46ddcd7b97d4cebf4a81b1e1fd54ac4457b0a769f15e30845e5b05a76cb9af8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e98cf0d7681a306e9a126923ac13a83f1b5f4726140ac73fb1991d2b905bac312675d212f5a1aa93ed617b3f30c1bbba0108459e41c2b11736a1eb2fcfa7b73b7c1771823ea97e9948f17a6c407a82d57cd2caafb07db0383607e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffba10fe22104d1cd9d9fda4453fe4b221ce951aadc0787343948ca6c84eaf89b974bc036563322bfc97847089716cf2e62f1471d45c4d6330e536affebd270feb5bf5a911cc87fb2e028b50da1361817beccb39a2c59347f7d01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43654d196f4890ebf62e4600f898b92e5db7ed003688669455ec61b375e3a4c7384481f5537f678f4d902b2e0a2953ecb14ee8d4aecba49ccd001c413fabeffcb51e935858fab382711915e1686eabb156f032f5963bde9aa33fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133bf9fa21ad521cb4281de3ada900e0c7aeb96260a71b4368b5d8032ce97ba2fb18f9d847544303788bf3df9e49d3545a2d271ee3d7a844aa8e4e5c3787494235f585975ba15d3caea222d5d0155dfb02fe5179f782654c1ef71a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e5585fe372170abea5007b6ddffe9728804bcd788fa60b5a377bb0cce1582057c64527277d17c16ec680b058313520b4089031c70dd67ba6337ba7f84d766f126302e31e4a3cd821a48f08b57b08520bab5207eaa93da15233b76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d4b3a94f38e262ac8eb31113709c1b706ea2eb83247b7b136417eac2858d29082c848a2b875ea360656188520b09d6052093d5a09519030aa2b9f8d0803abde9c6c45e3e020a345ff957b3c53854d2fb36838b719c69c917b76c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec90953c74b41ac4da6d6df945a31eef876767fae3deacbae284aca1349cf00ecee99a1e263b0508125f17fbde068022a16e99fbdbf826bad7083be8f4823e6ab13c64972545bfe80aef1f6bef98345fb1556814675f3389b71cce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h258a5863ea5519e790ed79c16a2ca7fc67c7fdc94b5809473f5ed7cf117e155ccd3c206133f37182dd338f526ba09e88e2a43196e2850c3e9fe46917d3a65abd6221f9e8e3621a3781e51d5617396cde55d6f7dc01ac876e14797e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148356d535fa67f93cc9aff66af3beea8397c2b524d7f1ce2714b50fcaa71f1dfe985f22edaa461b69cc80715cb97fa2f0257c88abbe651ac3b327ca4a8518bf8c57caa8bee78058d5666be94face24daf019d76ec67ad0f6703903;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168b10c52994dfb005b4200afe26d80b7fb2e0d8e5f9239c26148191e7a5e54ff0fe4080fc069ac043e712837c5a1a5544d705610d95f9a5b87c79cdf182cccdd64b210e3de2fdf8c88b9a355693f86ec4ac98ca6fab758035c7421;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1479c1a286fc161a5128efdefcd112b5d48e2c4d3215805e63c460b2b32225ca5d5ea24bf641d3ae318c0d20e996137c361e0637dab267e5cda61f26987b52db45883e4e061929e2e8c6d92529d02e387614389cddef98950246410;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8d7ebf47b4bb77e6340f691f7e7c327e011f5ccf06651eb566ea62de01fcedb7a831d5d88e646bfe4b6945a93a83171319737cd64bc023a328bacb0d48dd0cfcf8cdd10e77f7acd5e69d69b4c694b4ef035af5ce89bc6949b3fb8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181a71311daf3d45f62dc4649a9844c9c44ea6635e4f861e999b9a729751a25ecd1873d1e292c85f29ce676be1827f26d9cf097a3ede355f4afa042dc50368a2948a1e75e968b276e5d0bc41a691d3644a839b71a68a33b04cf0b07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64c6ef525642cb92349033041b18e1c363214f8bbe73f2a3bd0d046f64b14cbb5550615a57ad0197b16761867ff119a33668ddc36517e0b7d8de4e420868b41a8b8ce28a4a47fbee1d816ded53e7ab0583c0dc68cc9be0b105f91b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ef46322459563335055db111a79a544c131a4fbf1a7405dd55cb9ca09a14e512f9f38ba55e618018fbdb2d605261256d62a875830f258074e584f8179037b39927b3cdc03919a62939f882c458975d94bc2259658493b784da5a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183417a53b0b8a2b6c88f9c494d5a787be2cdc37c11415c941385224edb17337680822da7e45e8e96cbd83d50c3377a09d171fae62ad9c51affcf7a37fb70dcd62b97caa70f40117c2f2d3a61cc98094292cbeebace7336c631ba04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1198ce92882b63395780f4678f44c715d06ab3ad84d395e540b4c9f7f1ee23eb625b3b5f6a4bacd36498d684316165f802f242f1508f322316c5825db30f055b101148bb03206c718503d9f78f48b796ec9b4fed5b962b97e58fc32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dbdc591f8a441dba8d778adc385690f86cd56be2b6f94d20519ae2e842ef27a39ffe94602e88bd964d80abcf24d09a5d4e1b4ab43ec44cec1ad4e3ff3ed4f8a551543113e6efde5066ff0ef6a9c84784ca11027071d917b9746bd2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a83cbf650c7d50f467037162ea73a1c651f4ab0946486ba5fa7927052cd106e2618234149972a050e1dc37b1c3b1b117758450aedc3ad1ef98e0af30f70ed2333c22d6cc724cae4176633b56b32aae34205ffc5f52dbe396c30ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde4694e7e4e1391bf2a4c8807f956bf5a79cf8d4b312e6de0d597991ef8b3df626aa246da115e0e0c9aea6fe7a108d5df2bdcbfaa860e59ec92939f4377b879c6f5e9d367edcf65de0555e050a8042f34e3b649b2069d33ddc06b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d94d8299cd4b0966c5c389662cad04ad10aae7549b9ea4dd19bbbe48c27f9ec67aff9816408b5551836072c1e1f28fb5f90646d91c0b3807ce978957419fb7ff1a73dd8f560ca612b90fbf0e12c16f11fff6394898db7b9112201;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9515dfaa71a577db2edb362ec297651705c7433ac25b99875f1c71357be0d4cc76d1624f94e114f428418deca84bbc0e37c9e2325f9ac650bec912c2dcc348073ca3dc99c7d74c07a15f59c54effa820d5ac422ba3545eb96fc1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2f12532dd6d304ed6d1abe81da4625a92217f79e80567f93cc323f83578827a9b932f03dd57def236d497787564566bc7012488d14af2edc0d46c2fb9cb075ec3c4f9ee214b7b19cc2fed320ca94e02b5be1319d15394433d1556;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19800122e713eb9bcf8cd193e7103203632229347d99a8ef48f0f7b3fc55a312979442fe4542e7a02acc4b51d5655920cd55792574b00203d6cd3fbd734d6479c7b32af4a8af526fd171e3cab35d8d9692fb6baed0e44ab09e3734f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97b063b510374d17232673650bd2896e573a152544354081e6f32242c3b2c6228b9692fcdf8279115e7a33db323199ced7caa341996f220c273ef10547095f73cbb2fceb8d18af68244fb9e0bf50798ad233b863a0b0c16b404257;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cec9e2f0c39d34722f2e3c6227817ac630c6e5711e995cdcf7b323fc71e1b5eabfd3b70a3f54c9e8ed8ee9b55110799520cd321e9ccc6d978c3ab1f955678286d81c969e7b12075cdbbbbe1c20c98f41dfbe80191e74418a4ffc7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1874a159ad0fb0a41934b3a9fc71d9082d7c85bf124ff06bc14a394c9afdf70c272c2f8fa64e1ddedb75065a96642056d45eef28c12893f451e204d49d7b7be05849a9139326a560b6ea379257e4e373ce9605e7496af05aeb482cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h593e2f62d1411fd13f4450ca93bd3e979e47301f24f7467ea0988c4b262afdd20054a280146be0e9abe752e8b7bf52e89d527c2049b31fba9c086c82a718c78440628e94609958b89c4e4e9dc83c09083e5303a0467ed397d6c48f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6c2a9119e25a257d40f27505123db409708a879fc1d1a0be8580e415ad82c93165a1312ffc8ca7d4e492a3b0941e39c8ba1323b037053ee090e02fffa06be54efb83c22171dfa977678c68bb081f856182c72c568e8030a8e83c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb35519130d7fbf697b49d77cd09788cba54501a5be3539ff766f08e6725d0a1b6d3cf3765fff6ecdbc4c459c87ddfbc6c72a2b3c218116471f5407be11d057ac45b776fd7626c529de387c0374d73b293f498440478eecdc52f81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4efb10f6834af5d740228c2b59b275ac1ee7779cc8729ff76118041a67181767b13934c8509225203d253fa6e5b210693b1ac9cf8d34195c19e833bb468a6dde2123c8fca0f3ac11e2facfae87f5cdc7f4f9f33bc15cf0d2924fa3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he796123ed8d50d09efbeee202a51342e6e286feee2c2621baa25b37927d527d301c5f594116003a7b9a71bf7eda7eb7a99d8cc7873c1682316b8aa488fee50f8a636086a555bf617844389bffb55405634e9b46e500484a4888ccb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h223d24daea880606b9fd1dca633e5cbb6afb84de63b8f3b35292623688a8cd6dc30a6fa502ddd8a30455664d810bdbdd08abd59a81fe868261cfaeb288207fe68151cc363f40363236a015151136d53f199888b5680fd3e4d32727;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha94dd33c6a505587c9ea6da2913f7d9d21299f23a41c37a08876ea781023c0c3613074842f9bcefa51a46cc217b924dedf3c25f002a4416f2875f4af36d1a647ab885360b423339adaf18d6ccc6eca6ac2a93b50c0bc27f2ee9abd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d16d6c4c053418b3297dd1a74cda18e954fa7fe4e33cfd572ceee39108986460a38661b36116733f87a82c29ef4c430db94ad8fe7d4e13393fde353b348beae7834a1e96ffd39e0d5e009478833f613f464be723b8c0278c12391;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36661149731d22536781dc9176abf0095516bb3dbcaefeb2db11865884b1a6bc937d73cc4e7620c7f616909820cf4c00b80e4eb851646df9d50bf8d06666c4148599363950bd4481f8959b87f1db9b88b3c6d41aa95cf2b80d5cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c6a7eae6b25805f1783c9fdbf35a16fd50471e0c8b0c393c5719086e50cbae2c220087e38bdfefe959648444a1f46d7e6b6a3068b7b353958b46c5c9f37f31e1fcf144805ccccbdb34ae62411a16cddb1a1afd75e6a62f86a2c4ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1604415d1834c6b51fdadc6e5fadad94b6ad7898fc9ed8b1b143e4c7082f5fd775bb99e1b02f8793e1b4fd0e9757a215f2313d32beb0b4a7192fe489c206de9d69f59a776e60d81c02527c88687c4f99eb2ac4a7c113cd14b7566c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c4e6b51439d19fa340b6045272fdea826462adcae2f47a654e990e8da46ef317a896694d29006a3812a55da62bf7261a6842a19f41812338fbf3efe4efcacedff8b86a829655c5c50e3eed30eecb0bdec56ed5adc8df1f239c553;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164f6b687c173d104b6f9f01331043635fa9df0f7592a406f248338ed73948a223ca117109da739a454767d6996632b07e924dead3ca50782577d12c1b70c4f90e17726d89cc48689be8ce25eb0da63b8d52fdbd24f267fcd0bd6f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba5904203af3bc5a46bbf5659e7dfb4445c562304c7e2bd7263827b2d7f39296d0357f17ea653aa54f8dcc57e058db26e2cda5b7c526ccaefb5c2c5c4e60860c5bffc06d2470876d9ca5578d2f1ab008e5521f7a1d6c0fc590d4f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c447527cb2d95a267bed453a96b2fd629f367df01ee3c51ccd4ded90823a0caf5eba6d049335d7333b536eb1d035198fae4820af49b269f06678638ef120f3359e67c88f03fea20bf8dbdd135b0fef5d10ce5d17834365d883cad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b53a4345f71537046e52f3ea2d7eaa204a6fdf6683fb3f6ebfca721baefaf8cabf837729f123f4735fa797dfb3f45bf342d109e7b581c9b29c4f6d0cf79c5c40b374049a847562f076c18e97be241b2b8fe976d9c5da9026f536f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha039ca992419b57c010c76e20d227feb489ef89cc233f87096da3c91ae27cdae4b2effd552cacd91476f7b4718a5e5930401264faab3c6840edc6dc3643ad2e393a4364729136cd503c5d3de44066a851865a5d206c31b6fe21618;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd27f5dcabafd58e14358ab36d88e0351fa57a3a477e98f027de0ed51b60ce3af39c7976af7baf231d0f635ca15eda3b7320b590256c49f782cc9c51f21227f447ca48ae4776646930ccf9d339c3590680c96be6b5c18460668709;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1316e805be4107d34b7ba711a7e678299993d480f553fdfc8a4df5ecc414db62b2acc60c3a9b8eeaaa0e2bb3d04c2f97aa5d8f73526f3fc727f8afdd0c854ad4b34adb4ce51e3aba8c1791d0933c2e60285d4a806bf35e40ccba5d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ff6b396b8af6e2b6ad32be38dfc70b9959d2e4519190c702f798cb6b9db1404b310d4a9af8c9ca1f29fe816dedf016a15e8e743c3d71543cedad3a8843b2b066b71f80889eda31ce06e51d6cc821e0bef034a54862c9cd4bd176b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb763c91a6320f9dfcd42b9759f276514de4cd56bac9222640fdbffe6db0e6e4996804a13413e13322aa8b2b677413286cb47667294915c2daf4e6b4db25b2444e511ded170d0a289ed308182ffab61b2b109035ea0af680569c17e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1244e4fd78299c617182483ce0cdd3d31b28f6638db3c4c44734d71d848e27aca48378b03ce43f3e6f4abb1a54e34839dcf3b073096c3c0ace588cccb24e4dec850f455def81e16eaefddceb55e18a46027a1dad656154e72a17073;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7ae2e886f3af0b777f4858acd5756ec31ee5ede67615a625884a20d8ed6a2592d3b9daaf815d5741223cb114eee74053c858e6d4c9d115c1e52fd5633c1319706209742b3657872851b2415e0260f9c24fc81e9ea4f5772aebe65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1340f4306064375c63e936855af6701d6a03c7147917f7165f93323812ee2527c9c35ed364ee9d8a25c51701f16185cbe31c908a1ef70fb27fa51a1f058243e99f3347fa61927216ed4ab9909be639460c8ddbed9aa1ba657eff940;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a65c291078795bdf3b83db9d76ecba468d98735a2d0729d904a0ec813a9181c3bfe435818b7f86dfd76a2b3400140e30c95647dd2d600d8817fc4a0e9127eb8fbdf20fa34f1e77320c7e61910187be92496829bd5dae7ef7587665;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1900e9d166f8c7bb18e964a8e2464dfc5b33edd009baef50f85f7be5dbe302bbe295074c9a8ef83f7d3c59563908b71da777f693374f891016ce3ab0d4b802062005c2a7a5236da1a9feedae5f5f969fb5f9a42032d24a86d1d3ac6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1717987f165a3ec169f193196a04041f92cb7bfe06f9a25cf8cc134e390ac77c8ccb383e1ad9539040cba4ca18115f794615712eefcb7e7a59d829a8d69f59ab1fde0be6a57001f9b708804b93366a9e9f976f3190914f63f2c954c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9fd298b60f7324a0ba710894125195e235017b7b98a3f4878e9b26cf78de719486620b82a7c6c3b0a8da6e7416892f138c6e6e040a979a3733c14e57a1c3eb828605113b6922637fc70947731ae0fcc087f62f3288e315acc4cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h82ce09336326ec2bad1fca36ce4298a845581494ca1ebb1edb0dae13f946bc50c2ddf71eea11ae25d0c4f0cce8013d8053ad4a8dd490a6fda25056449d2e50e4e9ce051450a067db3532968bb5fd88e41d108cc6749b6a4160e79b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152937ed3df9ad9dc668333aa3bfd27f23510ce2dc170e78fc25c56fd0cdc5b27af85f173882ed91590f6b2beed12755ed8362dcbd152d2b94390c966f81be48c2028394dc9d4af82debcd180ccf69fe0c2128268530ca600c8aea4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6d25f7538bf84e9772f06e8e02a41ca25da4b6f96b0225d1d4288374e8f0da26f45ffa7698a2a9f0ccd9ce6b544af91a2af77e87f37371e5821e816b6a863375445f05150b178fa3bbb71baf93ace8118d201f7eab22310d5b0cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd440a325c700447ce7b3ebd709f8111eaf573652a8af48da2dcb1834a2179f52c9d49f0994b779a0847c42e7b3c31ad3279e9ef352a7d2cf1a49e59a7c0d5ad1f7c7c1fd5307714487d2744aab998825a7c3804d5bbb9c6961bbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197224a7307cede46ffbad71044683c03d32c20911a889221fb1561f52c9f30255bb0b0b3b9472d137b0f8edf03ccaec3f6b065f49592fe34fb8fc6028f74b31c89702e5dfebc383bd21d4e05f269cd11ae628f38611175ce284e8a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha59c93425e4bc1855454907c530bed235e2998ea796c255c04c6b6702d7e4552fc6fffe55f3993f0d688d87e51710002aa10466a5e37d58a44336ae416718438bd7d2a806c52b9ed601b229df1afefac629093328a8ed21c907aed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8fd33b91f9b902f29d09a4d552b5fe589da30dacd322520156f2ca69b32629b9c2b0750d19726d339c202dd546b54e67f0d61d8c6831ecb093f83feb7e8b020f068bccb670674438ac37e251b675d6fc619120a80fa411082a7ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4849091fa3d2eee9ec8f86f77eaaa2a55c6b91d6f2a74b0618e5e6ec7744213ec969f13cf92e9a08cf554be31fcbca77229754f107ac9f33d30ee56da8d34826d179fb87c09eb0eb1692a01847cf8a1b7fea32d36229fee5247d94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hedf7e28537236434a6f634752a399a93f54a312e1dff88e9c68e2466e8bf91d42e5be4d56d99a436c93ed8ccc677a936eb8a9727ad030016d86f713eb6c38a51723cdb09599910784b9ee2f50720186d0862bbd5648816146afdb1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20624527d3317416d24a16e2e2289998945db4bc363bf170067c02bae852576e2387697bad74a899a632b99bb5615986d9bc95ddd7254410b412a9733e93c95c5955a0109f322fa3e5b9440f6832e3a740450ab4b08668688ea4ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h303cd519c78047aefe5da4c0038802190b766cca1a05341cb68af2da113567d325561dc46be6447800511786659f80b3c73a4afef1c74564337f2ac09d6472349bbd8a48c0d35b74ab9a7fb0b86a106946959b1db96fee6fea5d76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ad3d68a8d01667779e5f2b0dd4169fdb4418e802d9e26c92852232f7c7337eb96ed2e00c1856cbe7e95dce1124a241cb0482720fdb51487cb7c5271e10f383d46eb69f8f31824caccd0e69745588ea70a51bdb808322c513af1de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7cbfe08ecce3b95fc435e099e19da7add07f7b40051e269df052a8830d5b102e258255ad05f4d1bd9218b453b902d3ebfd18c8c58e1556c10302918bca4914aa7eb538d064b8cff4cddcf1223df594cb6089614f770c8e9c87bd2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1d1ebf0a585027a574ce0cf5b7f6c78edadaacddcad38a53280efa545c1bb72a57b5a9ec21084e6bd6ffb8ba7eca055986ab88596a70f457c5510bb62bd5d0907a8fba6a6d08bb439adbe29bcb3c538d2027e89973bebddd3e93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13ab39575550b33d7faa78e354d599badbe3e8fb4bd70c59613b1cb4c76fa7b472761aa9af63108d705bfff29a5fe200b81953e9518094782a0154c5c00e2156ce890540dcf5f47ea8b355bf5c1a1d60adc6264e8f8fe8edc46a98a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc0034bad1c04b1819a919d122e9e7e169bc4f8d579f19e850897226d328608db373a2952af9e8c5512a004753a96873a2af69084365627b249a5ee0268edc1a16d304134f4d399eba5677dcc0719926892b0d92caae90708ec207;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf8ab9533ba69067285cf434eba0f7c3a1de2f9b6f934ca329c2b68023add28ed48b662532c158dff187f1a170b67b429235495162b205dfbdb7df7a9736be54d87f12236ff12969c48abf2c13cfb4c6be5cc0d6549a5c66271ccf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fab71c7f54c195885c324b5b9e9128ae47af20c007df134371bd35f3a15d5890de5031e34568c9b56f4712373d50c691f4d1360538cd497a4d60ded83f8813c65e8cda1cf1070181f2b6563ca232ca54075a4f925d25b1a070020;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f399de1a1ee4332cb77815ba8f57e4607ca4e73540eb7fff3f75465929c1e2c39aead6c2291c8ad1b16df39495e1356cc4f252862b5305fd3c63afdf834563e8b2465a28571cf065a6eceda5ccad4407c71590f3733246b7ead07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6db50a98cd1d90f35258ca5e6f1ee7ed87af9c28f2517809d8ce92a017d533b8c0b1fa8106737ec1bfb2c9049433d5f4a7f60a3f5a7858fd50dc1ede5503ad1e40102f0182bc9b8e1f28e483a774f85c0925cc04a2eee317383b4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cb233fa27e46593c832b08beb2635a293cf6b8fc6bb3eb4b1b0b5b1916877fda15221f00099d74a7b883a71467441ccab6b3494a930ec8953fa251ba15f0544d15800d09372aed8ce7db79fa9f44a04939b7ac0ba71000e77207a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf7f856b3e0aa19d2c24e694d6af169e16453666e776bd1aad83289d2e1462ad1ebd5bdfcb9e2c544f74c996565de80db9142793e1940da3bfea01875f466da4c7c2d10fd8b460b0f2b279fd50e970aa28a015e428db575ae28665;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e21819f81e4284930f6bbede3878317e155fc8dab0b7aaa6b67544e235140ebc4cef64dc4f177dd9d6c29a7abe1d1500f3d64e5cc343ca841747d179ef8afe81b100c737ba4c28de6ea3016bb73f5993bd24626da0d22d14963d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c35790faa9e843fb0ae6c7df78af0baf53d1eb98472640ba4e204e99b6448d8a4cf6aed93e85fab13dca6d14e34a889de57bc0cf8eded8100fcda1203c512e50ad6bde1739d4e46a9cd263b6ff4f7fdd6fd7460424823a0c0a86e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9f83de6c42058cc70542eda1cbecca267ee6d6746faa26d726d4bc3dead8466ede974e2db83ee000afeebc2aab4dec733dd2d4850ad9ac8b85bdf62daecf5b7c8520edcce891a4c6a3d923b38e2315a2102c3812f235f41eb226b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaa52dd8209e1edb4da730c7afef3b0debbd52f3e0286b1a9cb0e00ed6e0d105415fa976e2f50d3311e20d657aba2dcc9526c63f5fde3ba12c21e3e921ebab3fbd6022f741c46b40e6bec3e637ef9498ac9046cfee25f449926b29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f9d8a07ff9b6b42df1e63807261937994819fc8cd5ddbbc1f019a2bca9301729e4cf8fdef320fd7da8c64b800408474ab008f6ec1b4acb1a283cf2d8ab7fbb31cf40cd5f2dfe5527eb29bd9b019d50cffd53c40eb64e4905f7db7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192618a146a40a3efc3cf8924e4587d33c8b4f17d1d13cfab1927bbbf8bf81c142ed3c0e7bdeb261e8014785a86279cd9b2913e0ef9ca1020b65b5eddeab463738dc519c00be94f4bbe5c9b96d4980613c424a6b0ed1ac81391f064;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd0613de6ccf3e473303b2b92b48b5021eee51d0df8caba6127f10a87a0e23f19d133b2920676624c213ae66a52d8d342324431312f9d862dbcdf63927faee2d0b83794296566ae391302ec0a6366ca1c9ef4b6b1b55fbca6813fc7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a01c78cb973546e7e6c7254200e41edbd17e3b01f5b89d2a1e471a177c582b57648e815223e149be621ec73c3bad51226181b0ea38398d910a1e0c79c02f79283cb171e521f56e9d5bae3ea34b0a1f28a86b7964f7dd6d5401500;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaac2e865b656d6c31902a5508a3dca051eba40f9b6281381963760b6e217a2bca5e334c34eaebc5c42cbf7ff8bb67e2a605a7ab407da90c4d268afa3f42e4a90de0d788a996a45a31015c67c651fc29ea78d119bb874adbb8ae81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16dfff1dffb9185f9a741837c15261f09f18351a0dc49a2aa59e4953a2ca532fb5d5e4fc5284f6cd560b858994ea14e8ba9a5079cef8ae60cc923216679e7f1359ba0d8a5c619104a89112d4a397e32adf22e95e2c084bc9fdcceb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1318bdb754167d2a5fe5209c545d80bcbbc4ac92191d0e616f1de9fd01fa5af6851bbcf93189893660e9fc6e05cf07ff76022be0127b47225075da5cdb8502cd454d3bc5b67de66aac6a42d0140a4ca1cba30dc7a33c6853715cb8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he93ef3c379123414343fd72911afa17ed90859ccf4f903d874b4ef3fac79c341dc243898e2d6e7d08d8c408a92b47e5e0100c27f224ff924da309dc38111c61f7133c9861c4c1642d5362bc9d952debbf6d4cad7ee6759bcffdff1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a697fa151f1c0a22714844314bfafafc45f9eb76a132138122d8d895f492eb9158815c0a2abbcd1e3d0a839aa0621a2bb5feb53c8fcdb0218ef4434b1f1182d61dc9d58c4bb1d041fbf9d3f0ab6799d2ca085b19dd7666d756a9ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h885289b06a7990cec1733c835d4b37e606186914fcf480ebdae0c5c2622935f9b0b1f534d0bdbe074134d74795175e984267785bf455d360123860b6c4b155d7ea2fbc4ec8324b7ca9394c05c322f510751bc5fde7fe7874dde52f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133d031b4586af08f769caad3311fc94c608d5e7d57f16527a2ab05efa9e877988bd57a76fa0fd45c9742d3c95331d0687de62f3d061a3034c0b58dd90de1107e7324dc383585f519667ac23b97c68c13ebb0138f9c77d0b878324c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191fe08e3cb20e1d815ea7a5c0d14b3c758b956507ee153f5d6220163c4235ee8e2d096033e37bb1d3f9682cc844703725fffd604e79a44c43d9e41023439199e8ff42446fc4b99214a2e7dc437358cb64798313bb8ccdccc96474d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9308f50e2bee2ccab5a3c3745debe88498b195696a355b657c53720804486e6204b4084f6fe21e4fc4bfc2e87579f8389e1c552c6a8b4dfe0ba33bcd59930ee4871f302ecfac2c529c929157b8f810d6208c9518f09915d439d164;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6356ed28af0fd10c2ab36e9029cbed407b58c97030fb1dbb5c1a05c08c307a4c1e05dcbd9f91994911c582169dc413d1924cd9db639315387f69290dd6b568c9b83879adde7dd8287a17e5d68890eca41e03410ab7d1a76ee04fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113ea09cde5cbac01398f8647581e4a9afc15641c548c37b07dbf819b04a0442847d272075164c04ff662942c4fcfa530e8843fc40ce590d6edf750c28e77813ed1cdc8ac7749b8dc2e1b9f9732b44877ea4fc3858773383e7b2036;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79b36eb867b6e8b2b6049bd9be42145b87851a4ced75bbc565ab2e18e319ee85dd8b0911d2e3e7985d379dd34150d39d439f58ddafcc663311cb4cc3090b7584664f7f9aad2614713772ac2bbce2a0bb1e230243b50665b613b9dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2198e8ce218051d89c083d560e2dc1a99f6bbb22ad56c746322252b3d8e86bac97db1d16019590d575d545707bc16173b3e10dec98f05a65567b0cc9a443365a21843dc1a09354fabb453c240cfcb76db55fec6aab4c8b9f4b731;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2cdcf72c12b6132d5eb81384f90a44252dc84700762cacd3f0ce775d75bc62a213e81dacf32db791b248a952697a718aa0bb26e723d84c8cd7939b370bc901e65017cf0f0bab97d90cffffbc0380ace76a81d7a72d51aa33e56f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2b54c1c329ae1c929e0c88f927df5548397287d07b45e491aa99b6c3ca1b763aad9dba59b57d9576f63f0186bd3dc6e0dde5d23cd738250967e25720766940c687f7ad9bc5e923845a3dd7314d5f1e23bbfa92f050e8c66f910a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174b9ab4ad61cc49c0f66dcfd66dec6587802914f3fa88c4fecf16b7431fe17cd66d1251deb23a1a208c672b6f95bd4c222d11eb0617cc39bca30fb14cd7af797bc6694d1936b75b4973fcbe8c9ddf0a7b8032726de692097b733a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1130ffef02be0f741e492d1b09a9b1175dcbb29ec62fd95601ee76058656c5bfd47ce5e825185bad76f4853334487db813beb43dd621f0f0ef0b88598be93e89e877d82a3811105a81c539f9b18f804219bb9d3a8cd3724ec0a458;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7a1ad6b8eeb6c5baa415342a69444b2915343621c533dc7b602f6dc703ff04b366e34cd2fec2189df96dca1a9bfd24aa847dc146675f5dd9d482979a6aa0d3f371358caa4a5d7c39ab7d73279d8e9738280cc7dc1ab0c961d6938;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113ae47ffac56e26ac7ddb85d64b14544f59dffbbabd955929965d3354cc25bb2ba97f46e35ce58eb41a4f8e8b67c17eefe3c89b372f1b0ba8025e5b307a3359e4841bf316e044efc6491f335c1abbe58853e5199b3281f15599611;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63a51720c185f3afd396fbc7668b0e75d42684322d487258bb0e75fd4d8bd8731f8013d9d9cb913754e9c6e294d9a53c3b7e4a9b0487460b5ee49c3c399b6322f165aee448fa191ebb78562e1f31837a812e75b1bcd92f3883fe97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f65ee47b155f915be8e11075612f055f1a26b9cbfede3827582ba5b847b5d9eb6dd4efb655160e6600a8e3f03fdf542305480d6518eb8da4f57451ad37f9eb46ad6b5de3916bde19fa00dfb5846a710047ca34c76d41dc89c651c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c88a3ea68d4bd18c8f5436cb4ab3a14a733c0dc29e0790d1c9416c13d0a60dd446c349443f4886c21464ad2d65c4947759311e36276d5ae0bcb91e8d20066a8fde3b64d310eaec5bb94bf370bf12760f524f9e52965aa3d3cbbd0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32610cb094a525500837c67f9c1a83b9d9d447c2a68331923219d99bc8129f6f884ccda40876b1459aeb45d8b97ecb0b1e5c2f50f45a22f3aa7fe46c1419739e05531274016c8f808794ca9727697ff0f1c4a062424cd29baf2bdf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h293f713ef69bc07c8fd78c87fce039a506063b17853b8d3b98631881002340c2efeff9e8e782e602e5d0cd3077a87536c396d6b162780109da5ad60e00bb1bacf1524ed39bc2600a0e65ea8797a3ff70a3063cb85f0a050b66805;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b86fb8e0b44d0d68fc3e7b65949613c8709fc6527e1c8b59f3f34751a6a2283e0eb460d519759db58e7ba03c0e25559b130d0f2c9c736b19538a9b5dbbe72ce9ee6015679047141a8e5ce5aefb7760749b5c0eb51f60824db3de8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1460ba173303a386b847f6b4c66577e369cabd532376cb213060a8ecce940228f0ee07589862f9f75a7dc15666788fab5fb5222bb0335378aed5ab55ff348fa2fed181c6839f4436c2395e73208885c1b441416451148a1ff98fffb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14277c27b8dbbb03bce18f81f7d776e7c894fd4026bad22a0ef5418952e754ebe5db805b325f090a13155bb86b33b5e0b451a52bc141cdd187069a932085fb7fbc4c5effc6fd2b9aa73c602ace3cbf45008d6f82d09cf7b272618ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5242919c2cf79fb5783f95dece7171c0953e57f004d58867afd6b997cbbb863d138b962cebe85fe1449ce60ff5ba1ea4e8569a4164b6c1d9f69b25a60b407d35a08664488aeff876f5cb7df0165fcb3339d4e81f6a36574f44b6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha213a5f7a32f3107257cfa4fcda9bc80adcf7102f5496fffd5d33a20062c9018b4f035bce50bd5a69f32db543e9f3ddce5b34d33109c7454ca4fe6c7c4d2ff157c16440ffee64ba04cd3ccb4441e8b3582bef3963ebc2be474abc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf35fbd43fb7fbe1e3c1db7b197667e0cc9ea2837507a940fa802c7eb033f1aeedf17afc0cc8539e2b9d6b3ac95cc81deb088750052e8337ff93c776b0d1a14e6ac050b1028fe9949b775e5899f3195129c5071a7aeb6fbe6b3ea03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e64ba4af3f00e148590a9f6f4ae9cd0ae0f24a10e27e459bf4b3819f3b5ed2a02bc9888f27acd2f85bff140792b4a8ebeb81063aa1b1e4963447d3ef595dcd58bfea0e7e27504f0d20de76ed38cf89e5cc0ecd4f02b9be6abca41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd6b67be24f7a7325869bb6c59c1040b3a3c1327ac8ee86898a6702d0caff996b7b606b593a7645c1ff521820847b318026f1c8b7b71726b979a7c49d2d4751a1727932dc20f872b8e35155f4bbc49ef83e66b5e40ae366fe0f507;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c88f9506fe68415765266ae51303a8386a14843a05e3179b1ca720487155de0aa576eca07096f1a092e351bcaa065fd64010f0b335ef01574bef0ff2687a9c40e33066f5a05bf9f97e0dfe280158f38408108fe69332bf74b9be49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b2913c2bc087327a27f0d52f3d389471dbcc5bfadd8aec6baf077df03e7f00f14ef11e779460c80e824c945bddf0a062e79403da0ed4306e5a8cff9956174fc632de2bc1a652a9177412ca22dfc32e67d5364d9876d17e0b620f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1eb513ea61e1e15f8486e89d7fe7acaa8b5a2eb7b408fabfd84fd3c88e3c7891859bb350abcf35da7f0280b9d6b99c3f7e65f2fe52e5110a1e7404d5176a01bd04f859096d441bdd1caea9470641d7a03e86add8a90b02b5ed6206e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1476f63704dad78e922bc9312a3a9971d1ceae1a30eca1b98e8b2e791793b19e0039cb46054eac36c3bbb2514ae6e8acbbdb4fcd1ffd584fd7438e5013ccd1a025b63ff777cefe6d859421a415b190a76707d905a32b05b8f57bbbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f58136d136069b3b077ff3a0c1efe9227581c5ce7885608cee2704dd43ba0f5c294d7c064734bd97d68110bba04f7606fe394994ca8d990607845c1bcf644b7721dc894617cc7b60158e63d0ed101132255ea6b082819dc365aed5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ac956f5c87fda042204054a362af9e518af4c2471de764b693115d2bc50e0fb1e7e1947e4101767f58e0f4a5750f1435f1baabdf9180aa3aa5a4fe1c2e74d22f4cd93baa7e94c3ee7429482a532995ab56d6c5d71350ee95909c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc613a6f3ed70a5251d0873af1b39d4c1a5c511fb01adbf9051a84767ede3dffecffa5a31f7cb1568e6e5a0ebcdb9a339576e92d5b06ae69dc14e185240996a80b654816b0381458c7259a1fab191a1f0bce42c7cec2aef258c6903;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd074c2d3f788ee68a5ad2e34c3232c588f26344b0bb3bc29343d331c492c1020447f976bb0d4ba3136d98d014feb752cbe3e4c5c343a78b69d5be14c6daee3786cf28c114f178b81f992c79eb30ffa2c2ce715785015452b71db5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7af7af0b2994e7a92caa6d795b94988f9c620b59fa707f803046b3f6603f121dad6f39887ce26ff32d47a0663d9fc432a84ee50b3427eee52cbfc4ac2acc1bb0e663247a9a3f6586192e363be91f7e7528de5f8ce7d871343c7609;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c7c81536a7d2143e4e66db00bbf4de330e1036cafe37ea9a79e0da44f76e6aa293a7ce079e294ee9c01510378fa3af0fb03e617362a42a5ddc55ea72e7bc544a4ec1971b99ed85b66f7a7f8315459ff2cb6af0cfaea51295ab04b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f829c41fef47db116597f2f665dd95c746d307c5fd762a546b2489660d656b6836dbbef86a2652aff05a4b32709233b532c958e2854ed5b5032cd576e2e904f8af931155c9fe090c5da3453af50ea6040d9afaecf43ff7f688665;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h37b99a3fd307ccd3c53af5d42cefb3709d349248822d88c975a68c03c6bcdc89150b283e6e600b9cc2d6dae7756d6854fcb289c3e7bd42155f665efeb118fc7d8aa7de769192a2754a96bb99a8285d231b3e027ecc3701f69ee03d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc3bb740561ea217a331dbd950aba5ea5516311e122f925c9fcbedbbf7d60f1d36dac0c538879aec82bf170218e11593f0de1b74700342339d9749081dc90b61894ec66420773190748735195326228221f24c2b08f03dd99824a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5072c57dfe81d85e49e0b6428e2a6058dc4cb3b3804be40ef13cae6d11b203bf9efbab3713bcad329a9bf7cd7f33c3a59859f8f1487bc17d6faf761bddd0761aa59d26c95291c4ee1c99a6c905e8d845870cd12beac638c904a02;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17807598cf5ef079b3542f4737112426ea823dbf22ded1cd758b3cc735da4d25a5dc93da8ce45b3465072b72b9f77d57c8d4fcd6615212695936ea859b882c291333398b67032ed3ad9b19fd3bc225e3f7fd0aed846da25047e5926;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12119cd1f6a9437d45bf7df7a0e4b596b8a4dc8fd8d05ff6e41b568a9c9cf0e5ecd987f198cec333ef1dd0a79dbfd30d86abde2b85d324b38a9cc7b145f118df832472fa3296faed30f8cb7c8469629d4de67c612e1f97c44b7b0eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47d10aeab09dc517b82d0c76d18beef81c25de5223f61592ad79fca3de7d2446b48ec20cbab29fdb58e393c950fc2a1a548053c45362b40b841d2ca1326819b2172844f1c322c67de2ec9da3ea2ebe403e77f50f2b4c0e9ea2fe7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a4e8ec6cc5ae7a40924d6c4d13ab1c29b35ac771417a911e5963e808b37ea8b366b2018bc8c39f2de3f488510a33d3ac49ba987f73314a28a003823eaa134cb6f3de332f2fb918db8a24013ca137309ac4da9b1b5aa56df0b99dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5aabcd2f3d6ea25f88fc61eb18de2baccefb83d65e1e2dcb5849a1197eab13469b256ed450ff175885c99dc524503b4d8a549d359d04bf9cd2f6f61bd08799be59430d9bdffc863f289a2f6e9f10493ec39a0f9a7a4e945708af1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a28f16ea1b4ddbac6064efe30c1f6736339c16e2d4dbb2d225112e04c1bab8145f4c75c283ef42741d0a2b1e6ff6ad89a4d5062dce5bbdbb0e624e8206a7e390657280f3cca7e8e52170b23dce8a94d3aac99a709dccafdfbf9be6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b1978e7c00806e0dc81078078b2c7aecb13a4048583f0ff2a89e6be63c96f2a3c6fc8cf4b74ffa4aa01b592884774d946d51e8ad1710b3c8f71105c40bddb76955631f5606ae35b9a13ae094967d24c9a806331c3433c0a5f214c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4cc2e92d0a3d722246faa3eb8325eee19e46c97343429fee9536d08e758a6611d1ed6036e37f926b9e13fa97736dc653b52c5654cfcbbb655a0db8fe491457c72ffb4963bedea08faca377bdeed6eeafbc221ff8993616ffe0a95a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac4d6736c4fa1fe02c4bc8726b63ed57b6bd8b0a99fdc8332767fe1c721a9a14252f9efdcd3c0f24df205a03d9ca5579ef9f707590361ce7eb5c526ed2b73ef426d7960995aa95cac05385176ed2dd867f7bb55df5dab32f4e2240;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43c05aa1aea1a49d7d9de5880b31f7723de164ba56b7898ac0e4b94a8d3fc859abb26c2c3428e6ce28e58c931ee604ca5d6353d1b4da48245d28b709466bcb19322a325299f357c638b6a18cf9088069b2366d661fe15fadaa8fe9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1e45ae15e7928a09835c6a14746c9382121bdd82521ac5205d609cb003e06f1ec8b40ad3e53a47d2b181743a8f2895df5f3689c21531222a8430ca60221ff1769bcb51f4fe7aa60d78c7c2cf400ed47e38cca3e4ad419ac56093a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he848799e16e04deb6fe19b8e150073bba4700944e5e95818e4cb4f0ff4044393dd20af35931b369e06796413c9bdd5848da6bcd44511590202b5a266e36c2cfae8b14ca5c1e173c13b3a9bb39ff27f94a2e245a4032afa3de37352;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d3eb911518d9ebf5b2e4c6da23feb0dd6160fdd1ca1612d6b12ba51b493c1a61e28ed94d6f04dc40b50675b2e08be9bca824f524a2817a78a7e9a8f80607686bb4af7954e67d1d8d5d01bc52e06c496d9ab8a6bd2ebfb5922e546;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a62865d47d9fa46cdc8bcee84b2e104d5b07673e4b75a7f3160781c638338772926bde4b391ce64d43344423bbc3ba47f22403b12ce0f9d562d34f4d2dc58da0269b9bcc0d788ae3c9f16a0a23db480f05ccfaa41c6327ebb7422;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f523597c3d5c28e8ade063d8af3b89cefdd5d037eab1c2881a6609a7d31dced9c56cb8ddacaec61f84285e8d5937193a7ec68d4c867b4825ba43215092bbe9d547d92965d434f9e04eed9452bccdfe3377b7ca4ebddd66cea6ed2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5056c972ad00c0e33484ed0ab3bd3925f112770677932c68f85bd7e26747fb7736dd80994ec70a003569d84c54f6cb4e5ee49a0b7262c59da5ce0910e4f34c087d8ea71caf219340c03f1bf9ae690f6bb7280957bc0d2cee4b4310;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8008d1166da9f5e1e64ef09c65074038cad960de5a66a49c7d39e279f60f5c0fa41641a4563392119d1d29d39b0c3c48abc416dc242f0b70560febf1fade5b9a016a07ae64b410a87c62b49ef7c94f2597e01cb20eaa2e517bfee5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169c5ae1931953b8d610c728255d9a36280d04deb663b652a7978088e7d379d2bfa5310640647c2207b7e3f3f7e905c73a4927c21365c8c8706222badd5afc00096ac8ab02b1add34f318283ec66efb5adc9915479853c7ed3c2028;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31de87f749c639a09d57cc36aa93c48c2ee2e8aeea7c63200ea2fd80088d92c2f81c8b95e0034099248e91ce1cfe421b3f3c5ce07dbc8e361761af65a671321ce2d24ec8db46fcd788c3d425b4396e0082b4ee99cfd04ce9367b28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcb5c815d47e25393ec51569d7c6bfec85868a6cc892847c49b36c0bf4f2cc0625ccf0959d5750a66ef312d790f077390cf94169347832b7356ac0dd66d469e0d990bcb8afa36497ced51737443af693e73f3b27657820be3db4dc0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e9e4978a7d7b9a5273a56cafe97ddccd1ac24f643c553b64417e713ebe7775f083ae3281fb5257d6a75fbab1ff54c59f8c8f1f5bc203b45342a89a52e43f3980932cae4e9604f74e9ddb4dfac4c274b5f37d3590cb8755430f97b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113e1672594be3d3e190e0081251f3228733d0123169b56a5eb5a2b8b034aeec17e3540ab6c4115cef057a6c434647e1eda9dc3e3184efccb9dd9006cd3db4df6c77615678e84afddd2219b1543d6b492f6ddc54c87b03ed67d48d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc767b9032aca0f07cd1d3a26bd4fdcc56c36eeb63295bf3b30af7bca657f7e15a2fdeada34a85b5770da0105887b3521d7f868341df35dc81d7f189b12fa1c0dffca61dce2dd0efff28011cd17088cb19ab7e8659c69c6843ea0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1426de4636e2fad79b4bbf98007a99176abeac277fe41e03f2376f003afd1e46406e019b5b816204db0e378a23fee10ff4484bc770b99d5308fd2a50a043bcd531ab276e24653a61e99a0f9d8331780ad454a3152e5d4f80e2cd96a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4285091844beefa01d37cf10e5545c7e26cd02bb48fb77c95c662f73b26822a3a9f58e7d48df45bdcbb48b66f0435ab4128b9f77f075f87204eaf369e2541bb282e2bb18daac248efc41e526fd63e23259a6b6b5889c63aebc889f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a124f68305b043be659dba919efef5673986cfd99f8744d99f32ae56a30e8ad76e4964df7c21ba3f30e5678a8ee2e1cae1a0160319b79554d6676931e0aac1a76e15f2500ef803160ce82fdb2c7bb6b58eaae4e240f92a1d24abb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efac8f328a8ce5e67fccb9d773583ded9543b3f64ccfbc2dbafbf5886ab2cbf191b7dda9a29fa5c4682e059c4ded6f9dcaae4f07aa0a7ed1d890945b46bd8c00d6a8cb0ecc9550241b7f8dd7384c5dcdd8e061aa020cc8a9754517;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd34e343badad69d412b6aa0c0012c19677f2ec2502717a87fe80b3b50c9fe98f428ceb6b2f8286a3a421aa35d968dc00bb0f908c1fff0c6d1aad9fccb7c2974390176ac8808754c5625bfee29ea9abf192e82214a4ceb962fc7ab0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8d66b3c41a08429e950ba07c0e1b9f25a1567ef67f64265c79fb1fe310c9029cb7c9831d51b58e1bf96f0fd023be3fb67076a0bed3ab4b095aa02a1845acca775172ce95ebf422b8a47253b1484a32735481aa1f4602076da8cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79470480e2bafd61cfa4f448a8d56cdfb4b9dd1ed79ecffeee5cbb9d2b877f20e7b92b009ab7f6635ae2d48427479ce3bd3f968a8a8b01a9421e6596fc841a4c5d0f38a828f74ea186709e552b15955d5229ae9c3e44eb5ececb15;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e7cf277592f89e3985b221aabc31b43d4fd79fee7565be7cda7a9d7f104b6c6d73a76c9eaad253574cbd8f47e8350f636ef38793a19e945d08b382bcba1e728e7c52d97c099eeb3cda71acc0509dd59aa8074f66009fd0a8800f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189e3e3f3681437cb50ae15d6aac6da44b048f4450ed3dcda40b21d61d3e1384713da17a31054d97575f088111b2354d3f08e8586817335db19a579c99a7d7f2f82d9ec19bcbf45fd856b0be30c881e891b360cda0cc04c011bda8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18894aee5d08638bae56b1e299fa1c102014fb712ad34d58c52b83c7415f67fd5296fb9ea0d531d4518b62a9a281ebb4508047b2a07e0a0764f67fa11a2e40f7fd7849fa7e8b96cd6def71f9b7cb125b9b1f8f07b6145d150788abe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d64f7c68966a023592db3bb345fd47f33b5b60de4cea67710b5ab0efcc4732c98b16ae2596ef20daeba65dd6d7f8dcaedf0e13e0b11cba12dc8aa94507cff50b0e542a53984acbb50ade89d453ed4fa2a0a5c781bb63715cefe45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefca910f3d5c589987eb3d547a3c5e5d95a1808230d78a81e5f67cf6c891f0feb82dc40dc55a57114ed7de510a65b639285f224a4c2bba34919259a3cdfd40c30c3e55f819e99cafc96426e2afbfeb0fc2a6b43b30d7be7526d937;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d151c0b2a023b9f1ff788f3ff058dc31e3a6be6a7731b9b9f3091c063eb1875a1165ec5a53991ce14c458f4b232005c0eb537c80af875b769b8e8dbea926a6562260aaf584c3541f70221c795f78746e86d4c259a663e1661ec1d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80e11fe72f38373467fdc1f797e71ace70c3dd7a7babf61dbdabedeedc5c31ba5eef9aac5495ce0a27777cd05423b56cc648c9a53ed1a2b4dea9aa65b80386158858be9807c4ea076600a09a9e5cc4d1ac34617031a9c30d9ef76d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf321c414cf12e6383e43e27d4c01890fb39fd8ba8dc41d6f39eee67412753f35542ef34f3d53cc6ad9a9b525add39e50bcb7b9d1ac73c4b0b672bb6dce9c76331a0a17c0c56db57289ede14b87cd345336a7d2a254b625b6423b6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa4faffee793c53c64364080c557b9aeb32f4400660faa3a235a9f0c6a7aa4fd60ab4f7e4138a653154e36d131003976451b93f76f330935849c94626fc29f32f812bcde2e16782432cf21eac99903eb4ad2e943d0d58605d6c43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a4c891a05e4ef1ded3745594d75b2fe37bcf828847539dc3011a21c67e1dc243f4bde88787e59d48ddd919ac6f4356b70a565d9971f7eb11ce795f80dbba2f68b53639b9a6c10cf38f61404b7cffbb5143312af3a882708843ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11dcb1eca8e3a5a99237ecae48ad4a87e408509f14c25fa58bd504c4601c7d9e8407764d9904bc3801b3ac350ce7c427681bafddd8608e2d7a6a7c9627b80b53ea996ad997078bade8fea3ddf857ceb907b14f12aacfc69554bc5d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3a686339402cdcf96473fb14221ccbac89003f65b4dda7b1300a1ac00f99f1c314bdf6588b66561ca276cd80a4ddbc86abbee9d1bdb3eedf949eb5537d20c49b87eaab1080fdde9c25eb6a1400c0b479e3393bc8cd6d9d7450627;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h259fc2d6dbcfbb807c19a62a181b113a87fe830c08a5962ae222c4cb252c2069f3de96ab2565101be07a910e88a01d3c9ddedb17099a6bab789764f65bba6c71dbe2e73955dd946b9a2d2eb5be5888da5fca70c2efdbeda0afd3ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ccaaca3249ae69acdd7981f58e995f334500b4ba9edce8f979710c5573eb24bc52d6e2f2172b8c3dfed6010d17c2848e7af125d384a5de1d934bab93856010f11d47af1c30988a87e0cdf43ab9862611cb8bbff2a50cb8774b9ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121da441f164d5d6147775285bf5f6a77ff5f9c9598c84d76049bb058ede73be9dbd02a5931f6dcf63de57260b3fa116aa0c49fb7e257e6b09687a8704d9e54b013d881212454dd80f988be45c29eb55ea0923ca96bf496d078414e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5648108e01ae0b87e555bb390e9e616e20a680ee11e7cca6bbd407c5c4cbc5dd0b4960475a3ab0bc9585865a405f5826a6915c8a3fad57fd8bc0e5789c4fcf9cf8b34b193d067311e873124b00b3d0cff2c666f21525ae02bdfa9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfceb069f0c164ac89c242d97f9e78f7e0891db08bb0af5b6bbeda7df39a3c071885beeb5f4defb6d7cc377fa97e64aaacefe8f0281407730f1586aedd3fce79cda22c947aa62847ca18f75ca43ee374668283e1a40daa6c134a977;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6a24c9ee5d14d1d32884a773dd1647a2d33be3eefdc5a042a22e6f5411a919bb6f4408fe4f1e695bbc8b64ca1d120303d73d0ff096cb0f02399c51bdf3ef23befadfdb43761df5c917eadb5a281085150b589da6447073ad497ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106aaf18f0cb134573d60f849f3e7a1f2871e9d7027024164259aaa73202aea2b4104a5042b04e3098621230a976c95de1c0c3bec9a9e1fca149f621741ca32fc1a1a5cbed220ef0e334d30d8cd84116eef2d96e284329168d2a8ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89ccaf98c2ff4571cc79e5cedcfc2e6fa17b9a9f8a416fdc6a9a34b0b5d14508ffc8b6b738d126c8be1a78cc753454a2f7cb96a9ea290f341bb86535b6fde8b2d35bff4af97820287b648348659a363297b3a4523d02f345ab5d7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84b5d2569cc10263d1d0c2907dda0d806b2cec8bd9108c3d9652e57d4deacb6c3909ae695d7b90d8c123c563d600a237af68a93427e5317073939bf009a25e924d33ac4123d964f72c8cc1133e7734a5a75cb34a781e84be4c0656;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a94074e81ecc940d33383feb709c997d89b515eac03c472d350b8aadc0660d12c87ce6c127dc70c208755b8a3687d90c1ec90af6e2b0ba86a900fa4276b4b67287db228c4e33d1e435c993605cdede995c8f304903652dab5cfbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62cf0447db24c8051f5a0ac45bc5659cdfdcfce49a698d63edcb3f98b14d668a12d790040451bbf8b5da97512bf25b818b611af35197ac0f6ef9ffcb11bcfc16dd42c3ae0eec75640c087b80a3c0a7e5c435a0b988d522d95701f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d9ad15b04c084f59f5d26361f2871cf06378d94befd982cfbe3b1cd63a918f3380c28426008e456827f9854ab43a4d56c63e2ecef6e3149e83763435f95136e7bf7c0f2a66aff1fcd1ea324d69a8a88f198e52c8a489a652b67b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc628904fb28d21f54667016717105084e2da7bdcb18a7755ad309bccd04ecf92cbf7c5170daa23872a688a764532fd74d5b7ce4502437ec966782682c1095d2c54b382b96ba771f20f7c8f982c20c54ce0528a77f62ad175c91c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113f25f17e8fa0a08eb872ee1fcc70cfd9b1ba479b7a03b8f3a87435a9842390ba5496404249e635d3c0092edcdae674bdd1ff868bd081fba4b448bf0e4540c14bf504d02e7fff5a0b60f5dfd30f03a830e9f3486f7d49dab3d8b97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16de8219c020b4107e30d3e4288776007ff7d35fdc6b9aae0b5af4dda8de481e2074c0c7fe4d3b7d2d6e5f1a07348ee0660d1af49921f90984b683dc4fc65807da94457a2e0222260ec7d36fe8c518ae21559431ca17001df32e480;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b11ff981298dd6b621ed6fa575c700fb932b5551841355752fe8089a6a6184a4f159046a31db9243dc86d2ede013c1296ddff2ef826a760da6bc978dcd8269f67ed2ff5642fa3c968fe900e70dd11a936da14439a411feeaea99a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16469253a750a27165de73d1f062b680ad431e3501c6b3c916da69d5e612d26994681613a976a21e1167332cc6f3b6cb98e9515c79c99a11edaac2181ecb5ca85109ebed19542d4770df6bc9cbaea2d15fa8c2fc8ca28e8a0471283;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164ca9304aef793c6b2fb44a73619d40ce3d2583c9b2430d8335fc13079703d2f53b21e89f451c43eb1c8d7ed4f6a23c4bb0c9776d2ee8b04122f8ba7729dea7677739e46d608f15565866ce0bc26b8abf28b11ad5ce857db7ffc57;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he92d1cd296ca277be63c24940c2ae5febaefd8e6c5240fa6e3498f930cc2914d488e07434a05207ea3bac36e70734109392148e6620c29a08405b177a7147852c4ce13ee072a9adcbe13396b8366dec3819161da944563fba42c26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1188b375ea73741cb4d1b677e46c8977ffce7b6d7efa789e5f665a9f00b2b29062e3e753f93840c4c69b8b7df717e7341009b4e996728edbe142d1b5a999d56561900efbb4e7bc90d0455b01dd9b7ae76b18ef7b0dd03b00132b802;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8ce86ec6d7958d40140fa5bc5522876a89eb6ad5c09d23a72da27c4b48dcdb92df5732e2f5cffe8bcbe06a0ab3c0272b08af2007f6ba79a3fd17c0f061137563cc5c90c3f1ae7795fa72bfc7179df494e0b296ee8359bd0867609;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe3d85869f30b289b830f321317ab494c858a5098b5216a559eff36a1c7a4daf2a95a928a38a2d3d30df96bc747c56d3eb5c25d2b66bcd4c037a41b333c125224f89bb9e22952019cffecbadc0f1e4c26b2e55fe076205cd32e020;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1700b0f8cb39166b2700a03f2e4d20cc14dd8691fed8d5195b9ad8ffc6fa430bc0cee42a25386fb6b0e9c76e4293c10549bd0eed179e70d0b79b27aeaa10f872fcc9a2f12192355f0bc438d16107256eb39e26781fc8dcc7ed762c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9e6f3076732c1b491b751a1aef4b74910948562441d58f685f1506fc9ea7f7ee4a2eb868c94b43b648651dd383baa9291058194c6c5fa9f51e80543cb098b2afabb2077e530d81150ed084253ac7bb94e432953ceaf088b8761ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc733f672ffc25d32e7da8d78a05b699d4437d388c255adc8cbc3cfe6a995d00d6c7c85ce6f20d752c24b3f62dffbbbb8d06c4f62d0826279c9849ed22f27568a5bad06256294e0d8ea37f3fb06772d6f6145f0fdf144ad72c2dde;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146103728ac49026fba263bc2ad3db1b5c0a3dee7c8ab1da3d97a17168f35f062fb37d55b8532c2ceeb3709df12b762f9e5a7c52c7a1c015090089f507c00b475387a887f425ce456f9a4572f870f58c93a75d5f7e01f7964184358;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135bad3c0d39f1bd83200f45c19ce9ef3295108e2681458a9cb983fc025cf033b0cff5bdb9225abb4dd63879442ef985c62ed9a82824438bdce20510fa8403db4e7bbfbf7843d5f1a1dc6a94bc3db83b58432a65065b76e0ce09712;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22474482d2e3bd2c19d559a83e87ad4509e90fce6b075ec0a6c0e322131991c39d9665f620fb64f61a0901ae1e5f0f3d3d91a05f54f52af10ffe53d6c252f6d55542ecd00cad527cfffdd4116cd80516c1ed17649e4b658a0ac413;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h797267995ecf8beaa0f994e65ca9e1e4c82c3f48fe3eca5c1aed8373a13feb30c87f301ef3e01178d56d809fe470eefe4ccaac6a41f0b946f3f0f15c7b8821bac493631a239167e4f615a13ca94377441c4c5c1e8763579279ee2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae52f2014532bb84f6a0b434aedd44b6d5af55bf4d61226f956a07e442d0a9703a083ff0c36902a90064484015c7ae272a9a49e2d6d4dde60cde32f86ed1a1f89ff1cbe7a02ad360a8ef40638e9c269f700502579ffb53892f0aa6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97e350f5e7e0016142cbd0b2fa7ffe39030fe9e5c927b41fd9e15ca2ce7965f8d0dc602dd031a55699adf02eef7a8dadbcccde7f479ab9d1e93c334ee8f60f0e574ceb4c5eb7e5392e62b663b6b7ccd917ff4ca7523e42812268de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8f4b3106c5f4f9d6d3584a6ccb7a7b25523135692555d59ea091656dc40281eb91007e6080fcdef4c00b5f66efafb416ced471e83fe661a1dc34735e1ebd3ac8f839bd9377614c15a01c6b9c835eac82c655446bb585dd17bcfb8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1fc0d81105c2c52c434402c181cb0df93f8681d7a59fffd65a90ddc88b15f709f462c27cfd43d0dc376934be1f2c83557323e37795c469b172855e7e869d7b798d4491639926d221c30cfd64846b9e6168815915d1977afdb9634;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec6aac85069a069e5ca4ff2a2f6f72470bd31966db4b36cde8425d94fc3fa38dfdff2d76081969fa0f41411cb2a25010bfe16813e1644804c350dc9bff79cacd384617bf30972b8de5d0efe97609015dc63f64c0d7e6d049c098d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11200efdaae19a09fb1ce85261becba1966588b30ebb5cc4b3a51cfc858bc22ac5d60efe1a9e98eccc6f227e49f1c741c5cb33301f82138ada9cf7ad47d92f4fcceca47208eace54f0ae40421e9e2e9b3b7ad1b34654fe3a5287701;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13204f7fab4802cb8347debdd4599e193070d586fa93cb75c189dca10e854b3fb0ed8d54623c99ba98bab9e47849ddcfa8d964f852be90015dc3b67b3a12e2d9740ba7137cff5ae91a470e23cc3f442d2d3b990faa3bde772fabf9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14becf64242a76bfebeec351999e292e6899e3aedd9c1bf3ca4e6a367eae544ec901ad24be9187b124b729d721070b420f61a142ecd66210bf4bfa552b4c3b55dfe9db9a66b568a8b4e8dcb3ba4d1bc63097be7e374d790e20f5e07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcda5340a0d64cd1353ea36516cefd7878c8ed9a2921c14c5dc102a270f9b4dc1e21e07ef8f31becb218901bc64945bb0379e51a2897c32eedad4bb225430e3e2511454f4cb455f6bb55e70f863af5d1fe52791f9b3925c0cf8b429;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heff18879e7968c65904317950ed8f74b12d1b0460c7f14860d621f8a34e572efeb8ce4ba30e48770444dcf4c8b998d8fb854c3627cc8a9d08e2149d352bc01ba4c251a7251e62a192a652d649afab2c626823b225334d811c76eb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h570dc661b9519fd490f361f88099afecdc6aaef4bfc751a47d5e75779c0eaaca6166fbc3f95418f61b9db42d907112e7f571d3e2275c5a7331b5cbd9d1ed6cf398d68301e7499ebc4f00268a7090e24e39221d7e8063a76b0ad107;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8bde4ccaf9803cf5decbc4432c7b1042ce790d45ae898cae142dfc440c5c720f73d6cc2f9f0fbed11041368e62058e31a251fe13ce8168b69d23e99d844b4ff6aafc17abfe48162af3ee5edba546235d1514630fcd797313408eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f21486231c355c4f86ffd81cc68eb204a14365ae17752badf7775dda6a9fa75227105bf6e75756e0b73b4267219bb47f7b076ad7a4a35c57bc860074ac741ba468245f1416bf5e899161fa7b2ca4ee0085a61f03519e953236e917;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6e53f0eddb16666752b22e1c253d86dd98f4e083cc5bdc64b45de7c8118c401f6f9896fd1577d611a818fd860ef8e0e87906fe7432dfb7369be2b720007b99a69f1c68c8135b2041e6fbc68fdf5f2346d0237377f4646967691bd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12355872c7ade54335d192b6bb571ee9d570d281e2b9a60cada8951d9b03c11c5e1626542fcf4e2487fbc7c56fa18930216b0aaf3acf4011469906dc659a44da14bfd63b8a85072b40a460bd2d1fcffc8e5022ab402609e70d2f956;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190f2ea113380bc5ef8a6838d7851abfaf653365220c3ddb03dba1f90bcd423d0dd174890ce88e315297ffaa8478befc2ba464f7b6f0ac125be7136c4bec87e86e4b06775432540a54688aa015c4c86044a83837d8d04e246c9f9ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d32f7ac67fa723d51425b71831e3a8b15af5f0524eb3e75d8e107e6d76c29c9be1870e69f1565e8b1db3127e3f34c9c1f82b83e7ab7fa7638409eb3bfce928ddc37b0d6a2f960659b97ab8bd2903b851f3a353ffd286a80e9f134e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe26572b546f5d1accb75654db182497036c3dec5d2a633cb4f025325e86133fd839ef4f0a24bcb63f69c474d7380b220f7964e146ab1c4d8b968e59a412fa190eba73aa2b185c6e6efd39ce5f5bfc2f557c556e1807a295ba9927;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13809cd17095ceeabc129412bff1a8a3b6e0b378f97587baa1eb5eca69840bfad5c862a4cd43e3146da68dfc6d634bcf246ce69ad3c9cbcc832e4c958fba604bfe165d7838c98bd978667c22a5cb68b271b892af4b54c5a3d2e91ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f6ba625f75169260e6b5ad8f6fa44f01b5b164741e0984e706c45e88f853cfbff89d96c3943f3d5d37763a8d4173c4afb903f1e4927e15b052af8e97905b7dcdd04fb592abdfd31425f4e5204619f2c7a2517969196ea3f437da11;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf2c828d8a559dd4e88fed2c8466f25548e0e934a151b857e96a0d2dca3227f79f294ca3fb0794f1eafb01393d0efbc361794f17eba0af32a8e018cbe43c075da16dec1fbb4f9275e6fce8314f780c58919ccd76d1755b6b0df370;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126a98f1e14c286955919549b114387d3848db1ec262300c083ff132cbc364ef598612cfec10696e6c789f02b354242a9272111d08649443925038dd6fc19e1d1fc77c968815fcd230e3dac9585c2cca6d212bcc838ff8b565f33ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c664d7c2b276c0914cae6165e3663856ee556adbba2841ef6a184a809d3ba7f87148435f58d908dc19dbbc88afc59cc35f9a50d7b546509e559a2a1656be34cf29d143c40e2f1a61877bd62f3185afc4855bde94b57652a4652f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1fce8e962c0851008a1faf981aa55ec0806573fe9a0c628c7008f00650ec77e469c23fd56543f2ac95d42bc37af23919b20d3d952687b319a4499ff1ccc9fbb787f6b1ba2e0ca7e46e7f8ab4346fcc61e9d5e95f67eecbb5d2284;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87cbcae343308981e12b5d8292187d3370214a5f3eaecb01d5a3903c4fc49982165526c541c3fd6d7ae13702b55b1960521c2adf1fd4a3a90984d487fe7173ff577acfd7ea6ce64b8070d7e00a180a61a3a85920f21cf4bddd8f20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1289c2fb3e562dc14b5c90f9aeeae335f4a3b0926d6d044d993ae293fdf6ded98b6310f6c7cbaa7f856cfa8a8a4b12c8e5b4eaf0a3b505389d26cc757b02d958ab3fe08b21d3a28e35f6afd928768b4f606fce6367330e5032dcd5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15205b02db4a0f69c1576f1dec22ef3e64ae1333d76d470b2dc7e4f08e60360e36cd646ffe47b13fa6fde4eb5aea15d797a7b9aa76794c3f4ad4e1e49ae1b37932174224145bace53bca55a12640da282e35def242e19b48c1eaf9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8cce306440939a29c5d4f1f4af0ad0875610efc4cef86d36932397f0c0a244833273bbe363c802821437a0d471901ef5612c41c181a96fc85d50566da7b0389bc4e0c4a886b34dad3c47535f164e365c19f998e6b1ce3a0ef874b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee00d69997c3cf731157f794267390a7215aaafb46e9e24ec13e234e05f93edede7a281779e52e6a752480080aa8922ecfd1acf2f63445ea2798da87339188ad4f6181120496b9830b987acf309f627533b29567f542940be775c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f3f6a492445413002325b8b5ddcfa952a13f6f04b2e75f25653cc04ff51e0e2c937828092f505b566321d4279b6233e6fc2f4d7b36281c1eb25072ad13de875be11c8a1e96b5086755f306bb327c08faf5bc905d4519bba8a883d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae4c845c186231f6c9a2c17236d4d87593fee47449334b13166e64df529b8fc2d4fbc14cb4fda5db44da3fc59af4771a31983d6c49402c5a8abc370dee2301de03de86ff8c77ff4658210a2ea973517ea30b1b4737bcb7a2b2d6c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c9be4b58ed371166df6d8ca3f056fc430da6ac8761d6bff24f4ea264db21de177e01d5919e632c6a00cbab02c066eb4ece61e7cd67b494e212562d0e6d4689a3d0f003b5ce0bbe7f6e559c2fea417796d8aaa7e87247009d7a36f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c046b4bc727b1a74d721de7a7b5fd6031d9d50d49e1fbd37bbb38246368f16687f2d380bc464fa0e769d1ce0ad72b085ec683a5571b6e16351f250665d9357fe1cf50096fbc6cd31a0c82b47b24986c7db18624c247bb0946ef49d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6345e1fd91489bfa92d5db8bafb8d4ecedbda82d033fe95d55520294cf6477113b1b68b36fa067766a558162a4aec16d1a156560109305c1cbf48e2f4444ca6aef4bfc7a4e381c6dc5b021d3d9e003b5ee0c572ce032c55156ac41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4440757d7c40f0042cb600fa3ac99a9de40c9c6fb0f8b7e2bba135c3661bba9b1d037c0d928fb409a350938e608e93f364f361b84b7e135e13f30976c343a6daa97d6740b31ec8564c1141d3cc2c6070bafa5f13dd8b7263811d38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6af0e7f101d97234127cd8591e5b6b2479aeadc1ac5a48df40ebc4121af28ce59b72426d087ff6d00f72a54b2c806f19cb7615ce4e9a2fc5b241361380ec0e8530963f0b7fed1ed969de5bf7e870c9535e5613c8cd96b0c01f856a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde2f1b8e33d6ae8ac25fb482785c08cda7354e3da0b501fb04c78860733095a8e07c60ada7b01a682e1a1d74535ef254f3443a052a742eee66614377c8584f7030533706c64a049d7eed5d2d0257da89a835248d53e4a8406dfed9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he38985fae5377b1ccccdc38a4883cdb71325654713e91168c1ff3cece2b58d1d09fee30fe4a0cf413a330fd4292de0e4193b7816f6c4ff52846163c918d766e857f01605b814ed41f8a7612046889f04e32e84d0ea48531a07d932;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf093ff8ce118acaf77d8af20909754246e8b26344c273cdbbe5ae95b6a4f84101238a933b61162816663fd0bd1b00444dcc477a93cac57f8036c0d99fa8868127a2d8ee76fcd07c5a345f8f9b3af0066569a7faecbe056b78bf201;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fabb4503286266167b94cd49ffdbdbc3e65dcbec3ec57529391bebc761e0d7d8dcc5bc414364c497a7adf7140a3e670569156ba64f885b00fc4b418891915ac986ebd1ce05ea1e8ea7a0edc5b7944a9edb35ba4d76f1e910df261;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had137d82c0e2cf34a48b4cc4f30933fd0f0878e0d8643c438e3ec0bdc144bbd71630e142dbbdea380de58f2fc1ade1a1787c4a513f9bcb3bfad8fa92e511c2d75d6c3778791193e1088649a1579f9ba448118e1de74612c9678677;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7568018cc0ebf44f1599f31c4beea278c978b70231cd36adbe4ce129456d0726275a943fc5befcc3184f957b62b3064bf63db9a49f15462e47ad12ec1026a5e2ca614f90beb5dae7a3fd453d84d1ea17efb64cd3b63768d49cbccf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h865b001ea5f4c546ea89212885f6a6a6e55d0021ac9e386491b2474fa3d77e9329eaf496ca00d077f9b8b1ed883c3f41acbf6613d7e9512b71ad5c78e93f1583c6b49736612cffebf12bfe416af7e74451c259a1bfe77aa57b1168;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4786a5e26090bb9daeff7bf4765ea27825ae8e55df01a2c86273307918b16329e5234e7d7a0c93f34bf3b77efbbeb888ff477b9811e967635e54632bb39564e9f89e5c13aa7b61f4cd406fa2fc3f66f0fc2d4076da5445dc3f0f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef416c4d8df99be8255c7deeeb0d602b29d171035f1425d7ad2e0875636818c380b25a26011acaff26d9361f051d0ba9f19a7a80bb7f54bca0333c626fbaa6deb08c65abd36d8bdcdd0e157379a876eb48a2643674335ac32a4081;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112fdeb57d1ce2a3b3a33867aea92ce098bdbd92fdfdf695ebf00917d43a88d964f62652c0255743fd350f1d9983326ab694d4ab755279d091e50989009f63b76b2eea6b7f411c22c550506177fe48841f86fe3d17b144b89944352;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6ff623af78b257e4bc376d6bde1e8327bf4c2931b19d75553d0f904935a7817a0bbd147d3eec9d8bdf862804ac2d396fa32c8c0dfec2e876f312928f895c4038287d6cd323a2ed7bce4c8479ac6c2545dc7d9ed3e3d62a60fd2b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h309eedace434f533fc9f53c948bc775c08c7c0814a46d9b23ad36e6e0c262cd296928e242395032f9544714b7b76bae1d2f97abc28faa92865e217f97464f430bd9b31a82435df0015ce6ab41c40bae2a55a5a63736cf007536019;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14827c97a7a7c5fed428140ec311a2979f175386c3c79ffff84551242872468ac943ea2b24282e35c5915d6e72f09649014fc89b1bc41db4cc244492a011a154d9ed96ab2ffb5527b25c5d5ad806569f510784e68926949349e77c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9e1430026fc42fb866d967704cdc9306444082ec21677d2bafa79d66e0609a95b2dbb39c98beb750155dc149a8006e222a68ab2dc06b339ddc3c34cdbdaf57b9214548ea5e08dfcf630e7e60e9663be09f681b470dcc61f72ba74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbb9e89c6cb32a428d9526dacbf451b7e92db28e7fab5e10bacd37fb2e80e9987f71c7dc13090a3762c185e2b021487a56e131aa857d980a2388b8571d81d923200deb25e87abb8bbca61b40d4fec09b0f8bd4a94863f0a8e6498f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h640f85ee03d46264b2579f2de35ee92abe70780178722c15d3ae7431418703d65f37f32c15e91645fffd4e731a4fc6c3042d74dbbb32dd6773f55adb493012dbef0691542f050c78ed1479346c3c6013671ab9d467ec61f99b820f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ee322e79970eed802973be809774d443c548eaeb2e5706687f0e99db37720fc81566f4a430893e1488184d884da86e82a273078ed47f73ea7022f2e7efd01a47615cc1d0b7225aba072c25242d3aab4ab87feaf97ed274e6c5ded;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ee8fe04130cb762eb683f78ffb9f651933110032345e34f463af20506856feb892fa72122918ed7517a316c3ba0ed9990f5b497cdfdfc6c44b12a44f73e2a4bc66545ae8738d1533402ffc6092ffe3206ce9e555b78779d34a472;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e48e192f9e4d8583efb57312247a0249a291b02a2ae6ad02eaf080c016ebb68c6da2225f4c67f627a644b943c540fd5162f990ba61cf3860b0d8885f83306ab524a4cc7f347ee6294cbc0d6dce22df2eaa7c389bfa50bdeab2aa86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc4b74cf92c7b99422d3850073c34781bc546f5c6cd6131eb9f39c94906190960de34338b1269e124c8268bc4decea7363439cbbbb7508ae5fb9112c2feb238bbd697e500e9ea2b85d657ee83d630df951934c4fb8de41a3736c5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1776c1d18a2b68c9f64a885a3ca9f65e873f2ddef91e3dc610a6755f6aa07048574e2e26759403ca218dba1b15d2269a809c567f322eb1acd3f680c5f766abd40970956c346f738802514870931455461675a9d42745078cdcc0f6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he45e313898aab751051ed29c2e595e81d88b853f7031d08fa568ceeffe01b1c3d5b600afa31edf93b166109335d939073418775fb42d8aef80fb09c8ab29e468639cee0c9a50115c42cead6f06b40d4f19eabac3c830bd1207d36a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa6ac9e33ff0a791e683211efe8f9d7431e3ae338fb0ec09f0ca48b4f1256d2f0c049a3545e9dd97f731ff4785c1fa72b7ee1d40f3f7cd2fdfb60f007fd14aca60ae5e1c75bb56a9c011bddb8e4f4cfccc123ff1fee24f305271d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3f60377ecb4d01f8f5fede02cc0853acc1bc59a977e6d8dc1a1c2506fcef37bb79e51f5f465922a39cb07c0bcef2ca50e8559458c9c3afb47f9adaf1400317a5224f3e16a8daed067951e4086e7a8603ae32250abb1b9e9a55b9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5130d2dedf38d139e4aebf2762cec6d8c1ef3765685284045135da05d5f29cbcaf8ee2607d931a3c0292446ef30bfd2c15fb1e733180135e3ef8cfbe0645f16b4dab92c8679ff7d24e48ef4cd0ce6229a1d86558de3b150eff5fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5cf8dc04565dd13a23ab219c3b0fd194e48359e9495915d48378ff51c41c93699baf959812907579ea7beb15edcd6fb8c280d600696c24994542b83db622270b5756896f07ee3ae14494a86ede3e8e6b444a5456f41dbf568535f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57235b7d79a6436acc2df76b5c8bf00f723eb497055cd29fc065a600f6df52e6a2ca7b56159ff116e2c0eb7d21a7f2e337d802497061b91ee5abaf894366d15172f55d9c4f00fd54383fb2298caa261fdb0e1791c7defaba39ddb8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16a01d28d74d8a3151fb4f78ed013883105ffeca2d85c655d5f7a90d15fae92a98129a2810aaa0b3f17bf3f2a41ee41a1f0f5497bc4bd1e86766c6b1f0622eee0dabd2721f1342ddc097a93090a2f8c1881b86e32b2ee1de4c430b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c011a24e45fc7ea9218965d27efcb659815a346c8f1e5bc2e9cc2e9e3351fdcf855ab9887ccc9f39ab7982b78db5866ebc15b9e73d47e284316b745ef56d6e0518ab534ff54ffa90a63b4cffc0b33cdbaaf5710684d15f8ae7ce0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hffae8a8a25d86d9455b40bdbd6e906bf5128fa37e606c3ef23c1a8c130f1f1b03f2ee0314a62c008b4db830a9abcc34a8616dcf497db9d640b8551b6475948db675f95779d68ab57c663e65c3678dd1ff3aa63bd3779d0eedfb073;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h77f6ddd0ef3999d0d82a3e101e6f270bf181ae6243c3d02543c0d5f24a2d9de64f3ac1a926c970113604b6b2d9c5f353f273608318bc1f7a9f7261384855bbc8de89c578ac9c516817b15f56ada84be95f72c3dd123369d9016535;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ab8ce1a27fb84d27771a038c0309c88effcb3c3cd06af4191ea33d38093470b1a98ff2dcfaa6af92642eb7cab5bb9446314a205c9f05f0b80fdf5fae09497534ce13ff02e8f2922bda6b115785a3fee7966ed0125bca488771557;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2b1aadf34a8042cdcf4329ee0a5df8deb1a592ccdbe56aece76353569318985e4266970957a7c09d017bf3b26ca319b6d338cdb50cee0925ac8ab44bc61df5708bb0bf9f0b57c9e3d4cbd3c08fff1bf2c782bae0674d9887b704f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8253c4b4460d3018cd1e428c48c187199f8d2fd774b04c76f622f879b14b94c6dac599a62eaf3c0b089ffc2970b6e20073c48f02115d4f82ca9df9d2da8f122fed94934876a9d3d1dd515f5837fb0871500d8d34e231ceb686ebbc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a68a3de56dcaae7d828a3a0f7badf3a3f60f1c85ee78782e15dffc6fcc292701e67c514420157bc65230fbc1f575515ef8db8588315baebe18bd530a9ad951df03132a81c038c8e3f919021573df85b86ccc43efd957f9243bd24;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffc63422be14d5d990eb37c66c83581d98cbcb76183931fe9677e4c0b70bb369d343fcb176553f4fda1a62b2bc204ceab67f4a280015f80aedb61dbde1c05938410f09527313993c983ea12f60314941a1d0249951762f2f0b087f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9310cfadda4f7f47dd0de0023e24b2889766dc590964a9e1589c2c395cb3f0b2725abf9cd5d2c1c0e815899852d9c868625db18cc5807a04ccb7e552964ecfc0d52064cd585a73382b723ec4a864895c59db040093aad4d400687;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb727977ec0938fb5f77136eae4739f9822d8eba2cebeec5c40accdf2633905fa1f14a3e1d742a474e6a6247a971c7d20d5df296daff796ab888322d76881a79d3e3650a9cd649f5f8e3f84e8cfa1146590e7a62eea2e9aae864a39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb99ca372c40c175a370ee9a35b2e0881c4b57982e031d60719c528ccda2c995381adf706b29696343daa133d2df97a263a602c37fdd002059f82f9d77aa5350e3e4b16c89ce578632c3f02a105e13c66ecdd2c9669b01304cc837;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5415bd5f9c71d9ba12ec828a18a52167e3a432c807523651bf9ef5051b4c9f3f2203ef9f7143a4c5672502cf89c6c21aebdf1725f0d07d965349f6128c5ff88b580ecb36b92984f972094111f7ac7ef953185d511ba16088d42a64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63b9a39da5015162ea219e28adcff1fc614881f957d3a953f2cea8cf007a3837940a4f4a21b38e666b658484df34b9564c1d3b7bb3f04dcbe8c8bd12ae272b4906fd36ee9fe34ea110b83dac94d02963fd965f6c9338197ef08b9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1815063c910c94da565dae94186604787f1ce13c6d7ea136dc9c85e11ba0a532f4e9d6a04b6f67cb7321355436d5815ae81c60830771819763f458098b212a9e7f74713fd22e386b0dfd0bb73c5f7154beff54ae3dd70f435057387;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14860d2131d2ea86afa4595f92da5c61c4b64070b7276ae58f604caa5aa93c039d1073c336a33e3f560153c424903c7e06e8ca4ec64db792073cf17fca18f0cc2f34ab5e2bf791ecdf110174a8af02963638459ef5e3778e65fd328;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1710dd84029b57a3b2021b59d06fa8ab1b9d5d978277e05f8beb4fcb1042270e41ead3679433f7c06618266632ff705c420be83993804bd9564ab20d058e6d221c2a72768b9edb2ca04da47ed11a8aad6296604f9d9319acfac2e56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f1ae7b62d64be09ac9aed90705f92cd42af24974697c293533860acf862e6e03d2aca0bee1771f2381cc4f542fae2dc0a759a61f97816a3634331a97606bda30cf41d82e26d810540ecb4ece939378f84b194251eb0587e1124a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb90d2b825fe0b5919aaa4c1c71365fae3b855b6993c271cb23d433c9b83b68fc7649fb2f1e27d406d6a23192efb94a639e66551cf3baf9142ef3ddcd14fbf9075edf10cd7add85f26960f1245e3775fad504f3823bcc0c9a670dc9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1480ebcd7e8f4737c7e91abd3c319a38945fe952d9f8f3ad33a82b2af1dd39bc65f9901b9e16821998829206a540ee0ddd5a95992f0c3d819acda0bd0147d853b6519cbaa4df9356b3dfa3138a26694177c6467879219de245343;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbba42b1a3549f90df67b800eb7b3ce38c63d91ae14aaa0f2815988c5381208f98c77405d19d5dfa9eaea2a96b68ef7378ebdcf7f481a73b8d5265e8dbd731ba401ca892a3e8f552510bdcaba950cb435918388db9323d86e1520e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc847f7cedd2563715a923e3b61b13777912f713fe7bbfb60ceeb3896815de6feebecf51ff20f3d1fbdd009da23ce6b5c9728da67820fef34471fac819692aa6c9c79f0c9ac671173d15c70842d3a56ff252d9ecb308bee8c9005f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf55564ea6444b1b0e1a8390667a0ba795cb181c92823a13623bd3715e15d632b2a1a7d98293749237f5fbaac441bceffe1228488520644b5473d217f3cb29eb16d945be3a0592ca19ec8a7a5fcbc7f36b8caf502df1c2a6a6c93b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd1bd70c927eb73fa2b7678c996524ea5c9024f63886e7ce45faae2f347fc1ca3e22c9d2bc958d4ec6e59bc07d32ea03d7a6a890e44c5ac52ece0efe177f0c8cb2d1acd637dc338ced1b66fcc7f5b3ce4edd6490a7c1567a70b289;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9d1e8fb95d5b5ba91250ba7ff1c3ec60d71d0c16b785406f7b560ecf687adab5dc847449eeee8eee139f636dd7f86916cd664a99ee43033c8e1efdbca524c1ccd832149a6efb0e2864406ae236eb749ed25b1457c19a87cc2d452;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3794233ac84262e0a9605466b119b6d9969d4cddd44ad0e2e2e4058e2914201baa40f3beefd6dbe50a4da83a0d70d1f498b975801605140a7dac74d5d28a2bc7bac885109e16afb594dd3ecb503d5cfe7b114e5a784c7e2755600;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1193451afec7944d36d3ed5fa837fce7d89ee8dd1ff13ef257af38de80b8e0302e0899f03df3d512bf8a1cb2cedddc37ba53b80b191520f9428b71277a988212309ab1a95dc52919da20415c98f769c5555f1809aa36e5ddb3e8204;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he161e7be1143244d613c285a92e60806a92ff376d2d0911c2afa075524d80d815b0a45dcae645902cac81fc29b1759379ee48970e39e002c2f3f3c74adc3bd3386a8a42b1c243acc78084ffb10198b67625b5af1a22054ccfabca6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e2e9d22292d303eb862a0eee0b454a2a14883b47d22cd54a2a6d702d22deb4ca8756d4bd6ed74562b05e27fe331142219861ef07c82d782024ac7da323692d718e39a6a1d017f04fab5b5026859e4ca1113fcf98ba7d1067af86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1816ee83866377dc961570d1271afb823d000b8f5e0afa9e525ed1e273c79ddcf9046c84e0f9a121276ee45bf1361c9786032fddc3eda2758fa4775b785d45baf9749897450bbea9ee30de0858182688ede44ea92203bf53e195a18;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197e9d7cf1778a1dccd1da1038e87a122942207369e73dd871dc0a2ddb1d1aa2cd04e081dc64f46ee9b05e024c056d9754761db1890d578e7b103d0c38f2e44f83e192d595d8acf2df1a1c26a899127a15e2d119a90667fb48975d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95ba8024677d3e4ff410ff9dbf37ed4613d22bc87bc49f88a701472409bc86d5ae400463175da5b4a9fbbe2793cc33264ba2a0e08b527e8feea034cbf4fcd947172c9b28d122a0815cbd27ae1bf12a550932bb984ed0214fb7d9aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2eba41755aaf9d6d5d680e9e35708a2f11ef4d3e304de0669775eff08f8b221a65feca02e0348dc393483716dad54122a6ab3ff9354106073979829832f5ac3f024c7c5609a57b8f22cb39272c3552374c23c0b42c9235ee6697d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1aa826a7304c1bd298afddb3463db9023c6210dea1a90dfb1a29c5f6f25fb231edeeead808e66570d32de8cd57311f24ed61bfe91a770e66de4e46aa1152cdf3aa17d5f6bed8c0b8c2b90b684e0175cfd9116f7d5a64e9a8cb88;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ee4b8fd4518b8c01db5f978803e4fb88557baa2771701c6f7ac18fe25d407ec6796e20f4857208029a471d7f9836398360fea49821c143064bcf5a6674708d2b15e89d07c572eda1117efb77250897703145a7b6e48d067df89f9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d3d9d0bff9165746704aee813457079ba5ec385d5a053534bba6120ed6ec97fa027a1189473b90806da7e448abaef9b2f80694455811f7a7e8a2674453421f169866e420c1b1e2b496a2ba6c235a31afdf540d6ac07d94274ae45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1964829513a085408dad5bfff91d17b893a814238ea8cdea9f049588f1fc05866beb92c4e1f651381b9f7cacda17c199509d3ad934c904614876449ea38fe91a747e14559533c066a0492d9368b6395aa1925ac522507584accbd69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c77be6232b94f301d885e60d7395e52b1a2e4ae4c17fe4a3d51bb37ec28ee165125c287dd04079256066d7523d7979fdb77ea33d4d696c6c030b3f1cbfc5dbfa45e07627a0905a6adf42059874496d65f882ec75f15a697665fe04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5142a2ebbae6a714007591189a9c6dbcbf4288305de90ddbee90b127dc3b688789b0683d48595e824b168f83601c8e9613cdd9e19e9a9942ff67b71e4e93e1ae5e2aa1cd3ba25a713404ac7394f3ec13845215c5c2317d4809f7e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19651e9f00e48a53ee3f0411ef940f5e8619a8edafa314e391c933ed6f476ab3d1abc7290e51ff4643cf177ec01ff66bd438516e1ea9f5bc67edf85e031a00aadc6ae07b186197c5a4977d860153952fd3302e865087b482813b2d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h195ab019fc589584527d066a4751e0b7cdde565c54c695c03a6922859413f2831ac18cd5d914aa99f48ee5fd746798ad924ca83880d33fdf55ff614013b0da708e0e1b86c527faf1a1ca9171565465794f34b9d50e11d11781c74c6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12714ff9208705e8df385f12b15a19f3136f6cf5067f6ac4c13c6e781bd7bab466f93d603b73c0e8f3e0a68b17371fa7cbef2efbc4a7a2433a49f89ed446ea9bcdb73557ff0184aa629aa6bd26e5658473044b240d9e457f50ec4f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b69a52789f04fd61a91003cc1b0f34d258ccbb107ec5f2bb9d2f93d4bb8b330ad69191cfe7be0567f628d430f10f42a8018a9e19f815e4ad9845b8b01bd28d57191470b532ff93de827eb69b1558707126cea1f70011d7c2cbd2ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a503b6d459d5eeeaad1e976301596e4eef810e6ebb04b359e74ef2d232f45bfb459998ba153727ebae5f5ac436dc8c33ac78b777cbd3b3d9f75514ef88575fddc5a90c976bacbcdfe7b9013066859f52de4770f0164ee43a180bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f17e7c3b238599a323200bf21eca98e35e9513a58e8a25238b29d6fa3f42568b7fbea8fc98af21eca2f36f63ba2881bb0a507d14eb99561953834b97a0f6e929f0d54430f614d51f41a721c179239f609e099c683b345d1850f9dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db9933e8baa4d6e504378b86e458a20c1c7eb6828cb2409093f5ac13a1d06d17243aee5fc9af4dea47c9dca08002c0a8bb69ea49f73da0e21a1c6b14e931b71b0c1286fb7a5db49d947159c95bf257a77280bdd4e62033751e52f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h880956c670bce7f41ff5c3db98e66940efe49b95b0b42f6c35b83d162f1d96558be2f7434e38279dc34358b992c9a1f1b680ecfc2d5121e8ec5fc29dd41a62c41a9451835ce430f206e283da5361dd74a93ea78ebd6bf865eab7d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1789e5b0acdaa9d85e4b7aa94656c5669a5215e1bc149414cace555e38b40b71a1dbc7369c456321d94135c4439422f37438cba7704774048f9adc3caedbfa00f6c2f6a21ab515208d9f3d4f22665a0f564fe952224923b31ad9987;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b438faea3daac0b417fcdc096b6ad9b3b63d9fa3c89e240d4e3e56984f666cdfae74636e33d327f3357efd8a40af7ae7d7230a0f1ac7420309651c1a3512cc828e5bdd999e5c074f4e86daf5138b5fc92fd8d07b2895fadc20b8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d7c50e139929605379b1669fb510471d0345e8a35a19ac804dc922b0b78ffbfaeb15d17a4bf367431369e501046a40b3b2771b331efe821aceecd76420caeeb8173cb3be9089d7aea5b8524491963264e849d2be05c67545ae48b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h482510a4c19e776f56f5b059938b643638147b4973fb9805a7f9b9df8435e7cb2405cbe44bf0d6dad79b5c67c1f3611ee5cedb21b1ad6a0f0cf2c59a3cb700a2390fd5684854a29352d3a7badd4be17f0b17b27cc904f65600a32a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5a6082ab70cab38f664e4d5a32d202e22dcfe18e9489be12672ec58b2a0553f8d183a24a4fee288b65f7fabd17ddd2d9ee6a96b09482e82c78795d86716847dc6f8e0d6f26cab36a9ead2c3b05e75a83cc31adecff5482fc1e427;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1274b61167ee8cc9a8d008fcef07a99dcea1689f603702699015ac765242b76560618e1f546f9de38c15f6a54b2515b11a32474b6f515cbeab891faf371bcb7114a6f08ff5a8fe2ed69afeb72950c124669a944b044c6bfca2e9e3a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45d5952786523713afd1dd9deed9fafb75a40f77543a44a645744482fcd72e847ed3db20d505f8acc197c6525895b283051f0f147009ef11a89d393d82248d43e74f14213187930dc779b826b014985ef3536463894cb530163c0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76c5c75fb7ee68288905c5539af3a0358e1d3e4afaae7d0f54452793282a1a0f2a7d2de424592b6d1407764d0a23682a977764ee4e83c675735bd4c394f655d2cc28a38139cf786b00889c4c8039bc0c30fb53b967a31aa628fc71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10007da9a0bed01d333d9e8c4f784cfa75141318ead3ecf6a6013dbd9bf691fcb8ee079d79abda09acad667e241b61ecba77a237d750698306b77aa6f68650f842bca7fb73c3aad6bc05512d0e9f4e9a44888dbaa41078eeb38fff2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf0e2a6da8193456ee1e863bfb92bac00cd550f7c237b229db7845c5aba97547b083a02608677a411a6a68749cda63832948c63868f490459a8e09c136042600a7ca6f7dfcafad4f8650375bee1b57c78402d6c4a77ce1d6a73589c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca14a484c78b3586faf1a187f0f723bcca95676d30fde74cf4707506f2ac8f43bc3fdc227d9122c6e3f271dae006cca5b250a0d9ea5105e6cd2d6ecbbb13f07818fadc55dfda62525acd25e986ae0eec22e8e9e0dbb1065331200;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h161d866895fe065544932f0d1425fa4cf30ef6df31d2608b835df56d56492e57dbcd107c2651e19b6d561c2fa22b32d0ba731e6e1c044c61d2337cac4ffedf32a2d808ece4d131784f205c82261923c996b55a966e6f04d4415176;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f1697ed9567718f901551dd66ca4ad7fa429ca5d5496067a68748c12b76d7c15ec39493aec30e1ec955099026d7f20107b8719e7926c0b37e466d58774f0d9130532a5c8e96d67cc68a321b5e7c376da63c49577ed9281ddc974a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be34bd36dd42f13bd330c731f58c32f2c846c43789c2389ce6617f911a1a34e38419ee9a9369e7ab5620d34bbb4d9736ae239eb48033bd6df4bb70b2a55a61b05389da11a7a1f4d4c5a4e767294cf0443b578539b5937ce16bb404;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc493228e95bf090ad4de027142012a924128b7fdd7612ecd8b1aeb9f508563b653e4161967f78e7529a542221572e519bace28e4579031f0deebc9e0745b89a2d378703527407c082df4101443bc65da7e4597cbfe061356b4ea56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d52ac2b0da456b382e56a97c5e06e08df7d0c31c70c97099d12c6fe04e4357c6262caf92fe92f1efa0473629b2da2855a97a3d80aa738e2d4cc95063033a8f5654d688b606c1d8cc556026c821e2e00fac6db82849204bed592b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160990b437807cbcc98cac1091ea4e161c1600f2ed7870b1c6e25eb046fe8ad1391352d952472c6f5575b79abd6d903dbd2fe3e52c96ad5bf0bb8155dc2768bb3b45d3bababd0f5d7cb37573fbf086e9b7731562fb2f332ebcb105a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h899ae1c6cdf62880e6e38ed92635b31d123069d3ae66e8ffb640d318677023a551b3d837bd7aab90041f79736f2086e28bda0f91a45e1a67aef0c72ca9a0ca15418539fc693a1732277f21e1a52968593590e73479b94528bfc681;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ba1d1625a61464aae948a82bcd60acf1ec88da148071c9ae68d9fd01fc4b176c7a2909f107a7f920c082e77a5ad960f8cb374543a64a8cfb146d1f581498a6b26f54a339ae543145032fb74144a6c4a1948e7d07baf29eaed706d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4c52a8f087edd2693074f99fa7f52f2abfd2607109e3f5d3e54d68a7da9ce5e3318c49bf69afe5deddaaf9c85be3eaf7377cc96ebd903ac412ac9236f1e11cf17885331dfbd21d90abfd4ca21d405a6b8f6cc6dfc1f9f4db966ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c46b40205b95297fee63fef4557a79ef254a495f14792d53e32ca115932d4f3c88745d7bdfb154bec5723c6de75b194851ff16dab09c05f8137a6c421889453c50ac609a5836a900a56d2fddf9ce16117981abcd8099fafb390cb6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h949917a7499dda77680f404a3dd19623b34a4253727d2ce8230912e649fb215bda55fde5c354d9f55fe632d44b1370c6b40480bb1ec5630bfa7b9c06bc7a80d151d128c244616c0f741c0158db2e28fc7c42f569f5e21e7b2c9666;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172bb8e034f9f8bd2a3f9656158e955625d3ba1ccc777b213597736d52bc161096b9b679dbde82963be85fc384065881bac3cb7661709e60c7ee51564d461febe3c2679e8c7da40017655bef7e91507464a716da65bc7db7e2cc3fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173bc4a3581330e656ad7e3fef4d55d8f5270fbe8e2ffa49852e46c0d085a3e5211030cfe7963d8950afb35670b14709d8dde6545b05d9f2dd0e03452e1bdfd4528bd385c7a220a68de1b0da924cfe710d46ff0de6d3190b3ae0a27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a25b24cfe6957aa0d868fa6c6b39a83ffaaed2dbab937a6f9fa9776c1c9d36d607135f26b3ab561433c51edc3c283350ff5da49bd0deae061869fd4c817ad0b6e3993722e500c6c9a863c58324a4dcae5deb9ae6c536c36d5d0ffc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5f7d03730404160555bfac7a6fc13aee5ab32dbd402e1a75e00de7b1ccea86b5a8af8ae0643736113ef95b6fdd7a11b4514b14e0d7f69cc4d61ad7fad337e7c5ac10c1ec894ca59b0734ce402fe77932d6f45d828a568140df809;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121c52ab35ac588e2807c155ef77a9e4e05b9e6d789a0fd24a260dc1e6650735ab4263a3a0df4762ed4e1809ba2698144cd0887c0f699c14f0d4abaad13aeaa8932f3cdce8587021a488982c4be45fdf2927c73ce62bdc2b4cb5953;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dceaea8bf2fe91debfcec8bbe0276eb6be9e4492e2ae13abd613c58861f6a912d0c697a6929fcdabf3d04a38b3702d76647df5b7c6049759902b8aecc1e5b8a1fd0d78f90c0aed59c8fbd7746fc9fe18efb28b9a4f8f8830a1d6d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb69346beb562dcc0e686de3c2809ce869505c903e4bf25de8499781fd9ebcd1f92587479807405337430a3f11a5a780cf5ee784dc2d67ffc325a14aa89787828f42ffabe92fb77ec12b63bbe46af2bf30c2105a9d31b70c69df422;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc663d2c9fd7b2d70f961daaa3bf587695f7d076cee7dcec7a9d74465934f6a55f3d3666d8e6b2ea8a6e40d063db778c151bf16d4b88abd140d0b9480ebf2380769f86c86191056db59fd3147c5b1183255747981e0661978949772;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfdc61420c6a99492ee5d53beea7801c5d44eaacd0192d7d08b69b287626f2a56b1a037e36fcd872178eb72a0b3119a4fa1975698f3cb5913fa7178e5b2f579ba5c8026f2e984d0e28c9d3235fc6861e6678d7a1c240984784f4353;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h337b6ec1162c366b738369aaf1ef9a2a8f3ef0b967523c54d23952025e54647d12cbe0a4d81e3a2bbafb9befb817ab182a98ce12c1bad228a03fb6e1458112d0ec326079afde9dded821640735c1f418872add7a2fcf6e9ef32578;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184d7304cd3706905c4d8ea75667627843a421f2d4300ffbb41b5fb9b833e0d695e71b84f8612d46f38d06080081126a694450be25583d457884ddb4c35482e18e0f53b7db7145f0a0295493e72c95563d7e2723f3c1c703f8f74b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb2f66016d6b13dbc1c780d28dfb56d230a55de77fb9629f29714d6785ecf6f5766451e46bfddaa3ff1b61627d588d5e095fe5e42e2b260509d9377776449be79df560f325e88031c9e80340cf80fa627b179bb77b3d2500e9c738;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53273e3cc163a134c485d33cbba3b5376d8a65a11e0883c6562e95d0dff0ae2a5b812b9a4e9173f5fc307443f00ffdc03a472513bbd6412ae348df7d0a6e78a946c53a8955fc32f014014f751daedc44993a8c55278e8627ea6e7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b359925a183713d21086f8130835c4c316ec06585a08c8050c54b7a5670626022b758541bfed86c2c349a38eef554ed426a4975481272a03cb0349c1c232c75c02f77b720ecb14f5a54840a0df3eb543fd5e3fae228adc6b8ce27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d9322312d366aa8a0e8c63be83c511b57ee0ae989c338f2e8776d7ab271053cfbc663d3a02ac90ba6109e3397440adbc5c263b5c0a5177eeec2c1cd867cd64270d59f2076cdb8ee162dc04115f8c2cbf268604566ee93a15c8008;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c694c2124a8859c4f8a3953cb2f3d5a9792ce63a91cced3f72d9e57208c561d50f027021270cb547e4004579e26971cc308413c37b3082323fa8051c23867c67c0da66164fe861b6a1d5fb97ac382c9cda1ab6f42ac61b1c217ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13be4b209aca750e1dfe518efd6cfebe1578b5e4df10227495bceca78e7a0aba03d630dde87d7fae280c201c82b90ad1e2de02b016a7e92482e492f20bb42547157c0c3a015405bbafaa3b0e7704e17cf61b81b0a5d62090d522ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1788b193eda72026d34d66ad1258ab93457625e022691318dd055188253629dab967507ca4c69ff0ce63ce25689e04f32fb5c8f3810dbed8e2013079c476e6e72f44888583c71ba11a7086beb2d1d680b42bd60eca4333777271f8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34065a9fb4e5851134bc3a7542bf1106d3726f5f7b86454fdf3cd7b8d1f3980c5b775f41bb044d067c5aa5c380050a4d28dd975c696b539196440ae5c71f728dcaa89de5c23faa3e3a7592bfa7b9473c9b48f31dc42c9324e80909;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc6556c5156823e27c298875a1bd80bd4af70c4f34fcc008e0fcee4e4083a1f52cd3633435b331f2cfe9184ce0660e3e900f4a9aa9d24fc37798fb54c07ebf96735db9b8329b387e73a6fbf0d9a59f2566ca1be86d9a018d747d04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e21c4fd7af23f86486100be3fdb952639bbcac77d00c0a0d9055a14ca4874f06c98123de7e0167b9cc902889f11eece540bc2da1a731831c4a9de8920a3dd7cb27c36d14d816417de7d093922e8b16c07c553701729b71946097a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b72c76f82f60b1b81fa13ba7968469639f9007e7ccbf7bb3243ae24b8b9a0b8a9c07a3a2c5d3db9877f790a4baf672e7a833198e529397f3ee5830ee35bb785ad5c33dbeefb6e133e8a45304d6f27132ce60bd1889c9c387a11994;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h756d3cb1525f5a48b9279eaa8805626f66fd51f6dc52a99a8323b7f1f5c1e64fd09b0f07ef92b2be9e5fd98ed15cb8fc4ddde73ac1ae8d00c55e3379eb043e3071508570c63215e40b9607c4473ba40abb5d3e9fca1a0920b0a2af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16eef822b7357511d4088fab8922c13570e39665bebafea72c723ff8b4068c5502e04604f643dd6d6a528db89a73187b84ef2fd90ea89cc0530cb577bd06088a14c47151d70199581637cf171e34f6597eeaf546ec3d2248c11e95f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5cb3839c717a3c32a495d200d1094d61f41e66565065247a0e8c961ac7e8cc673d8431f88d3cb62d8a9e1847ee6745287e7358a57ad772a604d57e06613580b2f0096b3fbd248e5ea2f011d9575b68517e5acf53f00e323b545e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1cb2692bf3e6d379d9bc6c7fc65646b2e06ec7b03c3767c142e3949c4f6e6c0dd4aab4889778af595a33eb64affe83284ed31811c54083d6040f18b44664d8bd46f90beb208e793810a37e38648a1c19625d7e32b73c07c4586a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12166ab5a2972bfbb3b9bdd13188d035a779b4ae597baa81ca59c080cd5a8a18a845bbc3cb536fb3bad6b3143b89c24f484ac215c858a6339385995b0582b287f6e614bed41bed09d9570ff9132eb9d105eecc8c2d9b2443e8f3213;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91791a26d436b04fa3b97b6aea39379253a4cb8af0bfc247246e2086ada255533e164d26ee86d6192db17141f4a9139761c7dd09e1e893dd995685a25f5b9978e3d384f7dab69e4a9862d34c1c9106d264810f951866ee77d53e19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2f32f1333a6348706c4127c97324b160fde6b4e5f57f236b6ecaa898b501cf465c2c7d358e4ae8ce0930e23c152ee114d2a56c42ed000f5c63a52c3658a563f8c0b8a6f7e1d53c453920837ef7edc70a058f080c3447a72e85bb6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb19031ba1087d58ea02f53f86de0d85ae5eac422b19bce467dc8b8408c7cb60605c984bef811c252d14989aab98c74b863f1661b98fa82be0a03c20922047f1c2302d005ef189b9f0727c4303bfa327d65c56201ad5b2c9564fb3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45648be5673f9391bcf4525bb0ca7895d7e94415b34d43aa3417670e60e4c1ca01d666ba683df6f46b618fca950bb413333e4b3d9ce26614f8b958918de0d9ebab17b57ea59f1038e1b79ac483b3cfc375c4e37824644984680487;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca871fa0afcd39d1b45a99a24b9e3d47b4392db63901a2685a16305461b0dbf499c52f9167ebe3a0ef00d68080a7e2ceb1f985d0e336413e4477e7d46cca9918a2c4a51be4c14a2dbf843b60df176f4d3fb4cc121768b6de7fc402;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b8282255f8f65ce4cbb78c1167ee872df2f3e30524a4ad1c5ab4df7adb09e2dae054c339361f7f964d17764d421a0021ba6a400f01de006558075358018c71d8d8491ccb9aa37b7b012619e56237bf11439c751459bae8728c86d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8807f101d20ec86955dbe7c72a2f3cb83f9108b033c12394bf0616a463e9ee9cd8666a59d5af7ff4d31434219db30000b145c871b2159187eae361d8ffa2b58adee41c74d3177194d301f0b49a4a66d986c9197e324047ca142f07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dfde9fde19d95310be76d107bacf30706f8dda93ee1df68c95fc83a5e14973c21eb0a5986529a6db09f40a3b442ba94cf00c14a48ad1a29599998665f02e654844fd413e0fefcb16f34c147c356c46303db7fa998af07ce4ab4a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24c4c0fd5abf9f0c947cedbc36cfb3ded3c2e7938ffb60361781b9bcf5f78aacae5d8b36bf02bb4d68d733d9c437ba807fcbb1d75d1c46e628d61a3a41e0fd60927ce5180000ecaef9fc7692e324919b27f87a93191e955f6a4eda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1125c2b6754aeb95ec522174dd6e2377e55ee57e0137c4337a51a69e1c787acf5283c0d428d07f06a38f6cee1f7aa4c87b9493a9ed1bff0b71dcb227414d0bebbca1b7675fac8a1dc7f32a9d98e03387b7c1f29c0bc7d7c11b79788;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f089e0fa0a7c0c2b4ecd4e07d5f44d1ed03ac6e9a38b65a0cad9ca2d9de6ad12611be697ccd4eb86b5cd6d40b3cd814211bac55d828210b6eccbf3576e0ce861bd27bf93fccc23a6fecb6c231200f68b6981ee2eb1579fa697e8b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182dd1d0d028a99a2a8f997b843186b238de1bae38c755e1b0ba37a94b425dc29262eebc5f233e762ccb10d3c081bcb490fd8d421c4ef623fc8655752569d115f958ffbd141bd05f02fa5b280cc6cf02e83279a930d82a102dee1f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a0458bcf17bfb17718382564c9abce9b651e078c823cca6fe2c6dd566314be5c610d79c7c5228d273716b87d5da7fdd8346ee3e92927e749fe7ae7959359ae2b35554f85ba9bb5c8df286e1bded8a8c9e7188a835a76eb6f20d25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57ee38b570f0557c58ece925796cd3cc649151f0255371a664ae9bbffba04e2096dded17af4e88ade63219efaf87a0d20c25d9d867a2edadbeee965cfc00a655a967094826e3bd697ddf5e4dd361dbc1563f658940c56a739fa471;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf51b9f180cc794682664dae7cb08f4c01f8e91637881b9d7831212b30945efe150c6a61dcf6f6c3d743527da33a0071c3e73dd8c5f36dd7afd0f2bab17920489b667fb2217d97539bfe7dce827252c95184625a1d6e298b042ec2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58037d7bc91b2409415849437bb227d33211d51a7e1cd4807b996e30f6100554aad98d4d99e9bfe597e9529211194cc55f416edc96681ac24aff5852c75ddfc764024c3bb0079d67b9962c8ba2bbd0bff1dbc8a648b40a87469c19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d71bb3d7c7189344be750fa1f189421a9e17528312a01546c128369dc433ed8fb5bafd86d61a7ece3defb494bb5e57132120ef912004a3fe17b5c8d25307242a34f4d3113052c76b70dd164a6e46fea54fffa022597378e68bd4a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1469174025842b959794c311284f8e5a62faf0f7a567db7b23f861144df8d308f291215f17d652881b7aeac7409c770def7adf4ac4c1b54a9fa18ee331784c2ba91fa1346da27ad5e85cdb7da9b7e9af70e62d04876da147254f4b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188159ffb6175b6b2146c94371cd4937210a3216b87a4412f6ddc5a7eeedc20dadce583d55b13ab7c250689db093e164508dffa441c267683434f23793d1416e325689a6687d0d6eb2152b88aa25828233bf8b4181d2ad498914d66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa5abf4a8cf87852db0e7f97ea0f11f14ded5f9a939ff943e8de9e0b8ef89596a34d1f4636a4aae0f466c73c97f3b9ee9570d00743b4bd1130f2dcb080470cdca8493f1b9bec70ab9f571bf379f0de49bf55af18f26236c1ddb2d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99a257b90b7268b57071c30de905edd5108e381844f20278a7651e14ce228419a7c21b2f387404d31ef2bdc472f2144ab81e7eddf33588faa5618d795ac31017daf01ad436284309a43726813eaa45d9a0451b4199725420554085;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2671b8a6a0361388a539097c2f5ff3275ce168ad852da216a02c3e772af436ed5148836a36c5c02117a40eff789923a258d6b307cf60d80fa6bb2d53a8b4a9a4ecadfab1a67aa324c44a46926730666699fca651f18ef230b62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d55b714abe4cfd832b189a1b560c7cd50af0610dc5358d0e43afc861899bf4baf3adff5a2971d6944682f7888c5704888f3323491a7546ae325b9d834d046cd927ea750191d45e34b1ccafcfa0430574a0d13715fdce3a0529f3f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf6b8a0261cfbf3efe0eceeae285e4fb2c4fe6d05c29c3effe7fb80596684a169ece9568177c969fef8063690d8957c6696c7de980d1c6825c03c1e5328fea3e13fdcfda612f4648ce52d3c33bd58a3efba00c55218da6cdcc548c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81a139c9a1eec015829e569c75aabad910a4f9ec000bded1f2b4a082117642b9c41393b6383d25cfd07e42dc2933614f3d2da6cfeda0d1e98ec8cb2e9c8b927d3e4033a9df4176a73a07a611505e04b875d31d22fb2265db0f9986;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f18c2e8b4cad32b83e9f071eafa7f593054313d5db253ee89fb2c1457a9aab7d88391c6bacff5d7ad5b42de2f2371712a7048b682f0e5f08bdd0ae316db2af38fa5f3e444ce614880f9b6dd086b479e1956484bcc1e9b2d9b61a1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ff635c2cc3e8aa77d62ffbf333483766f2059d2f38995653289327b16fb9cd021bb5c7c4488ef3a674cbbecb95a36188603e7c92e7b935029d8cfef95afcc74535f7c7dbb8ddc540d5bfbd785844b85384f90d5ae891c8793c614;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42c6a171eb7f8a6e3bddbee5d1e36fea28ad061bda52b3433af07eee23f081bb8753fc92db627f7da7ab5eac303955fce8bd020d4c4082ed7f2af169bbaca177ce0c11352c81f8d88af0fe37fafe4cbe5be790d11433a6be6ad171;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41ae2c3e770fbfd343a4dc55fbd2a57d22ef705f039ddefac87f3b3b36896c9834490dce1a8af36ea7986f9d994c1c8e91a45dc72c99abf040d29f6e9932919e0c64f12fe12b0befe35b4c24db030807cd741135fcc1cf727e6656;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec04f00900a642ff097bb7a1b4f3ab5d27670f2076e91164f345e383755ec5a2ec852d95bb0b04fa74067e6a5cf6afe3ca0485151596db6e2f86b281e43483be0c45a729633ea5884ce3af7c2a799fbee2236573767ed77453641a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15af087b58537b730e9174bae2c3fee599039e1f25cc18266afc32e00b2e89ec1b0a2d87c97fe4fd09f3287739d65ebf6a3e8a2a940f092971e5bf4db3c66276d253668fa3d9650bcdaa6ff487d4b97c3c91477944f360a42145644;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f168db49fc068b1dd4505f4b5c2c64d8367688d100db9d4907f48c855500419fc62110e6b4e17c6a31764ccad6237e533a204df5f662bd492dfac470f33d6d666fb8a5fd6d5d3a44e91a6958d495c91c2c7f81be06f53edcf2f34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131ad700918a0fe5e03fa6c75af2af2374346429b0e6eda714efb12e2493c457e0af227a1e78c54709f6050b11ca9acc0a45b7e6ec05a83c53841177cbbb29086e6cf2ad4f6e07e6a37cd135775ee1a1d5a49d984fd52f344b2328f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e5620327be7880b1e046eadd5ae40d5bd2c2075248c22355042f8e8162a0c610611084ea6c398866440f1e436f58c7e06ddfeb14e5f17ba5fd64ccc5ee6b375855883fb44eaf8fcfd45fb8c30bf98de524e43284127c28c7a0db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172d9a8843b5cc85bade18ab94f2be9d9242b8b019473a7dde881b31a5d77010e59916790f61fc3a56e3aa8cd9fed8ca8d0e6fc656b04b2d96b3e4978ea4cc93d2c8f6493f9d3509c5b9770ccf8c51090934044db720e6021ba7f7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2ef2eee63d392256d5d710cd5518ab775f1924c97a35f55663a58ad5a7d5c8b71228153a090d4f45ba3221c69f2042e0592f857821fc1cd540ceb6b1bc887753e9e3cd6ec62db976b289e4486c5debb403d5949b9aaeb77dfb10c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c48cd1c20bcbfb89153d491065532a1440765a29f14ab1b92a02b081771141ef8a5f80ca68661d5ac0dcc3410b9bfb40e98600b176485a5056ab72032bea2fa3a13021ae018e2125f3519056d9e92d9f60652e9eba8dffc512af63;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf2b44c9da13c9f3877fd22e4c16da6949aec8d539a8fe246872d0482d31e397669c368ce32819fe310fd39bf3d7289593abc07672f74700b026af87f2beca787e1c69c38e1cbd5ebca631adc408b8fd2fd95d40ac2bd98a3198b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1caac3b7039a6f9a3715865fd3b66d204bc3cdb54fa293e8dae95dc127e1486f42ccd47a8e7de5ea0ddcf7e9113e8c843ae8106282c6a527d4c6cac31a6c68829425ec7a1bc4237ecd7c6962c3c1437088fb820c162706e00746d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152f620d3d2dee4fc6dcefa0c6144372af2f2023c974df7741535f0c010e156edeea534d52f3c840472e54950414c39c966c2f718bd4a9a67de7c18b2b71eb60ffe4b426959bb884453504befcea2bd3d4c1b2cb8e8783528223a72;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a332d56bf04ccaa4408c1fbc9829133c43dd83e106d7189684e7d4036caac58d648a55a526779fb56e6e6f82f8452f5d0795b0cf9eeab2cab660d32d6a633f18892ec87b034e43930b78334d3be860c7dfab29e16a8a641efc4304;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9ee5d378747883836f79c899c97246524f49f9e8c16f48390db7713ff77385349c9a2382c6fc1b40cf1eb885102a04a97cb042a89b4f906a4b88da2ec50155d9f83955002bb4730ecef1b22512de48bdc9189650fcf2b9e3e2501;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h367ebdbecbb287a31276c0c76f7d48b99a9b2f7d65b0d159f6110d299536715b4a95c19f71769ad22eda0a9e5bf1ee057a74d130a954aa0dc218b45a45480cf9004a665c4c6f97bfacccd20bf00fc274b18df9928aaa96991d0181;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1bfdb2003874e5b714c046eaeca1a185caeb9f03cfaf84e08d5054503c3b7da808982c5f3a2939fea9c47126b1d949cadcd5d1f2dfd33cbecb35ee3dc2983692d73b723893b381f247d7caf9472a20a6149733a821bdcbb829b84;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb2f65fdadaa71fb5df414acc009cfd4d8873e56e0b0a362d8eb4306d710078852265c12e31b2f7c9cc32bf2088561d8fb31c2f9db0115100d19d77603e989c0cdbe74a6e70268fd8f4d6f02341ec8727bb8b4f583efe6d3c41b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf748d63ea8ab3a2346187f074c8931e3116719527eeeee02fee559ac48f2560c8224d8b6183907be54617bf0cd3b05f15c431f5c610a16e0131d14a0658147f7e9ec152374e5ad8231d0e67999c9ca05d48d8fdd31f05f9d6bc2ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40a64f479721b671429d15055a60b322ab67d72ddff6a1f4c28a16f4f0479a266698d968c6f08b8bcd22e878193fa232674196e847bc181e789cdfcbc9a4e53f79c22f653552be38302022a432ec2a1339676d1fe7d6a5c5db98d9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119314a090d3ce5153e2692824362233d4bac445318781f3ba4455450a21e7852f352c417d313e97553267ec043389edaef0235e08185cbdb1b80f25812727f3029e34b532d3630578d7c89ae15c362ff342b69dafbde3de4eca4a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12591a3d1c41336099b4529b4305d8a28dd37991662a18c80a8414fa3570445f3295c526ec49d262add97386a8c383fa8b58f92797037336e1f42c3688d84206efe5d726e9caf2b991ce10b78cd4b560a6ae29fca2ace6e47201b09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1552698cea0a23d8ba21a46a9e9e7441c80f5a15442ab941ad5922566ba3fef0c1c4f4dbce2796575b9f3e026607d58cabad36e1d3a53e2cba8dd3da7f82c500dcfc925ce9c3f8ec40d7c59c3fa8bbf756a5d62f953b2174c2b7a69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecff23ec41bc31685166e74e8c4d0974c3935de5e72110a0598a45eccb9a2508e774f82a6ab3a9a7cfe263d9f80245945fc2acc4cd46a6c1a07e339854c3cda8a477189529fad7f7b8884bb90a9ec58006aba2d1f79ec3dda36a52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131a3d06c3d4d535863654a797fb019ae1dc211e121d513be0d427bea97d77f4dda79b4a1d174cfef89d613ed285d3113490a58c36edf2b324132838bca31736665d5e59eebdc22afd5fecaa67b3bb7479714f4a28c5b8c92f9cda5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h818eacd3e8fa892104665afb6a1ed30e837cd48932dde261371dd802b8e7d79a20ff2385e217fa6e067e804429f50a06c69c79e552cf5247702196b46d2a77f1517856226a017f4b79f09a9baa688e076d6c4aec8c7ece1327b16b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce24cf67be700e8a0b7e8d177ace60fb380f9b92f94db597d52420230a7c2480a1b3e62e69b29419844fe64aa44e49f5c21de16c76c246eee6bf7fd8e374b04c705cd02865a45004b9edb8451c8a86a7a3f05acbc43e437b869e34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f557f7f2c6b26a29f2e24a1bdda155510c392c1e83af8f8c1e37ade8b26efe9aefa92cdacb3b6f135700205063995640b43079ce61e67ac509e9553f657fd8c18ad24bc1797b228eb45e4a043ccd5cbab102c967c8ac252f40b41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166aaa47fc9d765b97b950ae86db4e7439a8e7d670db9f51e5ccb67ded8ad684e5f6b4aa9ddd01b7112c1250c5565d0a13a936d23ca159eb53265ec95584532e6beba141aee7642d093d55651f7e1ed588b35dd2632811fc9512eda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8fe50bfa7e3d0d965be7ab495cd3d37c005b82c356108de2333dccd1f56763d02069ef193121ac076b48edc75e643c122f9ba2d213fb8b24f0deaf0e5c5654be37111ef6cf46e65630cfca452cca1aa702170fad66a50d1a437c6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bde2257b88ac25e22a5b069d736d42b1b9d746398f977c8f41151fda50872d9dff75b8c088eee1115237255e0ae4d46427909f79d72092e50f30242bb13a907b4111b3684fdec1061a418f87f9f14317eaea34c317d56a2b4f5f0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17460ce48d4562c4cd32da41b981a060e4d44583623ccb8ffecd1af042fa997e5351c0ba7ad7c901c9a8970e36b11a4bf2587c21c248b334ebe49b778411d49a340954fa5d3f994219bbab0c9d41dd7e632ed5e9e71b72892bda2f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h823ed35143588eacb12953cd4ee2fb208c158d90902562a9728cdebf46011b3c1da6fe32b37ea6cbf9d98a383a3182725d94bf1e61e19c94e9713347bbc63f7d4d59eca201db24deabfec25fb14452510be60a73f66f40bd45034;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ee961d7adc2ed7d87c77b57cc42df3d472e732350b3a3baddd5390f75631bc555df3857a7655687863a0fe3231c21317a805a3a0a62b69972f0dfbd39fd99d28457b6442a64d09eabd21e9344a20c2842f7364aa20cdd598a1f81;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1abbe425f78b5c405d3be59fd8649235c0199899b59897f9f27921a8d35dc458080315534f69616fc6d362df41369eda5b3925bf45fd2120a2cad2512ca204a3a21ae84ecb67c94f9c6c3756ab81e758df08c832e30ad9f07e97a97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7db35bc548fe558fca7904820e800709dfc928d0962fc0fa269f33103b99c3b5b310f0fedf598b2520216aa6c11ddde3476fd4904bd38081968aff5faa9df4dc52d605e3ae6397ff6192029314388b16e643283c50c6355b8c48d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c35893a0daba1beecad1d0ab892e8685cb00a24ac26e2a400f0ca025884b45871d4f8f30b9395fc24e2a53076b7442d02f5fcad074eb87726c7bc0f70371a9b15fb243bd4536827ad75baa1d67eaa15b8d5aa1b38591c44afbd8da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha72f1ce5d2ec14513bc70745999d9ea780680e35ca992336bce30d1ac3361dd833b6257f7cad0c31dd483551ffb718b83865038123712a4ecb6ba944e7cedcb91005f754464935f6ec57b888d9ce4b6826be099f7e9debbeaaf186;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16083c8dc4b9448a298123fee74b0a7fe8a436fcb2591517c68e3dc4c768adde4c5c8a29d62e2d7f3400bdd611a1a8be87c80ad7f08d262db754782dbccef1797d4fee0557fcb2fa64b2eecc18166d0fbc521b606b99e3e85934665;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb04840c1e9f17131ea2d48f1629273a594473778c728e0ca79886e1db3dc0f5d4f39a391603c59705788b3edb91b8e3b3a1b213da80736df2f40bd928ac537b513720311d641db7baa52135eeb8c26a0c801a7c7c28837bdb9788a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h161e4ae3fa5ce386354fb018a73de2ec45d74ada6812aa0accd24920447e66e55534c40e14e03b0452acf30ba9b8501cbbad2b06a11eda3aecc08a3c191f28d5fc05c22fc7b847a1bd4cbe7b43c4bb685f6a5f7547e8dc1cf98260d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17aeea8e5cf4140fb55986d6159f736a8ee9a56ad1eb9c7bfadc109b8150db5ee21f91cf9bcfd8e4409b86807566e35e8e0e41a9e706f296e8b9a6a225c353d8f9b6f1f1ffa649efae052784e2a45b1dc04addc11b1c7f9d07459a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1912d496d92e5c812653b9e557f698bb0839749ecb3fb1117756a80c57de92d77f7c6a36f7d513f524f78db916c865b5c9f0235915cdc2b563e1a279a9db7aa2614712eafbbb0c2888c0939cd79faa17051edfd8c085a44cf039ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46948985fa8fa98ab11fe24c1daba8ea4e5a54d06abcb8aabb8bc89b95554e6b74fcf1ddb6f6f911cd7ffdfc3181954580a56611abf53622f14aa785441ed3f4d96247fc04a18b991d5cd96dd30ceb398c9af588d55ffe46398fff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1641aeabb28faf8c2533f4b1b84fcea108bf647a2eb9f54c8bd792d6c61addbe34b49751d53789c5801c4ccc4155f1c6138a81f6351ff8512c74ceb6d0a7893b3e6ba3c316e90c9bbf5b91ff7fc3422cc5374ef1d133f6f707ead9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h556974bde84002f43186b3fa3847f2487699f98360977dda6c0b270b456a58cf5e75a59e83c62e5ee7d43dc600b05585f23bf2f42e8afd60a6380be49fbb5063263fa10fba417c83e26eb967a9d42470e483113c131aff7e575abe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h60e46edee59162dacde0964372d75527d16afdc8bdd8912f0f826a4bffe802b7ee2a6bb611453b61628e10ba44343bac015bf0b72ed73969847e85adf7c504355f485bb6eb97284b6764b437ec6e3bf47e3f99a4eae08e2b5c77af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf7325150c3ba4b439920b99ba71d0d9695a0b421d277f29060de924a0a20cfcfea2b400561e9e473a6924f3fa985bb23034902aee31fdce984e309472260e38ba4b52b3a3ef3af22bef0adb8d5c2b65611327eff73b1e8d1ba0eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0bacdbbb5e4f919c59558da0c772a486350fc97f5d7ee7a49ca601a2ea4a224f36548b346f4108341ba552b72ad3a920142e661ed2e14158e62414eaf55dec45aa802c8537d89847bd31d8caf7edbc143389a519544a54f3b1105;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62ac14a61e9ce3262b374d7a1ab7332e290649105245f12f0af34da45efd0fb067956d7fb407975f5d3b8cdba45e1c309bd3808e3edfee73ea512c3617902e598c0e0ca4140eeac1e1c6151c3272aaa2555ce9314b6e1dc569f255;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119cf8ce5d6b7bcd80697c21e1664d877529a3ebe49fdd7f18fb405525cd54335e952bd34ac98e5585b903cc0a89f89002138adbd0263f84a15b69657fc7d877cff3f2193653336e409393b461f30909da847ca108bdc26609bcc90;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b2d515725ef564b251d5a5c6074cb89f1db76a492bb5e5244ee0565b4e284a19ca53132092d58e1e886414bafe54a252d2c70fb8a1e18613d8eb502b1574ebc8d155995505f87d04c886aa2473d87059208a95ed976b6e200dcfc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ccea790784f52c17f6b23ab76d9eea108d667eafe3ce74c822cb8e95e81ba2a0f1b43a63a80453c5afe084cb7bb3ead0415bb2691a6ab8e305a09280327312c19d21c26fb131bf7e42a0600789429423158aacc9042a7adf126e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1eeac63786a6f32edb1011e4d2ab785a843f8439b2b9ea8aec273e5bc4827329270f79f78a0b23f694c932df6b90328a00abc0321bd64f12262fefd91e788602a6b4bb0a48d95f7417d0ec3bf4c0b30eac76872a6fbda30b54a70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h161ed60a4f16af25ff126b3df4d60a37fbb16b107d7743d60bfecadb7e13069037260f38db6fb5e7411378ad1a1c984aa1563eb7f2c1a7ab12c537fb922f9080c4685a900f79dc7ee83e9b38547a1458b18ee3b5578e7597d845f35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170ea3995e1f2def16e6b3525dce50274347aa1b76566fd0049a71c62b6c469615f8585178a396cd071220b221bbec03dafa07e5ffd79719bcb8e587acfcec8b3be1849489a33a1d51938599347982c213ef71a60bde45d5d738c9d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbc752f16ca133630a611919bbf924a6915a08ee9fc5211d7ccbd37a383707ef80a0944ecde7624d1db32ddaf41645a43d8d18f7a729da665ae886cc7579e37c6ba72f4cae9e97f3b5d18d4b9dc6b8fb7ab77561bd2fd2bfc612db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fcb01ae40e83b5d4c66657a448e5f8fb5c552134ddf19894a527d623fa46a75c3bf9f5d1734dbea8e1df186e6d31cb3960fce063ec0bb98ccfaf0582426077caa8b4e3835b0ef00dc8f4a5966ad2efe0c7b2886d2244ea7fe4d5e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h955c1f7bc61a3b836cb14b4259823603f3636ac3e75f9a2835169bbb07e1e7d30667051d9ca0f262bce9bc1e0e10287ec5174218fc2448e78bb1972c280011381746c0a8f0096c844d8198bc0501080fb1d549d8dabbbe89e99f00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h584510771272a04a56de75b7d6517b7c5de2441c1dff93c0f069497c7219c622a07995ab5c500e1461c4cea2c604bd459d921f3673b75236618fca239f01a9d82e6f335fc0eda0a95290a28acae9f237f31890a86eef5c12e69649;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58fdc877a020dd507aba343c863668d6aacdf9bbcf5e692c7f9a94e034b5caaeae6aab20384d34140edeec1368d848d67aa26316d5982d1c65e02f0317155d16dfa2dcdb1554dedbe7754be00e512f488fd09b70262895b3e1cae1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5769f2c43380479381a2575a9c18a42b62544d5e080e04b1e5db3cefaa93468fbf729f3eee3711b7c89a8ab75354034761286f9dd3be2c27a3b0690369d30a4d5b47a18a59de6859039fa9ced0eb728386a806288706567da1ceab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6070d3bcad47946408b0e6c6a35d6e41736401189f8bd9344e5982c5ed2682f1332b07471a61be1d62878799f7c66511940f9841c15ad503023ff23f6d77a9b4cc4e315367b03e671cadcc94101e42d02a514f4f3ca013aaefcf3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4358d06fa8a7f7237604bc8b283442b7e4e06245eeb554184cc4cbf22e7ed6931ae3c148bc76372c38486f1a29ca967fc8c5711dd5af78b68a95b6210f5d383dd3ada6d1853920164d9ab0b7a2578b0944879050db39295298f220;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6c247e38c15baf1408b1e94cccf29b6740978d27a957048847b3d2fc9dbc1811933731a97b123f6f905cf0ef532dce19d1dd18078acb1dd1d7526f043ff9d3d34d11f63d0c0e323ed3dbad918f9083a624249f289eef2191c8666;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79caddc9aac777f1e7814597cc7e4876f965c46cfda3747da2d12c37424ee102c9a9f40bddbad3793c2e2573b6b295b1176cf9154a92150b611c6c465c45fa818ca4713ebb90c54c38cf3115150755523e25df02885c7e839b9fd3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6ad6948d6c7f9a9ac295c45c7b05df6c2742424f0e2bca251f05cfe80cd35269efbec8b1497fab3028166bb3582262d326438627f2d3d04ab8ad190a8197c993be3d259d96ca313205f790abe303b19559f4b7e515fdc6abcdc01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90f388de77cbd2041a363f502020a5ba18b3433990cb98888463cdf3210c4a69e4486d86a82a40de3e5c3a251173becbd9a06d9055e0e5812ea4d04fbd16538acff5561a14f248c5cee41e85f3f4bc9405c6ef7615b0516650fa47;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5996c5bcced9f7f9294a0d0c184def8eed9a662d198879f44c834d0152e4c4b9234392af659a1dcb8d5203f21cf7e3a9c4e7b213bb945e755e05bdc4910c065dbf65fbc0feeebf42bd5e64d198a50cb534754fbd8253e3a18135b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c52c2efc9f5f3e12c3cbc9db6a09fa023c7bee28a3d1d763b1f31b49b33457a6a26aafa8f4c84ac11ae6cb2c76ebd20973a750734b4023d06fb1cfda0158fb949d6cfc68bc63b356b515c990e1f7f558c534bfacb31b4a337e62e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fb0110ea7695903a8209ae70f401aed924d6fb09a7ba7b42e645cb7449738b9e43b97250e5c618e52cce00a5f0a9e8e278daea6a8a40bc71b0b01f8d39b76aefbc27df09581be7c0ecb56a7ebfa0b53f6961b098d7c1fbe21e970;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1148c533dcfb35cce912771e5f09015a0be13d600d5c240b5b48034af097543cf79d56666ea257d5e36626f81e174c950a46e7eec636b79ef22ddcb45a1b167d784e035596aafe002c85b2ff62052b49501717eb1e238fd8e0daabe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5cf4b4288dec95fd25bc22b3d19cfdca0051e5b826b3470595565c174572e08eaba59f6b92a529ee42a80f9cb6096c4c472bc20be643299d60879700f5f3c345ad2c696303943d4d1f481e5b39f7a37ee342a400e633c2461d9fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8bdb18ff730277c74782bdaf11db995de289854b2af2c56c3fe88a3936e57c5eb1d995db2e71f897320ca2dd242761e5b6377235bfcf540d5b2cc76b085413a5b2f87c0f79b91c865b7237edb908df95f360c44a052a2d0aa3c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f59c134c9c6d73c79bea96c4fc8f86276cb29b4d7038fbeb00d2084b90cdcf919696d3af7ffa146fa57c0a3ee91df70793a075dd239834f078c2858af574ab61fc7f8681613a56fcb6d36c48038f164a9d0a3c7f6aa549e4e0f89;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3fda80d327a7d49576f3127c4f1ee4163d436a2e3c0de919493ea26ab3cf07491c70166fde7cad0ee3509e455390f9c782ab43d7696d5fa3fa55be02b25b20eb552ff260c54d98c74d22f13173ffc0202c5859a6a6381289fb0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h159c4e6c344a1902c1660749ee7b9b2539f2ab1b65a1d5e3e17d3493841a4368a2e01afb56d31b84c5daa7c2c22d87201cec3455bee7cefd516c654185b51b47f9dfda8155862f2342792de842166d49e3cc913d2778bc164676c8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2cd3ae2d6c01e7b57a11f96713ec1c8113f5e32746b2280f8a611213bf57f241d9059caf59656ff3ef1dcabac52e976b093ec3a67e68cc85de8f74906447d7fd45d2fb4d504f551db86237812098cf243d6bd87392020644a687d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd547346d3ab2107f6ce856990c8217f9fee04f91ded8f337a2724a04e94f931c44e19c381ad4a688a047f0191fa05f5e443f072ebb7559d2b48cb884b983c383ccf2c0040d88745cb2a31f2c48c1f9d9e606749105666d8ec2ca9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e824a2b0adf52579b548e98100429818a42f8005bc58c7865b4ed76e54b3e000f8fa3c4ab2d638e7bc157f3afb256b5596fc4d614a1335f9a5570b5641ba1b9682291f2ca7c03732aac9aac6abbaaaed6e1c5b6452eb5fea33dae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec7485b7cc3c6faae961384f2e9ef0df87bbf8b903983d02a034d2981b4462fc6b60c468a2688c7d1f9d086b6452ec47e6a2f8fdbdce0f5092f1b2d3218b5e7793531ec962edb91c1018a4c40aba63499df36c142eaaba3794bffd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128f86409cdc15ec84c4d892941ae038beeb91623a7e21b72e9a64928cab9fdca8711c43ab2f8595f18e2605e7d4ef05ab0c7cf3776f5b05d006e27ea42a558491510a6b7bf103e347d1bd6511a076407eac2712eec3ef50a3ddf7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b591e954e2d465a8938688787c66619c3f2538a982e0404fed63708265ee8aaf3d6478199b7cfcaf15b52c44c9c901c58e65895e6c83753c3e2978f25962260b43421adf8b1cf5cea1987f7da71e1d0ca44db5af48600dc7531c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149dc6ddd1f617b5bcadda7129d6cde0f81a7982c3a648a3bb8bf2f2c3bbfec6c14eb08b8f3c3be931277dbbfe2dbe7ef21da4131f1ea4d3b4f245c81642343be4adea889b4a84a9b088aa076665aa3ad9ba21bfc92634f417c87c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h896e71b200fe907c0c498399521474fcfd1a71213f600e06ddc3f8b23ab3568a5198911deb320e06ccad3ff9e8552ad0370272fc817d98ca19abfb903f10d27fad60ac4705e31397d00357e864cdf4e41dca6c05fc30d331363c7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf37620a9868dd330d48632bdb8c87b072ecf00f078b31c5280cc69d2deeeaf957cca4823a65ab494c8e3bca152bfe808ce2c7dc0a4bcef1f7182be76ed363c7cd11b58155e79e1b17df4ab94d5b563a11190e3158113cf3a42a5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7dc0ce1c9524c0cc96e213d8e4ae89a498ca7327a85e34c37510aee96271b33cd68823a4bc80a554989b3c5340d9712e2942cb903cd19b192b83d15db931f7c2c569b6e7cf7b668c65250fe6b21a53658518fb5977925a4b559186;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda2e584f0e56aa8f2c169d967f2f1c4f1f539aa837068cfe1814ee7824eac6195fef816376aedde25c5592778fb1ee248641b6939943f5d97c12de5ab6579d9dc447d95628a61794c439af4a1644b40c5bf871890f43d613209f01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c26d0dd05160dd83bc06ceb4ca3a816a8369678ba3fc47bbdf9876fb0fde4d8831976ec44c1e07703814730da43c94f0eaec3810bd09293aeb54ab7a10a702ba35ae4b1d45d1a22c8a11e3a7fde5c949c79b1a542a7f2791e4cf3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36bbd0d0818bcba9b70f1e3bc0a1a4b089d056718b0c5b19a990f019e74b88d6eeb628102878c5a8fe0a65b8de9973fe3240a54144609c378372688a3c966c43049c096863fa7b4e708e0d03dad68621249990a6873ca6174e7e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9631648217cbcbbb06409fa2125c418439329bd618a012daef43bf9a1759639b3a0bef419fcdfa8830d05e52dc7b90740c5727cf324eb233ca226de901338a2acfd1c626246907c2a435ddfda77bf2f2ce0ccee1ea5a17dbb81a6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1158dabd4cf9c937b8c9ad4af609c54aea5970f6b86b43c01ae0c477d95ce84a2c35b9a7742e1f37bf524ce8a5773f1ab83d311f2101c9aa2d10d726b15cb9f991d369d3467245a7c410d8293ee887bb0d8c2ad98a3974f35d2b661;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd58c6780ac06942b69f20b358bb330aea65f1d1ad07896304833ed7b1fb8c27a4bdae9c35ec7a836a0a2c190e3d4dc85d9f1b6c7c577ddd3cabc8a8650d1ae0e0e55871755fdfb2fdb14295c56e6044a5d6d152f0e1c42ca0365ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135978437789a72bbee877032a28e7c9f110035c0af6e7b9109b21f90c7d216f65b39d2f097075e37fbd236956daabdd45f0de4a3c40e3dc7f5e5ff12258e397a31898c1811aa5517906770e1ada6b6223224ef843ddf8d37e106ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc27e3241871c619bdb7fb34aa62825df07d5fd9b5749cf0fe149a393b766f044c16bab5c190ab1c17549a65ce74097700a76addf698670633e940b8b08944ccc8f5e9c40ccd52f4c315f5389bca784decbfbbdcc3c461726901b34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf377f88bcb596cf08d8c0fa49677f96bb69f30941335f6b546ba11f6ed3650a22a89cff9fbe6a576ce4c8ed7fb6929a2e23abdd25bf8efcd69201d97cb547d591c5f8aa36fa6a64dfded733bd60c04879d6ed91f8698f84cd5675;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4b1e79d685999db63bf69bb0cd0eb9e6bd3e1dabb14ae0783355532fb85325e33e18bd67a66f37be8282a582b86440a7af4a01665c4167a946c4d17362fdf2b8c5f28331519a7b8ef7bdca792d7d9bda904a3a54a615b30fa1d8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2029cf546a2accce7aa6fb8d503417d13be4481d693fabdd414f67581e2ce29553d8e53ba470de31d59a23617a1f7e10e50e7b39c86904619a1b6292a9f680469bafc87a9be7817676d7dff9e39c8768c1aaf0960a19c77494551;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h169b38d2c071716d63e33cb951ab1bb191076e3ca073c0057cd1877eb92958e1f34bd52cc9612394011f26da63b0de404050e6b31af646bb73a4709c3606023f8ec45d1012e8b9179f3ff677e6ee11d4a57142e6e03d27ca64c7e9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155e70076041a7f5225fdae4599eaad5c32350f38a406c5922ddb147537eef0849f3d880574b64ea65b3c4253442e5ed01bb5e140eaf8a92aad8f862f2648a81dd26db44365405b10ff4902efa3607876d42116adb70bd507553141;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41771937b6ee829b59e53a667619dc35ec4fe85a4a4abe8eba9761e0760a796a3266a10c1a809a04cc7b25c7b695cd992b73d989de8ea6088371699fea2d13f482143315e244bcb9e3898c236d81c03f5ad6bdf0e8436e06b53c95;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3ea30436d9abb612853acd36a2722ddbc466e3d051249bfcf263b0fc52efa647502cd59a2655e6040ba4f92799b61e28c24a9f43b898bbdcdc6747397a9ce2be155634a952e5d7550e63f701cbf1381c748dfe7d8016c9e9dd44a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3b22695ad888e16cd564cd7f0ea54bf6bbf1fcc7545fb24a603b7252149f16cca293d7623dc29a2c845fcdd1d9242d46e0ef1c8ed8fae0e7736c6fba7153f2e1430f27dec7bbc28826d6d7142a1e478d8ee46e6b58d14082441d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a46c760cd5cb0489e5276e770af3616d86c95b1528f1cea815076ff76ffde5ce06874559310c69dae56bd5c7bf0d6beb2befaacc1892dae195b02116bf82d2bd85bd2cfc2001dfa917315392ce92bbadcb8b797ac571bb7cfd6333;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17505237d17b15d60febef26d5e53b061e9afd9bcd65a75a00bab9d392c1fd418da127df55f4aec9a28422967a2ba56f6c91c3ede6af77624738470f8a67034f64fbd0c0d42447fcb4969e21308c5b0c6936b6dbd40c97649aa4017;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3435b5153d86fa02d69886d212b297496972b054c234fc1c3002e28c4de742c4ad062b0e5c021ed83233e9562eec32e724985e826c6b1912932ccedfa1b89f11247b7621a8c0af164b12c1faade2760f9d5dc4ade0cb3aeacf43a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fbc3c7e3a0cf3b0eda0e4467f584186574b818388b1dfda977abbff6d8f04781c40bc53ed44466e97e7ad2918f7770981eeb8071323cb9e4c6b1529f2ffb347e18001dcb0143a4e823b851e1e4d96773c487f349ed2e17c35fc9e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf9f0fbaf68fd2eaea9e9d9d1f16aa8031a533a17c5c41f2653215be7c7941e53606a07879f6bbd3e5a5dfcd09056f6f4a53a1472c9c307c92371a79ffdd9b611819a9f135be462e656b757c1b4058ebf8a8f02ede5f5f3dc467d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41521303b3cdd92a04bde74c38e7d4fbd871b6d45fbf4b664c63d3066e37e3b5b9b326dae4e8515402675b795a9b0361d04b80e176990f9f7cf2c0310ca5c6c92c7d889b8e52132eef6926f7faaccf95a29b0675b5c07ad2d88871;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdff2508aa893862f71d84eadf003b90bff4a5876db7aa3969a2589280a4ab14c5f868df1394df94a7fea3fe2cc1d650f7d2f62942a3ee1a66a65916118e804a9690235f6ec80498f1fffd6333a6e4bd1691d301573165c22c6ff79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9952962bbcd10388d41327d5ac881b2ec2476a17f35d7a26e3113e9433cdbff07c03574acf92f8f932deb8ef75930d9a3cc15df9400bc057757e7f3b8b56544b98856b0f91f011d5f4f135210243a9d531d87f1b11d08cd72a4a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48427474a6b245901889e077ee976a6219e6368991b99bc5638cff7c58c096c8f30c1d131ebe2c7f1bc1ff5090ae1dd21c2975add0d2de24e1529fd73346b87f33773908429f1cb2a2568b6a94f8a8917dfa94861ed9a28e86e8d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h580903f570fc893d9302354459ff05a86ac0d231cf7d2ff0851a9a4d3667f56d4d57c65a1e421b94159dd2a1575590752fe943d0b2b83e189e404359120fd5bf400cd162c5458bf22f3e533a7365d923f68d2396372b0b05fbf516;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h31778471b4b4863b993fa8ec2a845ef1b470c670913a3d6708001c49629a3b8df692b2e27ed62f1caa593576ab8bf6e5fa84dcd81b7f87c287326617cc19e4849ca49c48236619a4c02d20dfa4a4491fa2e4dd3856dd532033225b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be17795ddfeaf9e2736cf5e3b1fde6465e760f0405eaf093e8022b25da81d35c4b4ec6f55e835bdff954da9a489b60e58e813893a7dc05fd05f7db3c1fabac85add42f91f3d94e17b5807f3fd0b0ee2cade9199ce09ce74a6e5e9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf26717e495e5d38e7f68a542f765ea3b2822f6dc518caa6f025dd352d57444b353bc29bc05807b286e098e1866a40b219ab131731748dcccf249da717a731f0031622daed71e4b5a99c29c5251141f52d28c8e7fb9e94e8be95d6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81397f1f4d57d5e8c62a7957c0306116e2f387ae3fe512253b8e09addfa538cf58253f1f068cd6c0535473a4769c6fb8c1bbed0cfe84455e5bf86737c4b7a296a126897194258405f0b0e917de3708b8d7ed84667ffc0cdf62af2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9288938e6fe80dfb642b8e4d131b1b3ebba7ecd113f4490b415e823f38069a169f8c5bbff99efb57337537fdf9c6c79624beef1be3fedfc5d6618cd3c842207a906a111d7945fde19d51e6d6f7b20fc651035af8421a9796622d08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179263c55045dbcb2095e6430cf39030ac1f46ddbc2382026c49f2463aac79c8563e31ca47189a09c0d998559e0226f0e406565e67c202963a5d04cb9ae75bae3e60eaea3c790c21b759fbf55bb3c08f4622bb3fa6553cbf27c4a4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3c107b56a4a04135e7f1c1c9fbedad4494115a67aedb4227850bcd3252ceac55e0d2e61ee0ce580eb96850667babf4419691d4fb9ad8a40127bd06b121bd7dd69d336a89f69c921730a0a85db87ff7904c8646494dc02082d9b63;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86d1c1b7aeae720ed6edefc6fa3ed8d200d5be9db2ee5bee15994a7628a8382d2b53b1f0e1635a3b13e7dac063aa01f27d548a4391578dd0bc3bd95565fc770103a03c0535a2c0391d309bcba8f451655760aa5da4b05b58474fb9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbef98bb8c82d429edcf0814faf3298098f5aaa38a9f0404c3e2aebd2512b2bfc8db5dc83ef178b9a4c47aa1d9d31b801ab8878ec2c4e52258e6b82bd8f81d3a99e9b922ea2cf6611e59e537b00b8ef3396aeae52129e3d75a198;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2f2c540cc4c09dbf4e1e4b3716c8f30adb84505450a45d06a9a51122c3244af76a7c4ea86ec4792e1727409dc8a093564db682338dd26f8bb160a9a8c3d5d8a4fa6f51c83bef063267ebd138df33f5d7508ddb404b805317b20fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1708edb112ed3fc8bf36565ac242638d41abf7b672a0a05866c1e36da7c74329106cf8863f18b6758de1dbd16b6a213eabf8be6173421c4d2d75e00f767ae4302427803488a2bc08126abdca7c2077e90a550e088699365af8dc6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f96c8b216528b7269dd6e40f2cdf2d824bb33e074a643d1fe254f7892f050232a2851974b4ed3a48629adf5ad4a0362029409ea8b4ba0e1a1fbf2c7e03d109461ff0b3327862e58b5e446a1eec40a0c1e816d517c982db6d41efd5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c15aa543fb0da264983aebaca02f09c68f9b64027c2b7203406da5ad8516af2186e7149d556d6552edb63c807c4ca123a38054a8f0fed19c81a17f3753f4e7b9a4942b542d6cc8b91da12fe3f98df9f72dec4782108e29fd228e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f458ccd9b96af6430c9c4037661b3517ba9b855666b67998c459013bb0824632776ec13e6b4e37c27104b4ac7d2c3ec0d2e7c0c587f7125b24098c894378b6eb1350af311a4594bd7d4ec15481e919d24cf04b5780a257d516f16e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6aee517fbd7427a4dd73942be283c01305c61d26bbf0cd712058cac5258ffc7123bab2b6332b8fe7cc358fe200e8d8a715681728833d728dfca1cad0553b6a83e5fd1aa97d789a34cc658f632cec741a0da4e3c04ba54d8d6860f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha45b7853641028c13d51583c3b6d35337c69ad9b9e4fcbde3e7e394d423acd59c6a0896a2c2859957e2680124758db1ffc392794ef56048d2b18bfe8a996274136a76d3f407c28b621cf24f82476b49254ce941315770dfbc02ac6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127cb00cafc8cf6a2dc8233efc661bff0f2a3e7254c9015eb24315154bdb15a7f5ffe2615e4a25d7d5d8841db3328353e841c55dff76f7482cb08767a782a1e8a4977472707b8ec61a2b1ef15f1ea1f4a699d289e7e50f208f8a2ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1954195086a453305337957c7560202cd9d62ddee24bf9a6803bfc1994f484d26cf3e424b8701a5342589d858c1c5b74a9ac526cfdc1eefadcce516f4eaaf1f120cd9d7f3e86966846439be17fd0d59dcc84ae0d7f4d7796c145a22;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0c4d82cf1915e1f9872bc41eaec244268abf3a2cb6060019f78dea9e308c1819a80edc343cf21b66cf1e6be243ef86009a236a521235909ffffa591b65d8839bb20a9556d3e32f93514443505c16eba3df183e7f5d596f84b1f92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2b3c35d6cf3766f8a381c11a21133c9ac14d94def1b93558df29a02155668ab25bf84e435d667722f0576433415580243fc0aa72b4f1659b5bd4fee1e5086b447594a9da5bd580dae7eb928a0bacf8a0a2a39e578e302bc95c3c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d8084f467d59cb127e93c37f6ec301078030b9691313233d68c9dd427c981cfa11f5b058ca882afe62dc960dba41be4f8710c24f82159033cc94a18a9f6a332fc1f2e5fe074219e7e126085ef9e4e66b79d98ff64b392e6084db0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1669ab385d1c675b49fc0d7f4700183d81b6b86cfd91042709bd4c30b6dc66a6771eb53234c9bcf8683c8d53781a7052e2316429225e8b41fd7811fb8b8599de7a6f20393445ea3b2b96dc7264c41e8e90252a189a83a80250bbc6d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h56d047d837e104fa0884f5d723e0cbfedebcec07d3d81d366c19f92335433700766ee88013d99a82f35b23a1ccbe3b0b0d6f865890b22b4b770342d9094cccb2eec3a943f87dd172ca37150efa8486c0a94be90138b5708b11dfb0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h762a743765c4a53017c87ce52ed38049546b14748742e1251131c72b3c3100c3b95ab169d72d09f01c99e3d4dcbcb286083f687b9856c3641cc6966c7c1efbe3d47d5597ebff0395e4fa710d57138a54b290b291f3f004280557b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a0c43b535a31052bacd03fb36750bfa8021e9a920d3e7dc415fc6060351036f235672eabb045f050d85978fc0af3e76fe274d289046d0b524821a9395a8bf072195c107d9c7975542d4264f70f74b8ea7a7b66b33614234758533;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1714ec851bae8b37736798a3c9decd50b5120078dbe1d5d04426288ea9c6987d6b13180d1df08ba12305cf8f54bfaef3463dea9a47212bea6042bd591a615c001f001c4c6266d2fc5ebcbd02bf1011d0968fb09f7aff1233ee52b71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha08b8673f9a329019cad6f19c1a77615ca23d0c3aa98310beb8094a3cb56f260e4a14fcc43148d5948cc8c19faa3573b51ea73650fe691b74edca5fc3a0dcf8572682981bfc05910a726305e1aa973ae1fc4351905cf06ac3b3852;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1165fcbd3318bc443f8c45e1efec9fd064f3fde5fee7f15bc950bb34281b6dc72c7ba24f32a662e54f491efa0758069d25ed7f45065d6ed163fd5e61a8da2086f2dd93a831be12151985881fbe763894394b9e24fee3a370245c5ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130a1502cecb89e19cbcd7d65327d28a74e61622b39ef2999bda39afbd9f0037276523c13ee3b0d82071f7fad5909c2b6fc7d5964b86948917107185e736d8288e7b2b8a691950dc16adcd2f9d04bad7f624826de3fc75658af95b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2e04606d334759a7015b64000cad01ddd6b91375cdc4513a4be2dcc68025f02a435309a987f6cf6ce6487b2abcd9d983c8ce8ca3c6d12d48f1aa051f6d5697b407172a270f8d223d205e17c6a002afb9293e3b9da7c0c780767d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c68f607eb4719f47897e7be35d7f1059de92960ff6e8bde11b130b4cc1226c15b66273401e45f30c4e052d49c7e4d11bee7035f31f590f8792ac322e95b3b24a640487aac3dd7e17c26ceb481d3cef6e70073b239cb355b5514e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed74b439b13c2f0fea085421f31f15fcb8a882ada9bd33cbbfbe27ccd6cc5035442c70b9b7b5780a2082edb8d95c1e0d78df36e968979d41e3a824b0a5e9377fc4ed9e91b118aeb59ee6df9fd45a75c65cb7bf203d1464713b1391;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190be517f9c1576f4ffd406c7762675fcc91ab346c4217ffcb0f6419b7996fbbbdd798c2488e875e9d89141ca3355376fadc77f7970df84d7d3346d07fbccb0dc722966f41ef8d68141fdf1f12e211b209229a9e2990984552fdbfb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12711fd4910489d8cf69cfa58ef480ccd78d7590273269b12503f3180a6caedb138ec5a7abaf0152f18f0ec3f843a74f14a7af4083c1664c83e00261cc313ae13c65865044addb10557a17ea74f1d16e5cb07090c9e3891a74beb0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3a0dd59e0b85618404af27a396f7339a92e812d790321ac9a40c361e0f750aa89180e3396498cfd4f477a32f0fffc2c2ed7c3c954c8e1ba70922a7325bcea1d829dc9b4eb21d59ef64a7aa8b575663ed76671015e38834cd302c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd38fc7b1eadafc0f60ad9e211c6705448120c74b7f628bd5780ab4a4d9a823bad3514342c4473735676043f23191cf22fbf988069cfb7049764136a9f782223e8e383859c82bdf4e1fb9d433b326a4c96be7d48cef8c2a862a06c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1337c97b9eb792de362a3442051db6bf5ae41620012aa407193465b25247658c4dc1e1e9bc999b4d11e32f76e632353b4178a0ee9c918b4f06997fd8f5f780c67f469e464567e7036ed3ea9c29a7c712ed2ed29cb71e41a60097b09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h941a105d06c115570f71e06ec38a5b7a95383c09223ff5454894bff1bc90b9fc279e8faa0bf8050c872ec5c7b240cd025a6bb2dad39a91b953e7d589f5b5348b46f10fd934e5c3b72cf33a9f1e39df30a5f556a3024a37c60c76d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c981e52866921a87a371c86d16ce9eb3ae5bc5637405dd1c1df6e56cb0408a0320b0ae645d84b5d01e3a979d31bd7ddff3e1908eaadaa75ffa0f1b4ffa184cf0ce3fccd2937efdaa0fad3ed6a4eb2861d681606fc70dc7cbe09dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee84ae816fb2d72614515fbb6f47ffd769cea2971f3481e70157b9379a3fc60703fc32a0352d339db788a2ea9ace384601b6749fda43cc679038143dd903db7ac48463896be642143e36098a6f80636450f817aa7563898674105e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd46ef268f1cf52e2f37f44854fc54424b254703075563e820ea344790799fe534e5e0f586ae6469e36c1835e3fe2b74e9a741c010ec21d6e1f04b5d43096832e1c484230c519cc2e65e211927c6ff7592147f71b5c32f5c21d1f4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5b628fce9ea1d6bc0f9e438a92cefa440975637878ae5e6422372e7fee6ba00faeb9e6da14de1e37e77d0af96d16e16223d5dadda5bc8bb9f37d2a628c93a9f92d7fcb9e832a784145eb569faa5c82d15c6a204b59ede66334d59;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a3034e2fc62ee39af308160c6f35da7e93b08ef3919a0146c1f023144a958d85a101edb27254a9b955ed34a829d0089cc1c38699a52727e9fd55ff6888410e3974f5f67377811fa290483952326b74447636aad2cb93fe7bfa516;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16272f68f6cb305019bc474b9b7dd6fd5efe92d84ea03d2369d3aa639af95bc3ce468871144a96878564707105fa4ccfe5e3bce6862948e9882347a60269c3b67756f1467114a067d82586ac40292f79c60bd636df8461c103615ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be574b86eb13b3373f27ae588efd996de3fa44280b2f06eaf47624c76d424efcbf3ed5c2e99ac76392b8af885208308ee4af8416583857a1a0c060b92854e66fd6de53903814931148bd8822c723b576d7496941e5b7895cad79f2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91a6d778179a557461478929f239e9eb3621930b79351e792a7bbde952b6cb12ca9b251e0e18407cd5796ae3c666b309c8cb6f1db66172c0a972626698b5d491c2feb0659e5b86b9704166bcc1a83256758be704843fe302e67756;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71aabc5cc76a52ad5e2a7a717a3e994e5a03e73dd0ccbd64ad5313a433cf72d497b682389dbc4642c8c104ae76e68e1bcc4b9747b922a0491a6abbda4ad6c99200bb1494480134fb981c682f5057b2d6fec039996ee573a35b2b86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha00ee858d43a83aff31a9f18d609407f227b201e4b8cf39add3743ef0d687122a9b5d70ae2089cff147bd114f4ffec9463e908b79025249111902d99ab2f7f22936542acc78148b048bee2e5881545f786fe9fddb1f649abfde6ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96e0383bedcc808e0512426429b58a6f4211d7daad2477df626411afde3487603a53064cd3612f2419fa1e680f1e1435c921744e5d07e0114e0ab237a840d75a267dd3e6f458974a35296ede523544f1d81c003ba7700bd389350;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hac41fc6ba66be5937e77062cfe085a5d0d39396f66e49b1a92d8216e5d7e644336e3d924b25e22841cbcf71a4a5411f718da5e1a1df825c8ad634de3cdf90a2ba2c5d7a39e0574f145d0d2de35bdc15376a81f237634017c8d74d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee816c5ca5cc550f52fc8e5de1b2ed4b8a9910a9f53f88ec64b5bc343f638e63b97cf7ef238bb8dcf01acdb88daacaae1927692fe7862ae88e805a1c7a149469d840940eb834c3e87f5018d3510d51666329f6d17d2a8165f4a8a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13fac6058953cbd8d36a0bc2215bf6e8b34b0dd1eb6cfc56bcde6eff6f78c59b234c9b3274fecabecbdfe38e744dfb969b06b2079e7b1116508e865eb2618ab9eb5e4e537520c037d6ce281e7bd98f35ba6e0f2b3683e16b657a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca07f93086365a0a718f1b7a7b954d45295d624671a6dd1e92c56f679a952bd23a1b979968003e4cc92bf6a57f776e0d764672eff852522ffc532875e114aa35d396ce0401a31a3ed5b6a7d1940ea1a75b8174dd7c384775c5c6b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40d693da100d7fa8b70f866e501b80a6ae0e503a646e53442f213ae8d39788683ef23559ae642cbd2c7188ec7294beebc3dbd69aac3f1cf61aaa3f03307a64b6ced231bbd7a955ffc9a6d06dc4cf312221fa65514ca887e38d5cdb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c9f62defb5b66ede7b72857b49f98541fcdf9f5467b39dc9b71cc3a11f7f793b788d8c77b6af654b73f8340ba3e375c236d2ff4825efbe6efb76e29eb7789e690335e05c6ed4211478a9b4962742479a89127a2bd5094e732c8bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14845bd7ccecb8357fd0951c1343e29f9c35a9169508af35ba3f0995c1d0f9f6934eb856ea9f5abbfa70b78c220096c7c3331772f02183d0ea7d619c77d3c10542e2c8134a53b47adced163ec25e8464420089ab6332db63bf662f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15920f450226d772b71550d11d81e6adc1b8c61d8f8d94ea009ba017effd4f51618f15da2e3d83d489d692825113d303cb656c2b7dbc291122647a202c2075d5bdd847a777fa39359cfc62f5d525292852722c3fc6b5ace947bd3fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167080ff72988bf9233d0d26a2f9fbec80f4556bca00ffe43f7ceb5f773deaf9671c8f57d8b1a8632986a0a5c799f37df138f0b7e3f0c8b1035f054820681bc097f5f55d14aa17385b6397c378882d22807e83c4e1082fe9146ee84;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e6e0dd022a8ee2e50dc7f235001ac3fe6bf5fa6f2621299ba2584d88d64db5c36a61048a88752c51472960392623e0cf1d189da1924336551f355207b41ec311640375c95bea022daf20cebb26ff76cb58f37be0f0260933800ab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1249d26d78700f6c146d90fe60c121a5e268f5e25e4ebd0fb3c7abf3805dc2c082b827cf538d0b0a49effb26a4b54da846bf19d82e37a941f7949e17b23a09498cedaf9e7f064ad8b399fc4059e5e38d750269cf2763ec2e67c7119;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e5bc12276a54cd883f3285e78f550277ffaf2869c4145be79db80d450f21fe3092b0a59c64873138a93e340ba8bffdbb9ff7ab1e61c6e2664fd4deaff7474baeb8294c5015a2e49330947b2632ee10a87ef6cbb373f205a56ed8a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e38290e46543cce2f37d349f278305baa8b788c192ac25e6d7103e86edf55719d9671486ff0e7d779e069c55458d04b45c410279f5d5193210edee61695e48a4ba3f8d9970975aaad56b7984f6775c56021fb3ff1a1d9afd5c4a13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f4a9eea8a43fc1029911756e4ea1ef8668cd664c3fbac832ccf8ab5ed35abb29c8496058f59aabbf25839b7032a84a15220392d63efe09cd357d3812eb043a3a96a2f03d9ba8ce6dffbe96ea45533ad529ba9d1f3ef5e82df26da;
        #1
        $finish();
    end
endmodule
