module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    compressor_CLA512_32 compressor_CLA512_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
        src16 <= 512'h0;
        src17 <= 512'h0;
        src18 <= 512'h0;
        src19 <= 512'h0;
        src20 <= 512'h0;
        src21 <= 512'h0;
        src22 <= 512'h0;
        src23 <= 512'h0;
        src24 <= 512'h0;
        src25 <= 512'h0;
        src26 <= 512'h0;
        src27 <= 512'h0;
        src28 <= 512'h0;
        src29 <= 512'h0;
        src30 <= 512'h0;
        src31 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA512_32(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    input [511:0]src16,
    input [511:0]src17,
    input [511:0]src18,
    input [511:0]src19,
    input [511:0]src20,
    input [511:0]src21,
    input [511:0]src22,
    input [511:0]src23,
    input [511:0]src24,
    input [511:0]src25,
    input [511:0]src26,
    input [511:0]src27,
    input [511:0]src28,
    input [511:0]src29,
    input [511:0]src30,
    input [511:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [0:0] comp_out40;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      input wire [511:0] src16,
      input wire [511:0] src17,
      input wire [511:0] src18,
      input wire [511:0] src19,
      input wire [511:0] src20,
      input wire [511:0] src21,
      input wire [511:0] src22,
      input wire [511:0] src23,
      input wire [511:0] src24,
      input wire [511:0] src25,
      input wire [511:0] src26,
      input wire [511:0] src27,
      input wire [511:0] src28,
      input wire [511:0] src29,
      input wire [511:0] src30,
      input wire [511:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [0:0] dst40);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [511:0] stage0_16;
   wire [511:0] stage0_17;
   wire [511:0] stage0_18;
   wire [511:0] stage0_19;
   wire [511:0] stage0_20;
   wire [511:0] stage0_21;
   wire [511:0] stage0_22;
   wire [511:0] stage0_23;
   wire [511:0] stage0_24;
   wire [511:0] stage0_25;
   wire [511:0] stage0_26;
   wire [511:0] stage0_27;
   wire [511:0] stage0_28;
   wire [511:0] stage0_29;
   wire [511:0] stage0_30;
   wire [511:0] stage0_31;
   wire [110:0] stage1_0;
   wire [198:0] stage1_1;
   wire [187:0] stage1_2;
   wire [276:0] stage1_3;
   wire [244:0] stage1_4;
   wire [205:0] stage1_5;
   wire [242:0] stage1_6;
   wire [185:0] stage1_7;
   wire [348:0] stage1_8;
   wire [211:0] stage1_9;
   wire [181:0] stage1_10;
   wire [205:0] stage1_11;
   wire [221:0] stage1_12;
   wire [231:0] stage1_13;
   wire [231:0] stage1_14;
   wire [236:0] stage1_15;
   wire [213:0] stage1_16;
   wire [223:0] stage1_17;
   wire [202:0] stage1_18;
   wire [262:0] stage1_19;
   wire [213:0] stage1_20;
   wire [269:0] stage1_21;
   wire [273:0] stage1_22;
   wire [165:0] stage1_23;
   wire [220:0] stage1_24;
   wire [273:0] stage1_25;
   wire [190:0] stage1_26;
   wire [199:0] stage1_27;
   wire [247:0] stage1_28;
   wire [242:0] stage1_29;
   wire [206:0] stage1_30;
   wire [242:0] stage1_31;
   wire [149:0] stage1_32;
   wire [70:0] stage1_33;
   wire [62:0] stage2_0;
   wire [55:0] stage2_1;
   wire [94:0] stage2_2;
   wire [76:0] stage2_3;
   wire [118:0] stage2_4;
   wire [93:0] stage2_5;
   wire [95:0] stage2_6;
   wire [108:0] stage2_7;
   wire [97:0] stage2_8;
   wire [107:0] stage2_9;
   wire [94:0] stage2_10;
   wire [115:0] stage2_11;
   wire [101:0] stage2_12;
   wire [123:0] stage2_13;
   wire [69:0] stage2_14;
   wire [97:0] stage2_15;
   wire [124:0] stage2_16;
   wire [127:0] stage2_17;
   wire [72:0] stage2_18;
   wire [97:0] stage2_19;
   wire [109:0] stage2_20;
   wire [124:0] stage2_21;
   wire [94:0] stage2_22;
   wire [122:0] stage2_23;
   wire [89:0] stage2_24;
   wire [102:0] stage2_25;
   wire [99:0] stage2_26;
   wire [84:0] stage2_27;
   wire [170:0] stage2_28;
   wire [142:0] stage2_29;
   wire [91:0] stage2_30;
   wire [101:0] stage2_31;
   wire [73:0] stage2_32;
   wire [59:0] stage2_33;
   wire [34:0] stage2_34;
   wire [11:0] stage2_35;
   wire [10:0] stage3_0;
   wire [25:0] stage3_1;
   wire [35:0] stage3_2;
   wire [27:0] stage3_3;
   wire [46:0] stage3_4;
   wire [58:0] stage3_5;
   wire [37:0] stage3_6;
   wire [46:0] stage3_7;
   wire [92:0] stage3_8;
   wire [49:0] stage3_9;
   wire [37:0] stage3_10;
   wire [54:0] stage3_11;
   wire [46:0] stage3_12;
   wire [36:0] stage3_13;
   wire [55:0] stage3_14;
   wire [70:0] stage3_15;
   wire [66:0] stage3_16;
   wire [76:0] stage3_17;
   wire [34:0] stage3_18;
   wire [69:0] stage3_19;
   wire [29:0] stage3_20;
   wire [62:0] stage3_21;
   wire [50:0] stage3_22;
   wire [45:0] stage3_23;
   wire [60:0] stage3_24;
   wire [48:0] stage3_25;
   wire [50:0] stage3_26;
   wire [54:0] stage3_27;
   wire [73:0] stage3_28;
   wire [57:0] stage3_29;
   wire [70:0] stage3_30;
   wire [57:0] stage3_31;
   wire [57:0] stage3_32;
   wire [26:0] stage3_33;
   wire [26:0] stage3_34;
   wire [12:0] stage3_35;
   wire [5:0] stage3_36;
   wire [1:0] stage3_37;
   wire [10:0] stage4_0;
   wire [15:0] stage4_1;
   wire [12:0] stage4_2;
   wire [22:0] stage4_3;
   wire [23:0] stage4_4;
   wire [45:0] stage4_5;
   wire [22:0] stage4_6;
   wire [14:0] stage4_7;
   wire [28:0] stage4_8;
   wire [41:0] stage4_9;
   wire [17:0] stage4_10;
   wire [42:0] stage4_11;
   wire [23:0] stage4_12;
   wire [18:0] stage4_13;
   wire [34:0] stage4_14;
   wire [38:0] stage4_15;
   wire [19:0] stage4_16;
   wire [42:0] stage4_17;
   wire [28:0] stage4_18;
   wire [31:0] stage4_19;
   wire [18:0] stage4_20;
   wire [18:0] stage4_21;
   wire [30:0] stage4_22;
   wire [37:0] stage4_23;
   wire [29:0] stage4_24;
   wire [18:0] stage4_25;
   wire [22:0] stage4_26;
   wire [26:0] stage4_27;
   wire [24:0] stage4_28;
   wire [25:0] stage4_29;
   wire [26:0] stage4_30;
   wire [30:0] stage4_31;
   wire [42:0] stage4_32;
   wire [18:0] stage4_33;
   wire [12:0] stage4_34;
   wire [14:0] stage4_35;
   wire [10:0] stage4_36;
   wire [2:0] stage4_37;
   wire [10:0] stage5_0;
   wire [10:0] stage5_1;
   wire [9:0] stage5_2;
   wire [5:0] stage5_3;
   wire [9:0] stage5_4;
   wire [10:0] stage5_5;
   wire [12:0] stage5_6;
   wire [19:0] stage5_7;
   wire [9:0] stage5_8;
   wire [10:0] stage5_9;
   wire [12:0] stage5_10;
   wire [15:0] stage5_11;
   wire [10:0] stage5_12;
   wire [14:0] stage5_13;
   wire [9:0] stage5_14;
   wire [12:0] stage5_15;
   wire [14:0] stage5_16;
   wire [14:0] stage5_17;
   wire [16:0] stage5_18;
   wire [23:0] stage5_19;
   wire [13:0] stage5_20;
   wire [8:0] stage5_21;
   wire [16:0] stage5_22;
   wire [9:0] stage5_23;
   wire [13:0] stage5_24;
   wire [11:0] stage5_25;
   wire [13:0] stage5_26;
   wire [13:0] stage5_27;
   wire [6:0] stage5_28;
   wire [12:0] stage5_29;
   wire [16:0] stage5_30;
   wire [12:0] stage5_31;
   wire [25:0] stage5_32;
   wire [10:0] stage5_33;
   wire [9:0] stage5_34;
   wire [7:0] stage5_35;
   wire [3:0] stage5_36;
   wire [6:0] stage5_37;
   wire [1:0] stage5_38;
   wire [6:0] stage6_0;
   wire [4:0] stage6_1;
   wire [5:0] stage6_2;
   wire [5:0] stage6_3;
   wire [5:0] stage6_4;
   wire [4:0] stage6_5;
   wire [3:0] stage6_6;
   wire [5:0] stage6_7;
   wire [5:0] stage6_8;
   wire [5:0] stage6_9;
   wire [3:0] stage6_10;
   wire [7:0] stage6_11;
   wire [6:0] stage6_12;
   wire [8:0] stage6_13;
   wire [5:0] stage6_14;
   wire [3:0] stage6_15;
   wire [5:0] stage6_16;
   wire [9:0] stage6_17;
   wire [5:0] stage6_18;
   wire [14:0] stage6_19;
   wire [5:0] stage6_20;
   wire [12:0] stage6_21;
   wire [7:0] stage6_22;
   wire [3:0] stage6_23;
   wire [5:0] stage6_24;
   wire [5:0] stage6_25;
   wire [4:0] stage6_26;
   wire [7:0] stage6_27;
   wire [4:0] stage6_28;
   wire [3:0] stage6_29;
   wire [5:0] stage6_30;
   wire [7:0] stage6_31;
   wire [5:0] stage6_32;
   wire [5:0] stage6_33;
   wire [9:0] stage6_34;
   wire [5:0] stage6_35;
   wire [2:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;
   wire [1:0] stage6_39;
   wire [0:0] stage6_40;
   wire [6:0] stage7_0;
   wire [0:0] stage7_1;
   wire [6:0] stage7_2;
   wire [0:0] stage7_3;
   wire [6:0] stage7_4;
   wire [1:0] stage7_5;
   wire [3:0] stage7_6;
   wire [1:0] stage7_7;
   wire [6:0] stage7_8;
   wire [0:0] stage7_9;
   wire [4:0] stage7_10;
   wire [2:0] stage7_11;
   wire [3:0] stage7_12;
   wire [1:0] stage7_13;
   wire [6:0] stage7_14;
   wire [5:0] stage7_15;
   wire [1:0] stage7_16;
   wire [3:0] stage7_17;
   wire [1:0] stage7_18;
   wire [4:0] stage7_19;
   wire [5:0] stage7_20;
   wire [2:0] stage7_21;
   wire [5:0] stage7_22;
   wire [6:0] stage7_23;
   wire [0:0] stage7_24;
   wire [1:0] stage7_25;
   wire [2:0] stage7_26;
   wire [2:0] stage7_27;
   wire [6:0] stage7_28;
   wire [4:0] stage7_29;
   wire [0:0] stage7_30;
   wire [8:0] stage7_31;
   wire [0:0] stage7_32;
   wire [1:0] stage7_33;
   wire [6:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [3:0] stage7_37;
   wire [2:0] stage7_38;
   wire [1:0] stage7_39;
   wire [0:0] stage7_40;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [1:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [1:0] stage8_39;
   wire [0:0] stage8_40;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[11]},
      {stage0_3[22]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[12]},
      {stage0_3[23]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[13]},
      {stage0_3[24]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_2[14]},
      {stage0_3[25]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_2[15]},
      {stage0_3[26]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_2[16]},
      {stage0_3[27]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_2[17]},
      {stage0_3[28]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_2[18]},
      {stage0_3[29]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86]},
      {stage0_2[19]},
      {stage0_3[30]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92]},
      {stage0_2[20]},
      {stage0_3[31]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98]},
      {stage0_2[21]},
      {stage0_3[32]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104]},
      {stage0_2[22]},
      {stage0_3[33]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110]},
      {stage0_2[23]},
      {stage0_3[34]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116]},
      {stage0_2[24]},
      {stage0_3[35]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122]},
      {stage0_2[25]},
      {stage0_3[36]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127], stage0_1[128]},
      {stage0_2[26]},
      {stage0_3[37]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133], stage0_1[134]},
      {stage0_2[27]},
      {stage0_3[38]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139], stage0_1[140]},
      {stage0_2[28]},
      {stage0_3[39]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145], stage0_1[146]},
      {stage0_2[29]},
      {stage0_3[40]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151], stage0_1[152]},
      {stage0_2[30]},
      {stage0_3[41]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157], stage0_1[158]},
      {stage0_2[31]},
      {stage0_3[42]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163], stage0_1[164]},
      {stage0_2[32]},
      {stage0_3[43]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169], stage0_1[170]},
      {stage0_2[33]},
      {stage0_3[44]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175], stage0_1[176]},
      {stage0_2[34]},
      {stage0_3[45]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182]},
      {stage0_2[35]},
      {stage0_3[46]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188]},
      {stage0_2[36]},
      {stage0_3[47]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194]},
      {stage0_2[37]},
      {stage0_3[48]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200]},
      {stage0_2[38]},
      {stage0_3[49]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206]},
      {stage0_2[39]},
      {stage0_3[50]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212]},
      {stage0_2[40]},
      {stage0_3[51]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218]},
      {stage0_2[41]},
      {stage0_3[52]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261]},
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155]},
      {stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267]},
      {stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161]},
      {stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273]},
      {stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167]},
      {stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279]},
      {stage0_2[168], stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285]},
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179]},
      {stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291]},
      {stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297]},
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191]},
      {stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303]},
      {stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197]},
      {stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309]},
      {stage0_2[198], stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203]},
      {stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315]},
      {stage0_2[204], stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209]},
      {stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321]},
      {stage0_2[210], stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327]},
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221]},
      {stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333]},
      {stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227]},
      {stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339]},
      {stage0_2[228], stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233]},
      {stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345]},
      {stage0_2[234], stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351]},
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357]},
      {stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251]},
      {stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363]},
      {stage0_2[252], stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257]},
      {stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369]},
      {stage0_2[258], stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263]},
      {stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375]},
      {stage0_2[264], stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269]},
      {stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381]},
      {stage0_2[270], stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275]},
      {stage1_4[80],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387]},
      {stage0_2[276], stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281]},
      {stage1_4[81],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393]},
      {stage0_2[282], stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287]},
      {stage1_4[82],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399]},
      {stage0_2[288], stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage1_4[83],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405]},
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage1_4[84],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411]},
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage1_4[85],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417]},
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage1_4[86],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423]},
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage1_4[87],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc606_5 gpc88 (
      {stage0_0[424], stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429]},
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage1_4[88],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc606_5 gpc89 (
      {stage0_0[430], stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435]},
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage1_4[89],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc606_5 gpc90 (
      {stage0_0[436], stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441]},
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage1_4[90],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc606_5 gpc91 (
      {stage0_0[442], stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447]},
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage1_4[91],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc606_5 gpc92 (
      {stage0_0[448], stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453]},
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage1_4[92],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc606_5 gpc93 (
      {stage0_0[454], stage0_0[455], stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459]},
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage1_4[93],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc606_5 gpc94 (
      {stage0_0[460], stage0_0[461], stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465]},
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage1_4[94],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc606_5 gpc95 (
      {stage0_0[466], stage0_0[467], stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471]},
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage1_4[95],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc606_5 gpc96 (
      {stage0_0[472], stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477]},
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage1_4[96],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc606_5 gpc97 (
      {stage0_0[478], stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483]},
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage1_4[97],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc606_5 gpc98 (
      {stage0_0[484], stage0_0[485], stage0_0[486], stage0_0[487], stage0_0[488], stage0_0[489]},
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage1_4[98],stage1_3[98],stage1_2[98],stage1_1[98],stage1_0[98]}
   );
   gpc606_5 gpc99 (
      {stage0_0[490], stage0_0[491], stage0_0[492], stage0_0[493], stage0_0[494], stage0_0[495]},
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage1_4[99],stage1_3[99],stage1_2[99],stage1_1[99],stage1_0[99]}
   );
   gpc606_5 gpc100 (
      {stage0_0[496], stage0_0[497], stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501]},
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394], stage0_2[395]},
      {stage1_4[100],stage1_3[100],stage1_2[100],stage1_1[100],stage1_0[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224]},
      {stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58]},
      {stage1_5[0],stage1_4[101],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230]},
      {stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64]},
      {stage1_5[1],stage1_4[102],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236]},
      {stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70]},
      {stage1_5[2],stage1_4[103],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241], stage0_1[242]},
      {stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage1_5[3],stage1_4[104],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247], stage0_1[248]},
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82]},
      {stage1_5[4],stage1_4[105],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253], stage0_1[254]},
      {stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88]},
      {stage1_5[5],stage1_4[106],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259], stage0_1[260]},
      {stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94]},
      {stage1_5[6],stage1_4[107],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265], stage0_1[266]},
      {stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100]},
      {stage1_5[7],stage1_4[108],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271], stage0_1[272]},
      {stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage1_5[8],stage1_4[109],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277], stage0_1[278]},
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112]},
      {stage1_5[9],stage1_4[110],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283], stage0_1[284]},
      {stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage1_5[10],stage1_4[111],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289], stage0_1[290]},
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124]},
      {stage1_5[11],stage1_4[112],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295], stage0_1[296]},
      {stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130]},
      {stage1_5[12],stage1_4[113],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301], stage0_1[302]},
      {stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136]},
      {stage1_5[13],stage1_4[114],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307], stage0_1[308]},
      {stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142]},
      {stage1_5[14],stage1_4[115],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313], stage0_1[314]},
      {stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148]},
      {stage1_5[15],stage1_4[116],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319], stage0_1[320]},
      {stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage1_5[16],stage1_4[117],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325], stage0_1[326]},
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160]},
      {stage1_5[17],stage1_4[118],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331], stage0_1[332]},
      {stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166]},
      {stage1_5[18],stage1_4[119],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337], stage0_1[338]},
      {stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172]},
      {stage1_5[19],stage1_4[120],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343], stage0_1[344]},
      {stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178]},
      {stage1_5[20],stage1_4[121],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349], stage0_1[350]},
      {stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage1_5[21],stage1_4[122],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355], stage0_1[356]},
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190]},
      {stage1_5[22],stage1_4[123],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361], stage0_1[362]},
      {stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage1_5[23],stage1_4[124],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368]},
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202]},
      {stage1_5[24],stage1_4[125],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373], stage0_1[374]},
      {stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208]},
      {stage1_5[25],stage1_4[126],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379], stage0_1[380]},
      {stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage1_5[26],stage1_4[127],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385], stage0_1[386]},
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220]},
      {stage1_5[27],stage1_4[128],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391], stage0_1[392]},
      {stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage1_5[28],stage1_4[129],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397], stage0_1[398]},
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage1_5[29],stage1_4[130],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403], stage0_1[404]},
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238]},
      {stage1_5[30],stage1_4[131],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409], stage0_1[410]},
      {stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage1_5[31],stage1_4[132],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415], stage0_1[416]},
      {stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250]},
      {stage1_5[32],stage1_4[133],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421], stage0_1[422]},
      {stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256]},
      {stage1_5[33],stage1_4[134],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427], stage0_1[428]},
      {stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262]},
      {stage1_5[34],stage1_4[135],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433], stage0_1[434]},
      {stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268]},
      {stage1_5[35],stage1_4[136],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439], stage0_1[440]},
      {stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274]},
      {stage1_5[36],stage1_4[137],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445], stage0_1[446]},
      {stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280]},
      {stage1_5[37],stage1_4[138],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451], stage0_1[452]},
      {stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286]},
      {stage1_5[38],stage1_4[139],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc615_5 gpc140 (
      {stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399], stage0_2[400]},
      {stage0_3[287]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[39],stage1_4[140],stage1_3[140],stage1_2[140]}
   );
   gpc615_5 gpc141 (
      {stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404], stage0_2[405]},
      {stage0_3[288]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[40],stage1_4[141],stage1_3[141],stage1_2[141]}
   );
   gpc615_5 gpc142 (
      {stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409], stage0_2[410]},
      {stage0_3[289]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[41],stage1_4[142],stage1_3[142],stage1_2[142]}
   );
   gpc615_5 gpc143 (
      {stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414], stage0_2[415]},
      {stage0_3[290]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[42],stage1_4[143],stage1_3[143],stage1_2[143]}
   );
   gpc615_5 gpc144 (
      {stage0_2[416], stage0_2[417], stage0_2[418], stage0_2[419], stage0_2[420]},
      {stage0_3[291]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[43],stage1_4[144],stage1_3[144],stage1_2[144]}
   );
   gpc615_5 gpc145 (
      {stage0_2[421], stage0_2[422], stage0_2[423], stage0_2[424], stage0_2[425]},
      {stage0_3[292]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[44],stage1_4[145],stage1_3[145],stage1_2[145]}
   );
   gpc615_5 gpc146 (
      {stage0_2[426], stage0_2[427], stage0_2[428], stage0_2[429], stage0_2[430]},
      {stage0_3[293]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[45],stage1_4[146],stage1_3[146],stage1_2[146]}
   );
   gpc615_5 gpc147 (
      {stage0_2[431], stage0_2[432], stage0_2[433], stage0_2[434], stage0_2[435]},
      {stage0_3[294]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[46],stage1_4[147],stage1_3[147],stage1_2[147]}
   );
   gpc615_5 gpc148 (
      {stage0_2[436], stage0_2[437], stage0_2[438], stage0_2[439], stage0_2[440]},
      {stage0_3[295]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[47],stage1_4[148],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[441], stage0_2[442], stage0_2[443], stage0_2[444], stage0_2[445]},
      {stage0_3[296]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[48],stage1_4[149],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[446], stage0_2[447], stage0_2[448], stage0_2[449], stage0_2[450]},
      {stage0_3[297]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[49],stage1_4[150],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[451], stage0_2[452], stage0_2[453], stage0_2[454], stage0_2[455]},
      {stage0_3[298]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[50],stage1_4[151],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[456], stage0_2[457], stage0_2[458], stage0_2[459], stage0_2[460]},
      {stage0_3[299]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[51],stage1_4[152],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[461], stage0_2[462], stage0_2[463], stage0_2[464], stage0_2[465]},
      {stage0_3[300]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[52],stage1_4[153],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[466], stage0_2[467], stage0_2[468], stage0_2[469], stage0_2[470]},
      {stage0_3[301]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[53],stage1_4[154],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[471], stage0_2[472], stage0_2[473], stage0_2[474], stage0_2[475]},
      {stage0_3[302]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[54],stage1_4[155],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[476], stage0_2[477], stage0_2[478], stage0_2[479], stage0_2[480]},
      {stage0_3[303]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[55],stage1_4[156],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308]},
      {stage0_4[102]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[17],stage1_5[56],stage1_4[157],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313]},
      {stage0_4[103]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[18],stage1_5[57],stage1_4[158],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[314], stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318]},
      {stage0_4[104]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[19],stage1_5[58],stage1_4[159],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[319], stage0_3[320], stage0_3[321], stage0_3[322], stage0_3[323]},
      {stage0_4[105]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[20],stage1_5[59],stage1_4[160],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[324], stage0_3[325], stage0_3[326], stage0_3[327], stage0_3[328]},
      {stage0_4[106]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[21],stage1_5[60],stage1_4[161],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332], stage0_3[333]},
      {stage0_4[107]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[22],stage1_5[61],stage1_4[162],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[334], stage0_3[335], stage0_3[336], stage0_3[337], stage0_3[338]},
      {stage0_4[108]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[23],stage1_5[62],stage1_4[163],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343]},
      {stage0_4[109]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[24],stage1_5[63],stage1_4[164],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage0_4[110]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[25],stage1_5[64],stage1_4[165],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[349], stage0_3[350], stage0_3[351], stage0_3[352], stage0_3[353]},
      {stage0_4[111]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[26],stage1_5[65],stage1_4[166],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[354], stage0_3[355], stage0_3[356], stage0_3[357], stage0_3[358]},
      {stage0_4[112]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[27],stage1_5[66],stage1_4[167],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362], stage0_3[363]},
      {stage0_4[113]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[28],stage1_5[67],stage1_4[168],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage0_4[114]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[29],stage1_5[68],stage1_4[169],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373]},
      {stage0_4[115]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[30],stage1_5[69],stage1_4[170],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[374], stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378]},
      {stage0_4[116]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[31],stage1_5[70],stage1_4[171],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[379], stage0_3[380], stage0_3[381], stage0_3[382], stage0_3[383]},
      {stage0_4[117]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[32],stage1_5[71],stage1_4[172],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[384], stage0_3[385], stage0_3[386], stage0_3[387], stage0_3[388]},
      {stage0_4[118]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[33],stage1_5[72],stage1_4[173],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392], stage0_3[393]},
      {stage0_4[119]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[34],stage1_5[73],stage1_4[174],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage0_4[120]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[35],stage1_5[74],stage1_4[175],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403]},
      {stage0_4[121]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[36],stage1_5[75],stage1_4[176],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[404], stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408]},
      {stage0_4[122]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[37],stage1_5[76],stage1_4[177],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[409], stage0_3[410], stage0_3[411], stage0_3[412], stage0_3[413]},
      {stage0_4[123]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[38],stage1_5[77],stage1_4[178],stage1_3[178]}
   );
   gpc606_5 gpc179 (
      {stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[22],stage1_6[39],stage1_5[78],stage1_4[179]}
   );
   gpc606_5 gpc180 (
      {stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[23],stage1_6[40],stage1_5[79],stage1_4[180]}
   );
   gpc606_5 gpc181 (
      {stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[24],stage1_6[41],stage1_5[80],stage1_4[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[25],stage1_6[42],stage1_5[81],stage1_4[182]}
   );
   gpc606_5 gpc183 (
      {stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[26],stage1_6[43],stage1_5[82],stage1_4[183]}
   );
   gpc606_5 gpc184 (
      {stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[27],stage1_6[44],stage1_5[83],stage1_4[184]}
   );
   gpc606_5 gpc185 (
      {stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[28],stage1_6[45],stage1_5[84],stage1_4[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[29],stage1_6[46],stage1_5[85],stage1_4[186]}
   );
   gpc606_5 gpc187 (
      {stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[30],stage1_6[47],stage1_5[86],stage1_4[187]}
   );
   gpc606_5 gpc188 (
      {stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[31],stage1_6[48],stage1_5[87],stage1_4[188]}
   );
   gpc606_5 gpc189 (
      {stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[32],stage1_6[49],stage1_5[88],stage1_4[189]}
   );
   gpc606_5 gpc190 (
      {stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[33],stage1_6[50],stage1_5[89],stage1_4[190]}
   );
   gpc606_5 gpc191 (
      {stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[34],stage1_6[51],stage1_5[90],stage1_4[191]}
   );
   gpc606_5 gpc192 (
      {stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[35],stage1_6[52],stage1_5[91],stage1_4[192]}
   );
   gpc606_5 gpc193 (
      {stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[36],stage1_6[53],stage1_5[92],stage1_4[193]}
   );
   gpc606_5 gpc194 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[37],stage1_6[54],stage1_5[93],stage1_4[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[38],stage1_6[55],stage1_5[94],stage1_4[195]}
   );
   gpc606_5 gpc196 (
      {stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[39],stage1_6[56],stage1_5[95],stage1_4[196]}
   );
   gpc606_5 gpc197 (
      {stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[40],stage1_6[57],stage1_5[96],stage1_4[197]}
   );
   gpc606_5 gpc198 (
      {stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[41],stage1_6[58],stage1_5[97],stage1_4[198]}
   );
   gpc606_5 gpc199 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[42],stage1_6[59],stage1_5[98],stage1_4[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[43],stage1_6[60],stage1_5[99],stage1_4[200]}
   );
   gpc606_5 gpc201 (
      {stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260], stage0_4[261]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[44],stage1_6[61],stage1_5[100],stage1_4[201]}
   );
   gpc606_5 gpc202 (
      {stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266], stage0_4[267]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[45],stage1_6[62],stage1_5[101],stage1_4[202]}
   );
   gpc606_5 gpc203 (
      {stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272], stage0_4[273]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[46],stage1_6[63],stage1_5[102],stage1_4[203]}
   );
   gpc606_5 gpc204 (
      {stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278], stage0_4[279]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[47],stage1_6[64],stage1_5[103],stage1_4[204]}
   );
   gpc606_5 gpc205 (
      {stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284], stage0_4[285]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[48],stage1_6[65],stage1_5[104],stage1_4[205]}
   );
   gpc606_5 gpc206 (
      {stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290], stage0_4[291]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[49],stage1_6[66],stage1_5[105],stage1_4[206]}
   );
   gpc606_5 gpc207 (
      {stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296], stage0_4[297]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[50],stage1_6[67],stage1_5[106],stage1_4[207]}
   );
   gpc606_5 gpc208 (
      {stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302], stage0_4[303]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[51],stage1_6[68],stage1_5[107],stage1_4[208]}
   );
   gpc606_5 gpc209 (
      {stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308], stage0_4[309]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[52],stage1_6[69],stage1_5[108],stage1_4[209]}
   );
   gpc606_5 gpc210 (
      {stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314], stage0_4[315]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[53],stage1_6[70],stage1_5[109],stage1_4[210]}
   );
   gpc606_5 gpc211 (
      {stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320], stage0_4[321]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[54],stage1_6[71],stage1_5[110],stage1_4[211]}
   );
   gpc606_5 gpc212 (
      {stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326], stage0_4[327]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[55],stage1_6[72],stage1_5[111],stage1_4[212]}
   );
   gpc606_5 gpc213 (
      {stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332], stage0_4[333]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[56],stage1_6[73],stage1_5[112],stage1_4[213]}
   );
   gpc606_5 gpc214 (
      {stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338], stage0_4[339]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[57],stage1_6[74],stage1_5[113],stage1_4[214]}
   );
   gpc606_5 gpc215 (
      {stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344], stage0_4[345]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[58],stage1_6[75],stage1_5[114],stage1_4[215]}
   );
   gpc606_5 gpc216 (
      {stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350], stage0_4[351]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[59],stage1_6[76],stage1_5[115],stage1_4[216]}
   );
   gpc606_5 gpc217 (
      {stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356], stage0_4[357]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[60],stage1_6[77],stage1_5[116],stage1_4[217]}
   );
   gpc606_5 gpc218 (
      {stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362], stage0_4[363]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[61],stage1_6[78],stage1_5[117],stage1_4[218]}
   );
   gpc606_5 gpc219 (
      {stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368], stage0_4[369]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[62],stage1_6[79],stage1_5[118],stage1_4[219]}
   );
   gpc606_5 gpc220 (
      {stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374], stage0_4[375]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[63],stage1_6[80],stage1_5[119],stage1_4[220]}
   );
   gpc606_5 gpc221 (
      {stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380], stage0_4[381]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[64],stage1_6[81],stage1_5[120],stage1_4[221]}
   );
   gpc606_5 gpc222 (
      {stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386], stage0_4[387]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[65],stage1_6[82],stage1_5[121],stage1_4[222]}
   );
   gpc606_5 gpc223 (
      {stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392], stage0_4[393]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[66],stage1_6[83],stage1_5[122],stage1_4[223]}
   );
   gpc606_5 gpc224 (
      {stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398], stage0_4[399]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[67],stage1_6[84],stage1_5[123],stage1_4[224]}
   );
   gpc606_5 gpc225 (
      {stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404], stage0_4[405]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[68],stage1_6[85],stage1_5[124],stage1_4[225]}
   );
   gpc606_5 gpc226 (
      {stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410], stage0_4[411]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[69],stage1_6[86],stage1_5[125],stage1_4[226]}
   );
   gpc606_5 gpc227 (
      {stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416], stage0_4[417]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[70],stage1_6[87],stage1_5[126],stage1_4[227]}
   );
   gpc606_5 gpc228 (
      {stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421], stage0_4[422], stage0_4[423]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[71],stage1_6[88],stage1_5[127],stage1_4[228]}
   );
   gpc606_5 gpc229 (
      {stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427], stage0_4[428], stage0_4[429]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[72],stage1_6[89],stage1_5[128],stage1_4[229]}
   );
   gpc606_5 gpc230 (
      {stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[73],stage1_6[90],stage1_5[129],stage1_4[230]}
   );
   gpc606_5 gpc231 (
      {stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[74],stage1_6[91],stage1_5[130],stage1_4[231]}
   );
   gpc606_5 gpc232 (
      {stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446], stage0_4[447]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[75],stage1_6[92],stage1_5[131],stage1_4[232]}
   );
   gpc606_5 gpc233 (
      {stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451], stage0_4[452], stage0_4[453]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[76],stage1_6[93],stage1_5[132],stage1_4[233]}
   );
   gpc606_5 gpc234 (
      {stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459]},
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335]},
      {stage1_8[55],stage1_7[77],stage1_6[94],stage1_5[133],stage1_4[234]}
   );
   gpc606_5 gpc235 (
      {stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465]},
      {stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage1_8[56],stage1_7[78],stage1_6[95],stage1_5[134],stage1_4[235]}
   );
   gpc606_5 gpc236 (
      {stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471]},
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346], stage0_6[347]},
      {stage1_8[57],stage1_7[79],stage1_6[96],stage1_5[135],stage1_4[236]}
   );
   gpc615_5 gpc237 (
      {stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476]},
      {stage0_5[132]},
      {stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353]},
      {stage1_8[58],stage1_7[80],stage1_6[97],stage1_5[136],stage1_4[237]}
   );
   gpc615_5 gpc238 (
      {stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_5[133]},
      {stage0_6[354], stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage1_8[59],stage1_7[81],stage1_6[98],stage1_5[137],stage1_4[238]}
   );
   gpc615_5 gpc239 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486]},
      {stage0_5[134]},
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365]},
      {stage1_8[60],stage1_7[82],stage1_6[99],stage1_5[138],stage1_4[239]}
   );
   gpc615_5 gpc240 (
      {stage0_4[487], stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491]},
      {stage0_5[135]},
      {stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage1_8[61],stage1_7[83],stage1_6[100],stage1_5[139],stage1_4[240]}
   );
   gpc615_5 gpc241 (
      {stage0_4[492], stage0_4[493], stage0_4[494], stage0_4[495], stage0_4[496]},
      {stage0_5[136]},
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376], stage0_6[377]},
      {stage1_8[62],stage1_7[84],stage1_6[101],stage1_5[140],stage1_4[241]}
   );
   gpc615_5 gpc242 (
      {stage0_4[497], stage0_4[498], stage0_4[499], stage0_4[500], stage0_4[501]},
      {stage0_5[137]},
      {stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383]},
      {stage1_8[63],stage1_7[85],stage1_6[102],stage1_5[141],stage1_4[242]}
   );
   gpc615_5 gpc243 (
      {stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505], stage0_4[506]},
      {stage0_5[138]},
      {stage0_6[384], stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage1_8[64],stage1_7[86],stage1_6[103],stage1_5[142],stage1_4[243]}
   );
   gpc615_5 gpc244 (
      {stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_5[139]},
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395]},
      {stage1_8[65],stage1_7[87],stage1_6[104],stage1_5[143],stage1_4[244]}
   );
   gpc606_5 gpc245 (
      {stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[66],stage1_7[88],stage1_6[105],stage1_5[144]}
   );
   gpc606_5 gpc246 (
      {stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[67],stage1_7[89],stage1_6[106],stage1_5[145]}
   );
   gpc606_5 gpc247 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[68],stage1_7[90],stage1_6[107],stage1_5[146]}
   );
   gpc606_5 gpc248 (
      {stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[69],stage1_7[91],stage1_6[108],stage1_5[147]}
   );
   gpc606_5 gpc249 (
      {stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[70],stage1_7[92],stage1_6[109],stage1_5[148]}
   );
   gpc606_5 gpc250 (
      {stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[71],stage1_7[93],stage1_6[110],stage1_5[149]}
   );
   gpc606_5 gpc251 (
      {stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[72],stage1_7[94],stage1_6[111],stage1_5[150]}
   );
   gpc606_5 gpc252 (
      {stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[73],stage1_7[95],stage1_6[112],stage1_5[151]}
   );
   gpc606_5 gpc253 (
      {stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[74],stage1_7[96],stage1_6[113],stage1_5[152]}
   );
   gpc606_5 gpc254 (
      {stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[75],stage1_7[97],stage1_6[114],stage1_5[153]}
   );
   gpc606_5 gpc255 (
      {stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[76],stage1_7[98],stage1_6[115],stage1_5[154]}
   );
   gpc606_5 gpc256 (
      {stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[77],stage1_7[99],stage1_6[116],stage1_5[155]}
   );
   gpc606_5 gpc257 (
      {stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[78],stage1_7[100],stage1_6[117],stage1_5[156]}
   );
   gpc606_5 gpc258 (
      {stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[79],stage1_7[101],stage1_6[118],stage1_5[157]}
   );
   gpc606_5 gpc259 (
      {stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[80],stage1_7[102],stage1_6[119],stage1_5[158]}
   );
   gpc606_5 gpc260 (
      {stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[81],stage1_7[103],stage1_6[120],stage1_5[159]}
   );
   gpc606_5 gpc261 (
      {stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[82],stage1_7[104],stage1_6[121],stage1_5[160]}
   );
   gpc606_5 gpc262 (
      {stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[83],stage1_7[105],stage1_6[122],stage1_5[161]}
   );
   gpc606_5 gpc263 (
      {stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[84],stage1_7[106],stage1_6[123],stage1_5[162]}
   );
   gpc606_5 gpc264 (
      {stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258], stage0_5[259]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[85],stage1_7[107],stage1_6[124],stage1_5[163]}
   );
   gpc606_5 gpc265 (
      {stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264], stage0_5[265]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[86],stage1_7[108],stage1_6[125],stage1_5[164]}
   );
   gpc606_5 gpc266 (
      {stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270], stage0_5[271]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[87],stage1_7[109],stage1_6[126],stage1_5[165]}
   );
   gpc606_5 gpc267 (
      {stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276], stage0_5[277]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[88],stage1_7[110],stage1_6[127],stage1_5[166]}
   );
   gpc606_5 gpc268 (
      {stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281], stage0_5[282], stage0_5[283]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[89],stage1_7[111],stage1_6[128],stage1_5[167]}
   );
   gpc606_5 gpc269 (
      {stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287], stage0_5[288], stage0_5[289]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[90],stage1_7[112],stage1_6[129],stage1_5[168]}
   );
   gpc606_5 gpc270 (
      {stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293], stage0_5[294], stage0_5[295]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[91],stage1_7[113],stage1_6[130],stage1_5[169]}
   );
   gpc606_5 gpc271 (
      {stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300], stage0_5[301]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[92],stage1_7[114],stage1_6[131],stage1_5[170]}
   );
   gpc606_5 gpc272 (
      {stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306], stage0_5[307]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[93],stage1_7[115],stage1_6[132],stage1_5[171]}
   );
   gpc606_5 gpc273 (
      {stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311], stage0_5[312], stage0_5[313]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[94],stage1_7[116],stage1_6[133],stage1_5[172]}
   );
   gpc606_5 gpc274 (
      {stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317], stage0_5[318], stage0_5[319]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[95],stage1_7[117],stage1_6[134],stage1_5[173]}
   );
   gpc606_5 gpc275 (
      {stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323], stage0_5[324], stage0_5[325]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[96],stage1_7[118],stage1_6[135],stage1_5[174]}
   );
   gpc606_5 gpc276 (
      {stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330], stage0_5[331]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[97],stage1_7[119],stage1_6[136],stage1_5[175]}
   );
   gpc606_5 gpc277 (
      {stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336], stage0_5[337]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[98],stage1_7[120],stage1_6[137],stage1_5[176]}
   );
   gpc606_5 gpc278 (
      {stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341], stage0_5[342], stage0_5[343]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[99],stage1_7[121],stage1_6[138],stage1_5[177]}
   );
   gpc606_5 gpc279 (
      {stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347], stage0_5[348], stage0_5[349]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[100],stage1_7[122],stage1_6[139],stage1_5[178]}
   );
   gpc606_5 gpc280 (
      {stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353], stage0_5[354], stage0_5[355]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[101],stage1_7[123],stage1_6[140],stage1_5[179]}
   );
   gpc606_5 gpc281 (
      {stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359], stage0_5[360], stage0_5[361]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[102],stage1_7[124],stage1_6[141],stage1_5[180]}
   );
   gpc606_5 gpc282 (
      {stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365], stage0_5[366], stage0_5[367]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[103],stage1_7[125],stage1_6[142],stage1_5[181]}
   );
   gpc606_5 gpc283 (
      {stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371], stage0_5[372], stage0_5[373]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[104],stage1_7[126],stage1_6[143],stage1_5[182]}
   );
   gpc606_5 gpc284 (
      {stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377], stage0_5[378], stage0_5[379]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[105],stage1_7[127],stage1_6[144],stage1_5[183]}
   );
   gpc606_5 gpc285 (
      {stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383], stage0_5[384], stage0_5[385]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[106],stage1_7[128],stage1_6[145],stage1_5[184]}
   );
   gpc606_5 gpc286 (
      {stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389], stage0_5[390], stage0_5[391]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[107],stage1_7[129],stage1_6[146],stage1_5[185]}
   );
   gpc606_5 gpc287 (
      {stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395], stage0_5[396], stage0_5[397]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[108],stage1_7[130],stage1_6[147],stage1_5[186]}
   );
   gpc606_5 gpc288 (
      {stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401], stage0_5[402], stage0_5[403]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[109],stage1_7[131],stage1_6[148],stage1_5[187]}
   );
   gpc606_5 gpc289 (
      {stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407], stage0_5[408], stage0_5[409]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[110],stage1_7[132],stage1_6[149],stage1_5[188]}
   );
   gpc606_5 gpc290 (
      {stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413], stage0_5[414], stage0_5[415]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[111],stage1_7[133],stage1_6[150],stage1_5[189]}
   );
   gpc606_5 gpc291 (
      {stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419], stage0_5[420], stage0_5[421]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[112],stage1_7[134],stage1_6[151],stage1_5[190]}
   );
   gpc606_5 gpc292 (
      {stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425], stage0_5[426], stage0_5[427]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[113],stage1_7[135],stage1_6[152],stage1_5[191]}
   );
   gpc606_5 gpc293 (
      {stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431], stage0_5[432], stage0_5[433]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[114],stage1_7[136],stage1_6[153],stage1_5[192]}
   );
   gpc606_5 gpc294 (
      {stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437], stage0_5[438], stage0_5[439]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[115],stage1_7[137],stage1_6[154],stage1_5[193]}
   );
   gpc606_5 gpc295 (
      {stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443], stage0_5[444], stage0_5[445]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[116],stage1_7[138],stage1_6[155],stage1_5[194]}
   );
   gpc606_5 gpc296 (
      {stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449], stage0_5[450], stage0_5[451]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[117],stage1_7[139],stage1_6[156],stage1_5[195]}
   );
   gpc606_5 gpc297 (
      {stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455], stage0_5[456], stage0_5[457]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[118],stage1_7[140],stage1_6[157],stage1_5[196]}
   );
   gpc606_5 gpc298 (
      {stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461], stage0_5[462], stage0_5[463]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[119],stage1_7[141],stage1_6[158],stage1_5[197]}
   );
   gpc606_5 gpc299 (
      {stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467], stage0_5[468], stage0_5[469]},
      {stage0_7[324], stage0_7[325], stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329]},
      {stage1_9[54],stage1_8[120],stage1_7[142],stage1_6[159],stage1_5[198]}
   );
   gpc606_5 gpc300 (
      {stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473], stage0_5[474], stage0_5[475]},
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage1_9[55],stage1_8[121],stage1_7[143],stage1_6[160],stage1_5[199]}
   );
   gpc606_5 gpc301 (
      {stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479], stage0_5[480], stage0_5[481]},
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340], stage0_7[341]},
      {stage1_9[56],stage1_8[122],stage1_7[144],stage1_6[161],stage1_5[200]}
   );
   gpc606_5 gpc302 (
      {stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485], stage0_5[486], stage0_5[487]},
      {stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345], stage0_7[346], stage0_7[347]},
      {stage1_9[57],stage1_8[123],stage1_7[145],stage1_6[162],stage1_5[201]}
   );
   gpc606_5 gpc303 (
      {stage0_5[488], stage0_5[489], stage0_5[490], stage0_5[491], stage0_5[492], stage0_5[493]},
      {stage0_7[348], stage0_7[349], stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353]},
      {stage1_9[58],stage1_8[124],stage1_7[146],stage1_6[163],stage1_5[202]}
   );
   gpc606_5 gpc304 (
      {stage0_5[494], stage0_5[495], stage0_5[496], stage0_5[497], stage0_5[498], stage0_5[499]},
      {stage0_7[354], stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage1_9[59],stage1_8[125],stage1_7[147],stage1_6[164],stage1_5[203]}
   );
   gpc606_5 gpc305 (
      {stage0_5[500], stage0_5[501], stage0_5[502], stage0_5[503], stage0_5[504], stage0_5[505]},
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage1_9[60],stage1_8[126],stage1_7[148],stage1_6[165],stage1_5[204]}
   );
   gpc606_5 gpc306 (
      {stage0_5[506], stage0_5[507], stage0_5[508], stage0_5[509], stage0_5[510], stage0_5[511]},
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370], stage0_7[371]},
      {stage1_9[61],stage1_8[127],stage1_7[149],stage1_6[166],stage1_5[205]}
   );
   gpc615_5 gpc307 (
      {stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400]},
      {stage0_7[372]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[62],stage1_8[128],stage1_7[150],stage1_6[167]}
   );
   gpc615_5 gpc308 (
      {stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405]},
      {stage0_7[373]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[63],stage1_8[129],stage1_7[151],stage1_6[168]}
   );
   gpc615_5 gpc309 (
      {stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410]},
      {stage0_7[374]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[64],stage1_8[130],stage1_7[152],stage1_6[169]}
   );
   gpc615_5 gpc310 (
      {stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415]},
      {stage0_7[375]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[65],stage1_8[131],stage1_7[153],stage1_6[170]}
   );
   gpc615_5 gpc311 (
      {stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420]},
      {stage0_7[376]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[66],stage1_8[132],stage1_7[154],stage1_6[171]}
   );
   gpc615_5 gpc312 (
      {stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425]},
      {stage0_7[377]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[67],stage1_8[133],stage1_7[155],stage1_6[172]}
   );
   gpc615_5 gpc313 (
      {stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430]},
      {stage0_7[378]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[68],stage1_8[134],stage1_7[156],stage1_6[173]}
   );
   gpc615_5 gpc314 (
      {stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435]},
      {stage0_7[379]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[69],stage1_8[135],stage1_7[157],stage1_6[174]}
   );
   gpc615_5 gpc315 (
      {stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440]},
      {stage0_7[380]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[70],stage1_8[136],stage1_7[158],stage1_6[175]}
   );
   gpc615_5 gpc316 (
      {stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445]},
      {stage0_7[381]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[71],stage1_8[137],stage1_7[159],stage1_6[176]}
   );
   gpc615_5 gpc317 (
      {stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386]},
      {stage0_8[60]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[10],stage1_9[72],stage1_8[138],stage1_7[160]}
   );
   gpc615_5 gpc318 (
      {stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390], stage0_7[391]},
      {stage0_8[61]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[11],stage1_9[73],stage1_8[139],stage1_7[161]}
   );
   gpc615_5 gpc319 (
      {stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395], stage0_7[396]},
      {stage0_8[62]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[12],stage1_9[74],stage1_8[140],stage1_7[162]}
   );
   gpc615_5 gpc320 (
      {stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400], stage0_7[401]},
      {stage0_8[63]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[13],stage1_9[75],stage1_8[141],stage1_7[163]}
   );
   gpc615_5 gpc321 (
      {stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_8[64]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[14],stage1_9[76],stage1_8[142],stage1_7[164]}
   );
   gpc615_5 gpc322 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411]},
      {stage0_8[65]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[15],stage1_9[77],stage1_8[143],stage1_7[165]}
   );
   gpc615_5 gpc323 (
      {stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416]},
      {stage0_8[66]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[16],stage1_9[78],stage1_8[144],stage1_7[166]}
   );
   gpc615_5 gpc324 (
      {stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420], stage0_7[421]},
      {stage0_8[67]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[17],stage1_9[79],stage1_8[145],stage1_7[167]}
   );
   gpc615_5 gpc325 (
      {stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425], stage0_7[426]},
      {stage0_8[68]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[18],stage1_9[80],stage1_8[146],stage1_7[168]}
   );
   gpc615_5 gpc326 (
      {stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430], stage0_7[431]},
      {stage0_8[69]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[19],stage1_9[81],stage1_8[147],stage1_7[169]}
   );
   gpc615_5 gpc327 (
      {stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_8[70]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[20],stage1_9[82],stage1_8[148],stage1_7[170]}
   );
   gpc615_5 gpc328 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441]},
      {stage0_8[71]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[21],stage1_9[83],stage1_8[149],stage1_7[171]}
   );
   gpc615_5 gpc329 (
      {stage0_7[442], stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446]},
      {stage0_8[72]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[22],stage1_9[84],stage1_8[150],stage1_7[172]}
   );
   gpc615_5 gpc330 (
      {stage0_7[447], stage0_7[448], stage0_7[449], stage0_7[450], stage0_7[451]},
      {stage0_8[73]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[23],stage1_9[85],stage1_8[151],stage1_7[173]}
   );
   gpc615_5 gpc331 (
      {stage0_7[452], stage0_7[453], stage0_7[454], stage0_7[455], stage0_7[456]},
      {stage0_8[74]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[24],stage1_9[86],stage1_8[152],stage1_7[174]}
   );
   gpc615_5 gpc332 (
      {stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460], stage0_7[461]},
      {stage0_8[75]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[25],stage1_9[87],stage1_8[153],stage1_7[175]}
   );
   gpc615_5 gpc333 (
      {stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465], stage0_7[466]},
      {stage0_8[76]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[26],stage1_9[88],stage1_8[154],stage1_7[176]}
   );
   gpc615_5 gpc334 (
      {stage0_7[467], stage0_7[468], stage0_7[469], stage0_7[470], stage0_7[471]},
      {stage0_8[77]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[27],stage1_9[89],stage1_8[155],stage1_7[177]}
   );
   gpc615_5 gpc335 (
      {stage0_7[472], stage0_7[473], stage0_7[474], stage0_7[475], stage0_7[476]},
      {stage0_8[78]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[28],stage1_9[90],stage1_8[156],stage1_7[178]}
   );
   gpc615_5 gpc336 (
      {stage0_7[477], stage0_7[478], stage0_7[479], stage0_7[480], stage0_7[481]},
      {stage0_8[79]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[29],stage1_9[91],stage1_8[157],stage1_7[179]}
   );
   gpc615_5 gpc337 (
      {stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485], stage0_7[486]},
      {stage0_8[80]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[30],stage1_9[92],stage1_8[158],stage1_7[180]}
   );
   gpc615_5 gpc338 (
      {stage0_7[487], stage0_7[488], stage0_7[489], stage0_7[490], stage0_7[491]},
      {stage0_8[81]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[31],stage1_9[93],stage1_8[159],stage1_7[181]}
   );
   gpc615_5 gpc339 (
      {stage0_7[492], stage0_7[493], stage0_7[494], stage0_7[495], stage0_7[496]},
      {stage0_8[82]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[32],stage1_9[94],stage1_8[160],stage1_7[182]}
   );
   gpc615_5 gpc340 (
      {stage0_7[497], stage0_7[498], stage0_7[499], stage0_7[500], stage0_7[501]},
      {stage0_8[83]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[33],stage1_9[95],stage1_8[161],stage1_7[183]}
   );
   gpc615_5 gpc341 (
      {stage0_7[502], stage0_7[503], stage0_7[504], stage0_7[505], stage0_7[506]},
      {stage0_8[84]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[34],stage1_9[96],stage1_8[162],stage1_7[184]}
   );
   gpc615_5 gpc342 (
      {stage0_7[507], stage0_7[508], stage0_7[509], stage0_7[510], stage0_7[511]},
      {stage0_8[85]},
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage1_11[25],stage1_10[35],stage1_9[97],stage1_8[163],stage1_7[185]}
   );
   gpc606_5 gpc343 (
      {stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[26],stage1_10[36],stage1_9[98],stage1_8[164]}
   );
   gpc606_5 gpc344 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[27],stage1_10[37],stage1_9[99],stage1_8[165]}
   );
   gpc606_5 gpc345 (
      {stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[28],stage1_10[38],stage1_9[100],stage1_8[166]}
   );
   gpc606_5 gpc346 (
      {stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[29],stage1_10[39],stage1_9[101],stage1_8[167]}
   );
   gpc606_5 gpc347 (
      {stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[30],stage1_10[40],stage1_9[102],stage1_8[168]}
   );
   gpc606_5 gpc348 (
      {stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[31],stage1_10[41],stage1_9[103],stage1_8[169]}
   );
   gpc606_5 gpc349 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[32],stage1_10[42],stage1_9[104],stage1_8[170]}
   );
   gpc606_5 gpc350 (
      {stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[33],stage1_10[43],stage1_9[105],stage1_8[171]}
   );
   gpc606_5 gpc351 (
      {stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[34],stage1_10[44],stage1_9[106],stage1_8[172]}
   );
   gpc606_5 gpc352 (
      {stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[35],stage1_10[45],stage1_9[107],stage1_8[173]}
   );
   gpc606_5 gpc353 (
      {stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[36],stage1_10[46],stage1_9[108],stage1_8[174]}
   );
   gpc606_5 gpc354 (
      {stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[37],stage1_10[47],stage1_9[109],stage1_8[175]}
   );
   gpc606_5 gpc355 (
      {stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[38],stage1_10[48],stage1_9[110],stage1_8[176]}
   );
   gpc606_5 gpc356 (
      {stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[39],stage1_10[49],stage1_9[111],stage1_8[177]}
   );
   gpc606_5 gpc357 (
      {stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[40],stage1_10[50],stage1_9[112],stage1_8[178]}
   );
   gpc606_5 gpc358 (
      {stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[41],stage1_10[51],stage1_9[113],stage1_8[179]}
   );
   gpc606_5 gpc359 (
      {stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[42],stage1_10[52],stage1_9[114],stage1_8[180]}
   );
   gpc606_5 gpc360 (
      {stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[43],stage1_10[53],stage1_9[115],stage1_8[181]}
   );
   gpc606_5 gpc361 (
      {stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[44],stage1_10[54],stage1_9[116],stage1_8[182]}
   );
   gpc606_5 gpc362 (
      {stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204], stage0_8[205]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[45],stage1_10[55],stage1_9[117],stage1_8[183]}
   );
   gpc606_5 gpc363 (
      {stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[46],stage1_10[56],stage1_9[118],stage1_8[184]}
   );
   gpc606_5 gpc364 (
      {stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[47],stage1_10[57],stage1_9[119],stage1_8[185]}
   );
   gpc606_5 gpc365 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[48],stage1_10[58],stage1_9[120],stage1_8[186]}
   );
   gpc606_5 gpc366 (
      {stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[49],stage1_10[59],stage1_9[121],stage1_8[187]}
   );
   gpc606_5 gpc367 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[50],stage1_10[60],stage1_9[122],stage1_8[188]}
   );
   gpc606_5 gpc368 (
      {stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[51],stage1_10[61],stage1_9[123],stage1_8[189]}
   );
   gpc606_5 gpc369 (
      {stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[52],stage1_10[62],stage1_9[124],stage1_8[190]}
   );
   gpc606_5 gpc370 (
      {stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[53],stage1_10[63],stage1_9[125],stage1_8[191]}
   );
   gpc606_5 gpc371 (
      {stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258], stage0_8[259]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[54],stage1_10[64],stage1_9[126],stage1_8[192]}
   );
   gpc606_5 gpc372 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[55],stage1_10[65],stage1_9[127],stage1_8[193]}
   );
   gpc606_5 gpc373 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[56],stage1_10[66],stage1_9[128],stage1_8[194]}
   );
   gpc606_5 gpc374 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[57],stage1_10[67],stage1_9[129],stage1_8[195]}
   );
   gpc606_5 gpc375 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[58],stage1_10[68],stage1_9[130],stage1_8[196]}
   );
   gpc606_5 gpc376 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[59],stage1_10[69],stage1_9[131],stage1_8[197]}
   );
   gpc606_5 gpc377 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[60],stage1_10[70],stage1_9[132],stage1_8[198]}
   );
   gpc606_5 gpc378 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[61],stage1_10[71],stage1_9[133],stage1_8[199]}
   );
   gpc606_5 gpc379 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[62],stage1_10[72],stage1_9[134],stage1_8[200]}
   );
   gpc606_5 gpc380 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[63],stage1_10[73],stage1_9[135],stage1_8[201]}
   );
   gpc606_5 gpc381 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[64],stage1_10[74],stage1_9[136],stage1_8[202]}
   );
   gpc606_5 gpc382 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[65],stage1_10[75],stage1_9[137],stage1_8[203]}
   );
   gpc606_5 gpc383 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[66],stage1_10[76],stage1_9[138],stage1_8[204]}
   );
   gpc615_5 gpc384 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_9[156]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[67],stage1_10[77],stage1_9[139],stage1_8[205]}
   );
   gpc615_5 gpc385 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_9[157]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[68],stage1_10[78],stage1_9[140],stage1_8[206]}
   );
   gpc615_5 gpc386 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346]},
      {stage0_9[158]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[69],stage1_10[79],stage1_9[141],stage1_8[207]}
   );
   gpc615_5 gpc387 (
      {stage0_8[347], stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351]},
      {stage0_9[159]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[70],stage1_10[80],stage1_9[142],stage1_8[208]}
   );
   gpc615_5 gpc388 (
      {stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355], stage0_8[356]},
      {stage0_9[160]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[71],stage1_10[81],stage1_9[143],stage1_8[209]}
   );
   gpc615_5 gpc389 (
      {stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_9[161]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[72],stage1_10[82],stage1_9[144],stage1_8[210]}
   );
   gpc615_5 gpc390 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_9[162]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[73],stage1_10[83],stage1_9[145],stage1_8[211]}
   );
   gpc615_5 gpc391 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_9[163]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[74],stage1_10[84],stage1_9[146],stage1_8[212]}
   );
   gpc615_5 gpc392 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376]},
      {stage0_9[164]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[75],stage1_10[85],stage1_9[147],stage1_8[213]}
   );
   gpc606_5 gpc393 (
      {stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[50],stage1_11[76],stage1_10[86],stage1_9[148]}
   );
   gpc606_5 gpc394 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[51],stage1_11[77],stage1_10[87],stage1_9[149]}
   );
   gpc606_5 gpc395 (
      {stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[52],stage1_11[78],stage1_10[88],stage1_9[150]}
   );
   gpc606_5 gpc396 (
      {stage0_9[183], stage0_9[184], stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[53],stage1_11[79],stage1_10[89],stage1_9[151]}
   );
   gpc606_5 gpc397 (
      {stage0_9[189], stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[54],stage1_11[80],stage1_10[90],stage1_9[152]}
   );
   gpc606_5 gpc398 (
      {stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[55],stage1_11[81],stage1_10[91],stage1_9[153]}
   );
   gpc606_5 gpc399 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205], stage0_9[206]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[56],stage1_11[82],stage1_10[92],stage1_9[154]}
   );
   gpc606_5 gpc400 (
      {stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210], stage0_9[211], stage0_9[212]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[57],stage1_11[83],stage1_10[93],stage1_9[155]}
   );
   gpc606_5 gpc401 (
      {stage0_9[213], stage0_9[214], stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[58],stage1_11[84],stage1_10[94],stage1_9[156]}
   );
   gpc606_5 gpc402 (
      {stage0_9[219], stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[59],stage1_11[85],stage1_10[95],stage1_9[157]}
   );
   gpc606_5 gpc403 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[60],stage1_11[86],stage1_10[96],stage1_9[158]}
   );
   gpc606_5 gpc404 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235], stage0_9[236]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[61],stage1_11[87],stage1_10[97],stage1_9[159]}
   );
   gpc606_5 gpc405 (
      {stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240], stage0_9[241], stage0_9[242]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[62],stage1_11[88],stage1_10[98],stage1_9[160]}
   );
   gpc606_5 gpc406 (
      {stage0_9[243], stage0_9[244], stage0_9[245], stage0_9[246], stage0_9[247], stage0_9[248]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[63],stage1_11[89],stage1_10[99],stage1_9[161]}
   );
   gpc606_5 gpc407 (
      {stage0_9[249], stage0_9[250], stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[64],stage1_11[90],stage1_10[100],stage1_9[162]}
   );
   gpc606_5 gpc408 (
      {stage0_9[255], stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[65],stage1_11[91],stage1_10[101],stage1_9[163]}
   );
   gpc606_5 gpc409 (
      {stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265], stage0_9[266]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[66],stage1_11[92],stage1_10[102],stage1_9[164]}
   );
   gpc606_5 gpc410 (
      {stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270], stage0_9[271], stage0_9[272]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[67],stage1_11[93],stage1_10[103],stage1_9[165]}
   );
   gpc606_5 gpc411 (
      {stage0_9[273], stage0_9[274], stage0_9[275], stage0_9[276], stage0_9[277], stage0_9[278]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[68],stage1_11[94],stage1_10[104],stage1_9[166]}
   );
   gpc606_5 gpc412 (
      {stage0_9[279], stage0_9[280], stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[69],stage1_11[95],stage1_10[105],stage1_9[167]}
   );
   gpc606_5 gpc413 (
      {stage0_9[285], stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[70],stage1_11[96],stage1_10[106],stage1_9[168]}
   );
   gpc606_5 gpc414 (
      {stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295], stage0_9[296]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[71],stage1_11[97],stage1_10[107],stage1_9[169]}
   );
   gpc606_5 gpc415 (
      {stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300], stage0_9[301], stage0_9[302]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[72],stage1_11[98],stage1_10[108],stage1_9[170]}
   );
   gpc606_5 gpc416 (
      {stage0_9[303], stage0_9[304], stage0_9[305], stage0_9[306], stage0_9[307], stage0_9[308]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[73],stage1_11[99],stage1_10[109],stage1_9[171]}
   );
   gpc606_5 gpc417 (
      {stage0_9[309], stage0_9[310], stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[74],stage1_11[100],stage1_10[110],stage1_9[172]}
   );
   gpc606_5 gpc418 (
      {stage0_9[315], stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[75],stage1_11[101],stage1_10[111],stage1_9[173]}
   );
   gpc606_5 gpc419 (
      {stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325], stage0_9[326]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[76],stage1_11[102],stage1_10[112],stage1_9[174]}
   );
   gpc606_5 gpc420 (
      {stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330], stage0_9[331], stage0_9[332]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[77],stage1_11[103],stage1_10[113],stage1_9[175]}
   );
   gpc606_5 gpc421 (
      {stage0_9[333], stage0_9[334], stage0_9[335], stage0_9[336], stage0_9[337], stage0_9[338]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[78],stage1_11[104],stage1_10[114],stage1_9[176]}
   );
   gpc606_5 gpc422 (
      {stage0_9[339], stage0_9[340], stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[79],stage1_11[105],stage1_10[115],stage1_9[177]}
   );
   gpc606_5 gpc423 (
      {stage0_9[345], stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[80],stage1_11[106],stage1_10[116],stage1_9[178]}
   );
   gpc606_5 gpc424 (
      {stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355], stage0_9[356]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[81],stage1_11[107],stage1_10[117],stage1_9[179]}
   );
   gpc606_5 gpc425 (
      {stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360], stage0_9[361], stage0_9[362]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[82],stage1_11[108],stage1_10[118],stage1_9[180]}
   );
   gpc606_5 gpc426 (
      {stage0_9[363], stage0_9[364], stage0_9[365], stage0_9[366], stage0_9[367], stage0_9[368]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[83],stage1_11[109],stage1_10[119],stage1_9[181]}
   );
   gpc606_5 gpc427 (
      {stage0_9[369], stage0_9[370], stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[84],stage1_11[110],stage1_10[120],stage1_9[182]}
   );
   gpc606_5 gpc428 (
      {stage0_9[375], stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[85],stage1_11[111],stage1_10[121],stage1_9[183]}
   );
   gpc606_5 gpc429 (
      {stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385], stage0_9[386]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[86],stage1_11[112],stage1_10[122],stage1_9[184]}
   );
   gpc606_5 gpc430 (
      {stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390], stage0_9[391], stage0_9[392]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[87],stage1_11[113],stage1_10[123],stage1_9[185]}
   );
   gpc606_5 gpc431 (
      {stage0_9[393], stage0_9[394], stage0_9[395], stage0_9[396], stage0_9[397], stage0_9[398]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[88],stage1_11[114],stage1_10[124],stage1_9[186]}
   );
   gpc615_5 gpc432 (
      {stage0_9[399], stage0_9[400], stage0_9[401], stage0_9[402], stage0_9[403]},
      {stage0_10[300]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[89],stage1_11[115],stage1_10[125],stage1_9[187]}
   );
   gpc615_5 gpc433 (
      {stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407], stage0_9[408]},
      {stage0_10[301]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[90],stage1_11[116],stage1_10[126],stage1_9[188]}
   );
   gpc615_5 gpc434 (
      {stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413]},
      {stage0_10[302]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[91],stage1_11[117],stage1_10[127],stage1_9[189]}
   );
   gpc615_5 gpc435 (
      {stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418]},
      {stage0_10[303]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[92],stage1_11[118],stage1_10[128],stage1_9[190]}
   );
   gpc615_5 gpc436 (
      {stage0_9[419], stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423]},
      {stage0_10[304]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[93],stage1_11[119],stage1_10[129],stage1_9[191]}
   );
   gpc615_5 gpc437 (
      {stage0_9[424], stage0_9[425], stage0_9[426], stage0_9[427], stage0_9[428]},
      {stage0_10[305]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[94],stage1_11[120],stage1_10[130],stage1_9[192]}
   );
   gpc615_5 gpc438 (
      {stage0_9[429], stage0_9[430], stage0_9[431], stage0_9[432], stage0_9[433]},
      {stage0_10[306]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[95],stage1_11[121],stage1_10[131],stage1_9[193]}
   );
   gpc615_5 gpc439 (
      {stage0_9[434], stage0_9[435], stage0_9[436], stage0_9[437], stage0_9[438]},
      {stage0_10[307]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[96],stage1_11[122],stage1_10[132],stage1_9[194]}
   );
   gpc615_5 gpc440 (
      {stage0_9[439], stage0_9[440], stage0_9[441], stage0_9[442], stage0_9[443]},
      {stage0_10[308]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[97],stage1_11[123],stage1_10[133],stage1_9[195]}
   );
   gpc615_5 gpc441 (
      {stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447], stage0_9[448]},
      {stage0_10[309]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[98],stage1_11[124],stage1_10[134],stage1_9[196]}
   );
   gpc615_5 gpc442 (
      {stage0_9[449], stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453]},
      {stage0_10[310]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[99],stage1_11[125],stage1_10[135],stage1_9[197]}
   );
   gpc615_5 gpc443 (
      {stage0_9[454], stage0_9[455], stage0_9[456], stage0_9[457], stage0_9[458]},
      {stage0_10[311]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[100],stage1_11[126],stage1_10[136],stage1_9[198]}
   );
   gpc615_5 gpc444 (
      {stage0_9[459], stage0_9[460], stage0_9[461], stage0_9[462], stage0_9[463]},
      {stage0_10[312]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[101],stage1_11[127],stage1_10[137],stage1_9[199]}
   );
   gpc615_5 gpc445 (
      {stage0_9[464], stage0_9[465], stage0_9[466], stage0_9[467], stage0_9[468]},
      {stage0_10[313]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[102],stage1_11[128],stage1_10[138],stage1_9[200]}
   );
   gpc615_5 gpc446 (
      {stage0_9[469], stage0_9[470], stage0_9[471], stage0_9[472], stage0_9[473]},
      {stage0_10[314]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[103],stage1_11[129],stage1_10[139],stage1_9[201]}
   );
   gpc615_5 gpc447 (
      {stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477], stage0_9[478]},
      {stage0_10[315]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[104],stage1_11[130],stage1_10[140],stage1_9[202]}
   );
   gpc615_5 gpc448 (
      {stage0_9[479], stage0_9[480], stage0_9[481], stage0_9[482], stage0_9[483]},
      {stage0_10[316]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[105],stage1_11[131],stage1_10[141],stage1_9[203]}
   );
   gpc615_5 gpc449 (
      {stage0_9[484], stage0_9[485], stage0_9[486], stage0_9[487], stage0_9[488]},
      {stage0_10[317]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[106],stage1_11[132],stage1_10[142],stage1_9[204]}
   );
   gpc615_5 gpc450 (
      {stage0_9[489], stage0_9[490], stage0_9[491], stage0_9[492], stage0_9[493]},
      {stage0_10[318]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[107],stage1_11[133],stage1_10[143],stage1_9[205]}
   );
   gpc615_5 gpc451 (
      {stage0_9[494], stage0_9[495], stage0_9[496], stage0_9[497], stage0_9[498]},
      {stage0_10[319]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[108],stage1_11[134],stage1_10[144],stage1_9[206]}
   );
   gpc615_5 gpc452 (
      {stage0_9[499], stage0_9[500], stage0_9[501], stage0_9[502], stage0_9[503]},
      {stage0_10[320]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[109],stage1_11[135],stage1_10[145],stage1_9[207]}
   );
   gpc615_5 gpc453 (
      {stage0_9[504], stage0_9[505], stage0_9[506], stage0_9[507], stage0_9[508]},
      {stage0_10[321]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[110],stage1_11[136],stage1_10[146],stage1_9[208]}
   );
   gpc606_5 gpc454 (
      {stage0_10[322], stage0_10[323], stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[61],stage1_12[111],stage1_11[137],stage1_10[147]}
   );
   gpc606_5 gpc455 (
      {stage0_10[328], stage0_10[329], stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[62],stage1_12[112],stage1_11[138],stage1_10[148]}
   );
   gpc606_5 gpc456 (
      {stage0_10[334], stage0_10[335], stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[63],stage1_12[113],stage1_11[139],stage1_10[149]}
   );
   gpc606_5 gpc457 (
      {stage0_10[340], stage0_10[341], stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[64],stage1_12[114],stage1_11[140],stage1_10[150]}
   );
   gpc606_5 gpc458 (
      {stage0_10[346], stage0_10[347], stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[65],stage1_12[115],stage1_11[141],stage1_10[151]}
   );
   gpc606_5 gpc459 (
      {stage0_10[352], stage0_10[353], stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[66],stage1_12[116],stage1_11[142],stage1_10[152]}
   );
   gpc606_5 gpc460 (
      {stage0_10[358], stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[67],stage1_12[117],stage1_11[143],stage1_10[153]}
   );
   gpc606_5 gpc461 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[68],stage1_12[118],stage1_11[144],stage1_10[154]}
   );
   gpc606_5 gpc462 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[69],stage1_12[119],stage1_11[145],stage1_10[155]}
   );
   gpc606_5 gpc463 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[70],stage1_12[120],stage1_11[146],stage1_10[156]}
   );
   gpc606_5 gpc464 (
      {stage0_10[382], stage0_10[383], stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[71],stage1_12[121],stage1_11[147],stage1_10[157]}
   );
   gpc606_5 gpc465 (
      {stage0_10[388], stage0_10[389], stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[72],stage1_12[122],stage1_11[148],stage1_10[158]}
   );
   gpc606_5 gpc466 (
      {stage0_10[394], stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[73],stage1_12[123],stage1_11[149],stage1_10[159]}
   );
   gpc606_5 gpc467 (
      {stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403], stage0_10[404], stage0_10[405]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[74],stage1_12[124],stage1_11[150],stage1_10[160]}
   );
   gpc606_5 gpc468 (
      {stage0_10[406], stage0_10[407], stage0_10[408], stage0_10[409], stage0_10[410], stage0_10[411]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[75],stage1_12[125],stage1_11[151],stage1_10[161]}
   );
   gpc615_5 gpc469 (
      {stage0_10[412], stage0_10[413], stage0_10[414], stage0_10[415], stage0_10[416]},
      {stage0_11[366]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[76],stage1_12[126],stage1_11[152],stage1_10[162]}
   );
   gpc615_5 gpc470 (
      {stage0_10[417], stage0_10[418], stage0_10[419], stage0_10[420], stage0_10[421]},
      {stage0_11[367]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[77],stage1_12[127],stage1_11[153],stage1_10[163]}
   );
   gpc615_5 gpc471 (
      {stage0_10[422], stage0_10[423], stage0_10[424], stage0_10[425], stage0_10[426]},
      {stage0_11[368]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[78],stage1_12[128],stage1_11[154],stage1_10[164]}
   );
   gpc615_5 gpc472 (
      {stage0_10[427], stage0_10[428], stage0_10[429], stage0_10[430], stage0_10[431]},
      {stage0_11[369]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[79],stage1_12[129],stage1_11[155],stage1_10[165]}
   );
   gpc615_5 gpc473 (
      {stage0_10[432], stage0_10[433], stage0_10[434], stage0_10[435], stage0_10[436]},
      {stage0_11[370]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[80],stage1_12[130],stage1_11[156],stage1_10[166]}
   );
   gpc615_5 gpc474 (
      {stage0_10[437], stage0_10[438], stage0_10[439], stage0_10[440], stage0_10[441]},
      {stage0_11[371]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[81],stage1_12[131],stage1_11[157],stage1_10[167]}
   );
   gpc615_5 gpc475 (
      {stage0_10[442], stage0_10[443], stage0_10[444], stage0_10[445], stage0_10[446]},
      {stage0_11[372]},
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage1_14[21],stage1_13[82],stage1_12[132],stage1_11[158],stage1_10[168]}
   );
   gpc615_5 gpc476 (
      {stage0_10[447], stage0_10[448], stage0_10[449], stage0_10[450], stage0_10[451]},
      {stage0_11[373]},
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage1_14[22],stage1_13[83],stage1_12[133],stage1_11[159],stage1_10[169]}
   );
   gpc615_5 gpc477 (
      {stage0_10[452], stage0_10[453], stage0_10[454], stage0_10[455], stage0_10[456]},
      {stage0_11[374]},
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage1_14[23],stage1_13[84],stage1_12[134],stage1_11[160],stage1_10[170]}
   );
   gpc615_5 gpc478 (
      {stage0_10[457], stage0_10[458], stage0_10[459], stage0_10[460], stage0_10[461]},
      {stage0_11[375]},
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage1_14[24],stage1_13[85],stage1_12[135],stage1_11[161],stage1_10[171]}
   );
   gpc615_5 gpc479 (
      {stage0_10[462], stage0_10[463], stage0_10[464], stage0_10[465], stage0_10[466]},
      {stage0_11[376]},
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage1_14[25],stage1_13[86],stage1_12[136],stage1_11[162],stage1_10[172]}
   );
   gpc615_5 gpc480 (
      {stage0_10[467], stage0_10[468], stage0_10[469], stage0_10[470], stage0_10[471]},
      {stage0_11[377]},
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage1_14[26],stage1_13[87],stage1_12[137],stage1_11[163],stage1_10[173]}
   );
   gpc615_5 gpc481 (
      {stage0_10[472], stage0_10[473], stage0_10[474], stage0_10[475], stage0_10[476]},
      {stage0_11[378]},
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage1_14[27],stage1_13[88],stage1_12[138],stage1_11[164],stage1_10[174]}
   );
   gpc615_5 gpc482 (
      {stage0_10[477], stage0_10[478], stage0_10[479], stage0_10[480], stage0_10[481]},
      {stage0_11[379]},
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage1_14[28],stage1_13[89],stage1_12[139],stage1_11[165],stage1_10[175]}
   );
   gpc615_5 gpc483 (
      {stage0_10[482], stage0_10[483], stage0_10[484], stage0_10[485], stage0_10[486]},
      {stage0_11[380]},
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage1_14[29],stage1_13[90],stage1_12[140],stage1_11[166],stage1_10[176]}
   );
   gpc615_5 gpc484 (
      {stage0_10[487], stage0_10[488], stage0_10[489], stage0_10[490], stage0_10[491]},
      {stage0_11[381]},
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage1_14[30],stage1_13[91],stage1_12[141],stage1_11[167],stage1_10[177]}
   );
   gpc615_5 gpc485 (
      {stage0_10[492], stage0_10[493], stage0_10[494], stage0_10[495], stage0_10[496]},
      {stage0_11[382]},
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage1_14[31],stage1_13[92],stage1_12[142],stage1_11[168],stage1_10[178]}
   );
   gpc615_5 gpc486 (
      {stage0_10[497], stage0_10[498], stage0_10[499], stage0_10[500], stage0_10[501]},
      {stage0_11[383]},
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage1_14[32],stage1_13[93],stage1_12[143],stage1_11[169],stage1_10[179]}
   );
   gpc615_5 gpc487 (
      {stage0_10[502], stage0_10[503], stage0_10[504], stage0_10[505], stage0_10[506]},
      {stage0_11[384]},
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage1_14[33],stage1_13[94],stage1_12[144],stage1_11[170],stage1_10[180]}
   );
   gpc615_5 gpc488 (
      {stage0_10[507], stage0_10[508], stage0_10[509], stage0_10[510], stage0_10[511]},
      {stage0_11[385]},
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage1_14[34],stage1_13[95],stage1_12[145],stage1_11[171],stage1_10[181]}
   );
   gpc615_5 gpc489 (
      {stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389], stage0_11[390]},
      {stage0_12[210]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[35],stage1_13[96],stage1_12[146],stage1_11[172]}
   );
   gpc615_5 gpc490 (
      {stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage0_12[211]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[36],stage1_13[97],stage1_12[147],stage1_11[173]}
   );
   gpc615_5 gpc491 (
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400]},
      {stage0_12[212]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[37],stage1_13[98],stage1_12[148],stage1_11[174]}
   );
   gpc615_5 gpc492 (
      {stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405]},
      {stage0_12[213]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[38],stage1_13[99],stage1_12[149],stage1_11[175]}
   );
   gpc615_5 gpc493 (
      {stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_12[214]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[39],stage1_13[100],stage1_12[150],stage1_11[176]}
   );
   gpc615_5 gpc494 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415]},
      {stage0_12[215]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[40],stage1_13[101],stage1_12[151],stage1_11[177]}
   );
   gpc615_5 gpc495 (
      {stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420]},
      {stage0_12[216]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[41],stage1_13[102],stage1_12[152],stage1_11[178]}
   );
   gpc615_5 gpc496 (
      {stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage0_12[217]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[42],stage1_13[103],stage1_12[153],stage1_11[179]}
   );
   gpc615_5 gpc497 (
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430]},
      {stage0_12[218]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[43],stage1_13[104],stage1_12[154],stage1_11[180]}
   );
   gpc615_5 gpc498 (
      {stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_12[219]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[44],stage1_13[105],stage1_12[155],stage1_11[181]}
   );
   gpc615_5 gpc499 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440]},
      {stage0_12[220]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[45],stage1_13[106],stage1_12[156],stage1_11[182]}
   );
   gpc615_5 gpc500 (
      {stage0_11[441], stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445]},
      {stage0_12[221]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[46],stage1_13[107],stage1_12[157],stage1_11[183]}
   );
   gpc615_5 gpc501 (
      {stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449], stage0_11[450]},
      {stage0_12[222]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[47],stage1_13[108],stage1_12[158],stage1_11[184]}
   );
   gpc615_5 gpc502 (
      {stage0_11[451], stage0_11[452], stage0_11[453], stage0_11[454], stage0_11[455]},
      {stage0_12[223]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[48],stage1_13[109],stage1_12[159],stage1_11[185]}
   );
   gpc615_5 gpc503 (
      {stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459], stage0_11[460]},
      {stage0_12[224]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[49],stage1_13[110],stage1_12[160],stage1_11[186]}
   );
   gpc615_5 gpc504 (
      {stage0_11[461], stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465]},
      {stage0_12[225]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[50],stage1_13[111],stage1_12[161],stage1_11[187]}
   );
   gpc615_5 gpc505 (
      {stage0_11[466], stage0_11[467], stage0_11[468], stage0_11[469], stage0_11[470]},
      {stage0_12[226]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[51],stage1_13[112],stage1_12[162],stage1_11[188]}
   );
   gpc615_5 gpc506 (
      {stage0_11[471], stage0_11[472], stage0_11[473], stage0_11[474], stage0_11[475]},
      {stage0_12[227]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[52],stage1_13[113],stage1_12[163],stage1_11[189]}
   );
   gpc615_5 gpc507 (
      {stage0_11[476], stage0_11[477], stage0_11[478], stage0_11[479], stage0_11[480]},
      {stage0_12[228]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[53],stage1_13[114],stage1_12[164],stage1_11[190]}
   );
   gpc615_5 gpc508 (
      {stage0_11[481], stage0_11[482], stage0_11[483], stage0_11[484], stage0_11[485]},
      {stage0_12[229]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[54],stage1_13[115],stage1_12[165],stage1_11[191]}
   );
   gpc615_5 gpc509 (
      {stage0_11[486], stage0_11[487], stage0_11[488], stage0_11[489], stage0_11[490]},
      {stage0_12[230]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[55],stage1_13[116],stage1_12[166],stage1_11[192]}
   );
   gpc615_5 gpc510 (
      {stage0_11[491], stage0_11[492], stage0_11[493], stage0_11[494], stage0_11[495]},
      {stage0_12[231]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[56],stage1_13[117],stage1_12[167],stage1_11[193]}
   );
   gpc615_5 gpc511 (
      {stage0_11[496], stage0_11[497], stage0_11[498], stage0_11[499], stage0_11[500]},
      {stage0_12[232]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[57],stage1_13[118],stage1_12[168],stage1_11[194]}
   );
   gpc606_5 gpc512 (
      {stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[23],stage1_14[58],stage1_13[119],stage1_12[169]}
   );
   gpc606_5 gpc513 (
      {stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[24],stage1_14[59],stage1_13[120],stage1_12[170]}
   );
   gpc606_5 gpc514 (
      {stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[25],stage1_14[60],stage1_13[121],stage1_12[171]}
   );
   gpc606_5 gpc515 (
      {stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[26],stage1_14[61],stage1_13[122],stage1_12[172]}
   );
   gpc606_5 gpc516 (
      {stage0_12[257], stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[27],stage1_14[62],stage1_13[123],stage1_12[173]}
   );
   gpc606_5 gpc517 (
      {stage0_12[263], stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[28],stage1_14[63],stage1_13[124],stage1_12[174]}
   );
   gpc606_5 gpc518 (
      {stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[29],stage1_14[64],stage1_13[125],stage1_12[175]}
   );
   gpc606_5 gpc519 (
      {stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[30],stage1_14[65],stage1_13[126],stage1_12[176]}
   );
   gpc606_5 gpc520 (
      {stage0_12[281], stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[31],stage1_14[66],stage1_13[127],stage1_12[177]}
   );
   gpc606_5 gpc521 (
      {stage0_12[287], stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[32],stage1_14[67],stage1_13[128],stage1_12[178]}
   );
   gpc606_5 gpc522 (
      {stage0_12[293], stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[33],stage1_14[68],stage1_13[129],stage1_12[179]}
   );
   gpc606_5 gpc523 (
      {stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[34],stage1_14[69],stage1_13[130],stage1_12[180]}
   );
   gpc606_5 gpc524 (
      {stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[35],stage1_14[70],stage1_13[131],stage1_12[181]}
   );
   gpc606_5 gpc525 (
      {stage0_12[311], stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[36],stage1_14[71],stage1_13[132],stage1_12[182]}
   );
   gpc615_5 gpc526 (
      {stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321]},
      {stage0_13[138]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[37],stage1_14[72],stage1_13[133],stage1_12[183]}
   );
   gpc615_5 gpc527 (
      {stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325], stage0_12[326]},
      {stage0_13[139]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[38],stage1_14[73],stage1_13[134],stage1_12[184]}
   );
   gpc615_5 gpc528 (
      {stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330], stage0_12[331]},
      {stage0_13[140]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[39],stage1_14[74],stage1_13[135],stage1_12[185]}
   );
   gpc615_5 gpc529 (
      {stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335], stage0_12[336]},
      {stage0_13[141]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[40],stage1_14[75],stage1_13[136],stage1_12[186]}
   );
   gpc615_5 gpc530 (
      {stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_13[142]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[41],stage1_14[76],stage1_13[137],stage1_12[187]}
   );
   gpc615_5 gpc531 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346]},
      {stage0_13[143]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[42],stage1_14[77],stage1_13[138],stage1_12[188]}
   );
   gpc615_5 gpc532 (
      {stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351]},
      {stage0_13[144]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[43],stage1_14[78],stage1_13[139],stage1_12[189]}
   );
   gpc615_5 gpc533 (
      {stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355], stage0_12[356]},
      {stage0_13[145]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[44],stage1_14[79],stage1_13[140],stage1_12[190]}
   );
   gpc615_5 gpc534 (
      {stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360], stage0_12[361]},
      {stage0_13[146]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[45],stage1_14[80],stage1_13[141],stage1_12[191]}
   );
   gpc615_5 gpc535 (
      {stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365], stage0_12[366]},
      {stage0_13[147]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[46],stage1_14[81],stage1_13[142],stage1_12[192]}
   );
   gpc615_5 gpc536 (
      {stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_13[148]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[47],stage1_14[82],stage1_13[143],stage1_12[193]}
   );
   gpc615_5 gpc537 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376]},
      {stage0_13[149]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[48],stage1_14[83],stage1_13[144],stage1_12[194]}
   );
   gpc615_5 gpc538 (
      {stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381]},
      {stage0_13[150]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[49],stage1_14[84],stage1_13[145],stage1_12[195]}
   );
   gpc615_5 gpc539 (
      {stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385], stage0_12[386]},
      {stage0_13[151]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[50],stage1_14[85],stage1_13[146],stage1_12[196]}
   );
   gpc615_5 gpc540 (
      {stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390], stage0_12[391]},
      {stage0_13[152]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[51],stage1_14[86],stage1_13[147],stage1_12[197]}
   );
   gpc615_5 gpc541 (
      {stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395], stage0_12[396]},
      {stage0_13[153]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[52],stage1_14[87],stage1_13[148],stage1_12[198]}
   );
   gpc615_5 gpc542 (
      {stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_13[154]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[53],stage1_14[88],stage1_13[149],stage1_12[199]}
   );
   gpc615_5 gpc543 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406]},
      {stage0_13[155]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[54],stage1_14[89],stage1_13[150],stage1_12[200]}
   );
   gpc615_5 gpc544 (
      {stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411]},
      {stage0_13[156]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[55],stage1_14[90],stage1_13[151],stage1_12[201]}
   );
   gpc615_5 gpc545 (
      {stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415], stage0_12[416]},
      {stage0_13[157]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[56],stage1_14[91],stage1_13[152],stage1_12[202]}
   );
   gpc615_5 gpc546 (
      {stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420], stage0_12[421]},
      {stage0_13[158]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[57],stage1_14[92],stage1_13[153],stage1_12[203]}
   );
   gpc615_5 gpc547 (
      {stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425], stage0_12[426]},
      {stage0_13[159]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[58],stage1_14[93],stage1_13[154],stage1_12[204]}
   );
   gpc615_5 gpc548 (
      {stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_13[160]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[59],stage1_14[94],stage1_13[155],stage1_12[205]}
   );
   gpc615_5 gpc549 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436]},
      {stage0_13[161]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[60],stage1_14[95],stage1_13[156],stage1_12[206]}
   );
   gpc615_5 gpc550 (
      {stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441]},
      {stage0_13[162]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[61],stage1_14[96],stage1_13[157],stage1_12[207]}
   );
   gpc615_5 gpc551 (
      {stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445], stage0_12[446]},
      {stage0_13[163]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[62],stage1_14[97],stage1_13[158],stage1_12[208]}
   );
   gpc615_5 gpc552 (
      {stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450], stage0_12[451]},
      {stage0_13[164]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[63],stage1_14[98],stage1_13[159],stage1_12[209]}
   );
   gpc615_5 gpc553 (
      {stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455], stage0_12[456]},
      {stage0_13[165]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[64],stage1_14[99],stage1_13[160],stage1_12[210]}
   );
   gpc615_5 gpc554 (
      {stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_13[166]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[65],stage1_14[100],stage1_13[161],stage1_12[211]}
   );
   gpc615_5 gpc555 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466]},
      {stage0_13[167]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[66],stage1_14[101],stage1_13[162],stage1_12[212]}
   );
   gpc615_5 gpc556 (
      {stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471]},
      {stage0_13[168]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[67],stage1_14[102],stage1_13[163],stage1_12[213]}
   );
   gpc615_5 gpc557 (
      {stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475], stage0_12[476]},
      {stage0_13[169]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[68],stage1_14[103],stage1_13[164],stage1_12[214]}
   );
   gpc615_5 gpc558 (
      {stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480], stage0_12[481]},
      {stage0_13[170]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[69],stage1_14[104],stage1_13[165],stage1_12[215]}
   );
   gpc615_5 gpc559 (
      {stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485], stage0_12[486]},
      {stage0_13[171]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[70],stage1_14[105],stage1_13[166],stage1_12[216]}
   );
   gpc615_5 gpc560 (
      {stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_13[172]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[71],stage1_14[106],stage1_13[167],stage1_12[217]}
   );
   gpc615_5 gpc561 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496]},
      {stage0_13[173]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[72],stage1_14[107],stage1_13[168],stage1_12[218]}
   );
   gpc615_5 gpc562 (
      {stage0_12[497], stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501]},
      {stage0_13[174]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[73],stage1_14[108],stage1_13[169],stage1_12[219]}
   );
   gpc615_5 gpc563 (
      {stage0_12[502], stage0_12[503], stage0_12[504], stage0_12[505], stage0_12[506]},
      {stage0_13[175]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[74],stage1_14[109],stage1_13[170],stage1_12[220]}
   );
   gpc615_5 gpc564 (
      {stage0_12[507], stage0_12[508], stage0_12[509], stage0_12[510], stage0_12[511]},
      {stage0_13[176]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[75],stage1_14[110],stage1_13[171],stage1_12[221]}
   );
   gpc606_5 gpc565 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[53],stage1_15[76],stage1_14[111],stage1_13[172]}
   );
   gpc606_5 gpc566 (
      {stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[54],stage1_15[77],stage1_14[112],stage1_13[173]}
   );
   gpc606_5 gpc567 (
      {stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[55],stage1_15[78],stage1_14[113],stage1_13[174]}
   );
   gpc606_5 gpc568 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[56],stage1_15[79],stage1_14[114],stage1_13[175]}
   );
   gpc606_5 gpc569 (
      {stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[57],stage1_15[80],stage1_14[115],stage1_13[176]}
   );
   gpc606_5 gpc570 (
      {stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211], stage0_13[212]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[58],stage1_15[81],stage1_14[116],stage1_13[177]}
   );
   gpc606_5 gpc571 (
      {stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[59],stage1_15[82],stage1_14[117],stage1_13[178]}
   );
   gpc606_5 gpc572 (
      {stage0_13[219], stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[60],stage1_15[83],stage1_14[118],stage1_13[179]}
   );
   gpc606_5 gpc573 (
      {stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[61],stage1_15[84],stage1_14[119],stage1_13[180]}
   );
   gpc606_5 gpc574 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235], stage0_13[236]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[62],stage1_15[85],stage1_14[120],stage1_13[181]}
   );
   gpc606_5 gpc575 (
      {stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241], stage0_13[242]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[63],stage1_15[86],stage1_14[121],stage1_13[182]}
   );
   gpc606_5 gpc576 (
      {stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246], stage0_13[247], stage0_13[248]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[64],stage1_15[87],stage1_14[122],stage1_13[183]}
   );
   gpc606_5 gpc577 (
      {stage0_13[249], stage0_13[250], stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[65],stage1_15[88],stage1_14[123],stage1_13[184]}
   );
   gpc606_5 gpc578 (
      {stage0_13[255], stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[66],stage1_15[89],stage1_14[124],stage1_13[185]}
   );
   gpc606_5 gpc579 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265], stage0_13[266]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[67],stage1_15[90],stage1_14[125],stage1_13[186]}
   );
   gpc606_5 gpc580 (
      {stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270], stage0_13[271], stage0_13[272]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[68],stage1_15[91],stage1_14[126],stage1_13[187]}
   );
   gpc606_5 gpc581 (
      {stage0_13[273], stage0_13[274], stage0_13[275], stage0_13[276], stage0_13[277], stage0_13[278]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[69],stage1_15[92],stage1_14[127],stage1_13[188]}
   );
   gpc606_5 gpc582 (
      {stage0_13[279], stage0_13[280], stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[70],stage1_15[93],stage1_14[128],stage1_13[189]}
   );
   gpc606_5 gpc583 (
      {stage0_13[285], stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[71],stage1_15[94],stage1_14[129],stage1_13[190]}
   );
   gpc606_5 gpc584 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295], stage0_13[296]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[72],stage1_15[95],stage1_14[130],stage1_13[191]}
   );
   gpc606_5 gpc585 (
      {stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300], stage0_13[301], stage0_13[302]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[73],stage1_15[96],stage1_14[131],stage1_13[192]}
   );
   gpc606_5 gpc586 (
      {stage0_13[303], stage0_13[304], stage0_13[305], stage0_13[306], stage0_13[307], stage0_13[308]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[74],stage1_15[97],stage1_14[132],stage1_13[193]}
   );
   gpc606_5 gpc587 (
      {stage0_13[309], stage0_13[310], stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[75],stage1_15[98],stage1_14[133],stage1_13[194]}
   );
   gpc606_5 gpc588 (
      {stage0_13[315], stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[76],stage1_15[99],stage1_14[134],stage1_13[195]}
   );
   gpc606_5 gpc589 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325], stage0_13[326]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[77],stage1_15[100],stage1_14[135],stage1_13[196]}
   );
   gpc606_5 gpc590 (
      {stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330], stage0_13[331], stage0_13[332]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[78],stage1_15[101],stage1_14[136],stage1_13[197]}
   );
   gpc606_5 gpc591 (
      {stage0_13[333], stage0_13[334], stage0_13[335], stage0_13[336], stage0_13[337], stage0_13[338]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[79],stage1_15[102],stage1_14[137],stage1_13[198]}
   );
   gpc606_5 gpc592 (
      {stage0_13[339], stage0_13[340], stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[80],stage1_15[103],stage1_14[138],stage1_13[199]}
   );
   gpc606_5 gpc593 (
      {stage0_13[345], stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[81],stage1_15[104],stage1_14[139],stage1_13[200]}
   );
   gpc606_5 gpc594 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355], stage0_13[356]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[82],stage1_15[105],stage1_14[140],stage1_13[201]}
   );
   gpc606_5 gpc595 (
      {stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360], stage0_13[361], stage0_13[362]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[83],stage1_15[106],stage1_14[141],stage1_13[202]}
   );
   gpc606_5 gpc596 (
      {stage0_13[363], stage0_13[364], stage0_13[365], stage0_13[366], stage0_13[367], stage0_13[368]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[84],stage1_15[107],stage1_14[142],stage1_13[203]}
   );
   gpc606_5 gpc597 (
      {stage0_13[369], stage0_13[370], stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[85],stage1_15[108],stage1_14[143],stage1_13[204]}
   );
   gpc606_5 gpc598 (
      {stage0_13[375], stage0_13[376], stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[86],stage1_15[109],stage1_14[144],stage1_13[205]}
   );
   gpc606_5 gpc599 (
      {stage0_13[381], stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385], stage0_13[386]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[87],stage1_15[110],stage1_14[145],stage1_13[206]}
   );
   gpc606_5 gpc600 (
      {stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390], stage0_13[391], stage0_13[392]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[88],stage1_15[111],stage1_14[146],stage1_13[207]}
   );
   gpc606_5 gpc601 (
      {stage0_13[393], stage0_13[394], stage0_13[395], stage0_13[396], stage0_13[397], stage0_13[398]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[89],stage1_15[112],stage1_14[147],stage1_13[208]}
   );
   gpc606_5 gpc602 (
      {stage0_13[399], stage0_13[400], stage0_13[401], stage0_13[402], stage0_13[403], stage0_13[404]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[90],stage1_15[113],stage1_14[148],stage1_13[209]}
   );
   gpc606_5 gpc603 (
      {stage0_13[405], stage0_13[406], stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[91],stage1_15[114],stage1_14[149],stage1_13[210]}
   );
   gpc606_5 gpc604 (
      {stage0_13[411], stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415], stage0_13[416]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[92],stage1_15[115],stage1_14[150],stage1_13[211]}
   );
   gpc606_5 gpc605 (
      {stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420], stage0_13[421], stage0_13[422]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[93],stage1_15[116],stage1_14[151],stage1_13[212]}
   );
   gpc606_5 gpc606 (
      {stage0_13[423], stage0_13[424], stage0_13[425], stage0_13[426], stage0_13[427], stage0_13[428]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[94],stage1_15[117],stage1_14[152],stage1_13[213]}
   );
   gpc606_5 gpc607 (
      {stage0_13[429], stage0_13[430], stage0_13[431], stage0_13[432], stage0_13[433], stage0_13[434]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[95],stage1_15[118],stage1_14[153],stage1_13[214]}
   );
   gpc606_5 gpc608 (
      {stage0_13[435], stage0_13[436], stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[96],stage1_15[119],stage1_14[154],stage1_13[215]}
   );
   gpc606_5 gpc609 (
      {stage0_13[441], stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445], stage0_13[446]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[97],stage1_15[120],stage1_14[155],stage1_13[216]}
   );
   gpc606_5 gpc610 (
      {stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450], stage0_13[451], stage0_13[452]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[98],stage1_15[121],stage1_14[156],stage1_13[217]}
   );
   gpc606_5 gpc611 (
      {stage0_13[453], stage0_13[454], stage0_13[455], stage0_13[456], stage0_13[457], stage0_13[458]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[99],stage1_15[122],stage1_14[157],stage1_13[218]}
   );
   gpc606_5 gpc612 (
      {stage0_13[459], stage0_13[460], stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[100],stage1_15[123],stage1_14[158],stage1_13[219]}
   );
   gpc606_5 gpc613 (
      {stage0_13[465], stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[101],stage1_15[124],stage1_14[159],stage1_13[220]}
   );
   gpc606_5 gpc614 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475], stage0_13[476]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[102],stage1_15[125],stage1_14[160],stage1_13[221]}
   );
   gpc606_5 gpc615 (
      {stage0_13[477], stage0_13[478], stage0_13[479], stage0_13[480], stage0_13[481], stage0_13[482]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[103],stage1_15[126],stage1_14[161],stage1_13[222]}
   );
   gpc606_5 gpc616 (
      {stage0_13[483], stage0_13[484], stage0_13[485], stage0_13[486], stage0_13[487], stage0_13[488]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[104],stage1_15[127],stage1_14[162],stage1_13[223]}
   );
   gpc606_5 gpc617 (
      {stage0_13[489], stage0_13[490], stage0_13[491], stage0_13[492], stage0_13[493], stage0_13[494]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[105],stage1_15[128],stage1_14[163],stage1_13[224]}
   );
   gpc606_5 gpc618 (
      {stage0_13[495], stage0_13[496], stage0_13[497], stage0_13[498], stage0_13[499], stage0_13[500]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[106],stage1_15[129],stage1_14[164],stage1_13[225]}
   );
   gpc606_5 gpc619 (
      {stage0_13[501], stage0_13[502], stage0_13[503], stage0_13[504], stage0_13[505], stage0_13[506]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[107],stage1_15[130],stage1_14[165],stage1_13[226]}
   );
   gpc606_5 gpc620 (
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[55],stage1_16[108],stage1_15[131],stage1_14[166]}
   );
   gpc606_5 gpc621 (
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[56],stage1_16[109],stage1_15[132],stage1_14[167]}
   );
   gpc606_5 gpc622 (
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[57],stage1_16[110],stage1_15[133],stage1_14[168]}
   );
   gpc606_5 gpc623 (
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[58],stage1_16[111],stage1_15[134],stage1_14[169]}
   );
   gpc606_5 gpc624 (
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[59],stage1_16[112],stage1_15[135],stage1_14[170]}
   );
   gpc606_5 gpc625 (
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[60],stage1_16[113],stage1_15[136],stage1_14[171]}
   );
   gpc606_5 gpc626 (
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[61],stage1_16[114],stage1_15[137],stage1_14[172]}
   );
   gpc606_5 gpc627 (
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[62],stage1_16[115],stage1_15[138],stage1_14[173]}
   );
   gpc606_5 gpc628 (
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[63],stage1_16[116],stage1_15[139],stage1_14[174]}
   );
   gpc606_5 gpc629 (
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[64],stage1_16[117],stage1_15[140],stage1_14[175]}
   );
   gpc606_5 gpc630 (
      {stage0_14[378], stage0_14[379], stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[65],stage1_16[118],stage1_15[141],stage1_14[176]}
   );
   gpc606_5 gpc631 (
      {stage0_14[384], stage0_14[385], stage0_14[386], stage0_14[387], stage0_14[388], stage0_14[389]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[66],stage1_16[119],stage1_15[142],stage1_14[177]}
   );
   gpc606_5 gpc632 (
      {stage0_14[390], stage0_14[391], stage0_14[392], stage0_14[393], stage0_14[394], stage0_14[395]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[67],stage1_16[120],stage1_15[143],stage1_14[178]}
   );
   gpc606_5 gpc633 (
      {stage0_14[396], stage0_14[397], stage0_14[398], stage0_14[399], stage0_14[400], stage0_14[401]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[68],stage1_16[121],stage1_15[144],stage1_14[179]}
   );
   gpc606_5 gpc634 (
      {stage0_14[402], stage0_14[403], stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[69],stage1_16[122],stage1_15[145],stage1_14[180]}
   );
   gpc606_5 gpc635 (
      {stage0_14[408], stage0_14[409], stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[70],stage1_16[123],stage1_15[146],stage1_14[181]}
   );
   gpc606_5 gpc636 (
      {stage0_14[414], stage0_14[415], stage0_14[416], stage0_14[417], stage0_14[418], stage0_14[419]},
      {stage0_16[96], stage0_16[97], stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101]},
      {stage1_18[16],stage1_17[71],stage1_16[124],stage1_15[147],stage1_14[182]}
   );
   gpc606_5 gpc637 (
      {stage0_14[420], stage0_14[421], stage0_14[422], stage0_14[423], stage0_14[424], stage0_14[425]},
      {stage0_16[102], stage0_16[103], stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107]},
      {stage1_18[17],stage1_17[72],stage1_16[125],stage1_15[148],stage1_14[183]}
   );
   gpc606_5 gpc638 (
      {stage0_14[426], stage0_14[427], stage0_14[428], stage0_14[429], stage0_14[430], stage0_14[431]},
      {stage0_16[108], stage0_16[109], stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113]},
      {stage1_18[18],stage1_17[73],stage1_16[126],stage1_15[149],stage1_14[184]}
   );
   gpc606_5 gpc639 (
      {stage0_14[432], stage0_14[433], stage0_14[434], stage0_14[435], stage0_14[436], stage0_14[437]},
      {stage0_16[114], stage0_16[115], stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119]},
      {stage1_18[19],stage1_17[74],stage1_16[127],stage1_15[150],stage1_14[185]}
   );
   gpc606_5 gpc640 (
      {stage0_14[438], stage0_14[439], stage0_14[440], stage0_14[441], stage0_14[442], stage0_14[443]},
      {stage0_16[120], stage0_16[121], stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125]},
      {stage1_18[20],stage1_17[75],stage1_16[128],stage1_15[151],stage1_14[186]}
   );
   gpc606_5 gpc641 (
      {stage0_14[444], stage0_14[445], stage0_14[446], stage0_14[447], stage0_14[448], stage0_14[449]},
      {stage0_16[126], stage0_16[127], stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131]},
      {stage1_18[21],stage1_17[76],stage1_16[129],stage1_15[152],stage1_14[187]}
   );
   gpc606_5 gpc642 (
      {stage0_14[450], stage0_14[451], stage0_14[452], stage0_14[453], stage0_14[454], stage0_14[455]},
      {stage0_16[132], stage0_16[133], stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137]},
      {stage1_18[22],stage1_17[77],stage1_16[130],stage1_15[153],stage1_14[188]}
   );
   gpc606_5 gpc643 (
      {stage0_14[456], stage0_14[457], stage0_14[458], stage0_14[459], stage0_14[460], stage0_14[461]},
      {stage0_16[138], stage0_16[139], stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143]},
      {stage1_18[23],stage1_17[78],stage1_16[131],stage1_15[154],stage1_14[189]}
   );
   gpc615_5 gpc644 (
      {stage0_14[462], stage0_14[463], stage0_14[464], stage0_14[465], stage0_14[466]},
      {stage0_15[330]},
      {stage0_16[144], stage0_16[145], stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149]},
      {stage1_18[24],stage1_17[79],stage1_16[132],stage1_15[155],stage1_14[190]}
   );
   gpc615_5 gpc645 (
      {stage0_14[467], stage0_14[468], stage0_14[469], stage0_14[470], stage0_14[471]},
      {stage0_15[331]},
      {stage0_16[150], stage0_16[151], stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155]},
      {stage1_18[25],stage1_17[80],stage1_16[133],stage1_15[156],stage1_14[191]}
   );
   gpc606_5 gpc646 (
      {stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335], stage0_15[336], stage0_15[337]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[26],stage1_17[81],stage1_16[134],stage1_15[157]}
   );
   gpc606_5 gpc647 (
      {stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341], stage0_15[342], stage0_15[343]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[27],stage1_17[82],stage1_16[135],stage1_15[158]}
   );
   gpc606_5 gpc648 (
      {stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348], stage0_15[349]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[28],stage1_17[83],stage1_16[136],stage1_15[159]}
   );
   gpc606_5 gpc649 (
      {stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353], stage0_15[354], stage0_15[355]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[29],stage1_17[84],stage1_16[137],stage1_15[160]}
   );
   gpc615_5 gpc650 (
      {stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359], stage0_15[360]},
      {stage0_16[156]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[30],stage1_17[85],stage1_16[138],stage1_15[161]}
   );
   gpc615_5 gpc651 (
      {stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage0_16[157]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[31],stage1_17[86],stage1_16[139],stage1_15[162]}
   );
   gpc615_5 gpc652 (
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370]},
      {stage0_16[158]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[32],stage1_17[87],stage1_16[140],stage1_15[163]}
   );
   gpc615_5 gpc653 (
      {stage0_15[371], stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375]},
      {stage0_16[159]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[33],stage1_17[88],stage1_16[141],stage1_15[164]}
   );
   gpc615_5 gpc654 (
      {stage0_15[376], stage0_15[377], stage0_15[378], stage0_15[379], stage0_15[380]},
      {stage0_16[160]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[34],stage1_17[89],stage1_16[142],stage1_15[165]}
   );
   gpc615_5 gpc655 (
      {stage0_15[381], stage0_15[382], stage0_15[383], stage0_15[384], stage0_15[385]},
      {stage0_16[161]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[35],stage1_17[90],stage1_16[143],stage1_15[166]}
   );
   gpc615_5 gpc656 (
      {stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389], stage0_15[390]},
      {stage0_16[162]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[36],stage1_17[91],stage1_16[144],stage1_15[167]}
   );
   gpc615_5 gpc657 (
      {stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395]},
      {stage0_16[163]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[37],stage1_17[92],stage1_16[145],stage1_15[168]}
   );
   gpc615_5 gpc658 (
      {stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400]},
      {stage0_16[164]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[38],stage1_17[93],stage1_16[146],stage1_15[169]}
   );
   gpc615_5 gpc659 (
      {stage0_15[401], stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405]},
      {stage0_16[165]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[39],stage1_17[94],stage1_16[147],stage1_15[170]}
   );
   gpc615_5 gpc660 (
      {stage0_15[406], stage0_15[407], stage0_15[408], stage0_15[409], stage0_15[410]},
      {stage0_16[166]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[40],stage1_17[95],stage1_16[148],stage1_15[171]}
   );
   gpc615_5 gpc661 (
      {stage0_15[411], stage0_15[412], stage0_15[413], stage0_15[414], stage0_15[415]},
      {stage0_16[167]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[41],stage1_17[96],stage1_16[149],stage1_15[172]}
   );
   gpc615_5 gpc662 (
      {stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419], stage0_15[420]},
      {stage0_16[168]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[42],stage1_17[97],stage1_16[150],stage1_15[173]}
   );
   gpc615_5 gpc663 (
      {stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425]},
      {stage0_16[169]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[43],stage1_17[98],stage1_16[151],stage1_15[174]}
   );
   gpc615_5 gpc664 (
      {stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430]},
      {stage0_16[170]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[44],stage1_17[99],stage1_16[152],stage1_15[175]}
   );
   gpc615_5 gpc665 (
      {stage0_15[431], stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435]},
      {stage0_16[171]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[45],stage1_17[100],stage1_16[153],stage1_15[176]}
   );
   gpc615_5 gpc666 (
      {stage0_15[436], stage0_15[437], stage0_15[438], stage0_15[439], stage0_15[440]},
      {stage0_16[172]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[46],stage1_17[101],stage1_16[154],stage1_15[177]}
   );
   gpc615_5 gpc667 (
      {stage0_15[441], stage0_15[442], stage0_15[443], stage0_15[444], stage0_15[445]},
      {stage0_16[173]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[47],stage1_17[102],stage1_16[155],stage1_15[178]}
   );
   gpc615_5 gpc668 (
      {stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449], stage0_15[450]},
      {stage0_16[174]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[48],stage1_17[103],stage1_16[156],stage1_15[179]}
   );
   gpc615_5 gpc669 (
      {stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455]},
      {stage0_16[175]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[49],stage1_17[104],stage1_16[157],stage1_15[180]}
   );
   gpc606_5 gpc670 (
      {stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[24],stage1_18[50],stage1_17[105],stage1_16[158]}
   );
   gpc606_5 gpc671 (
      {stage0_16[182], stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[25],stage1_18[51],stage1_17[106],stage1_16[159]}
   );
   gpc606_5 gpc672 (
      {stage0_16[188], stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[26],stage1_18[52],stage1_17[107],stage1_16[160]}
   );
   gpc606_5 gpc673 (
      {stage0_16[194], stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[27],stage1_18[53],stage1_17[108],stage1_16[161]}
   );
   gpc606_5 gpc674 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[28],stage1_18[54],stage1_17[109],stage1_16[162]}
   );
   gpc606_5 gpc675 (
      {stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[29],stage1_18[55],stage1_17[110],stage1_16[163]}
   );
   gpc606_5 gpc676 (
      {stage0_16[212], stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[30],stage1_18[56],stage1_17[111],stage1_16[164]}
   );
   gpc606_5 gpc677 (
      {stage0_16[218], stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[31],stage1_18[57],stage1_17[112],stage1_16[165]}
   );
   gpc606_5 gpc678 (
      {stage0_16[224], stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[32],stage1_18[58],stage1_17[113],stage1_16[166]}
   );
   gpc606_5 gpc679 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[33],stage1_18[59],stage1_17[114],stage1_16[167]}
   );
   gpc606_5 gpc680 (
      {stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[34],stage1_18[60],stage1_17[115],stage1_16[168]}
   );
   gpc606_5 gpc681 (
      {stage0_16[242], stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[35],stage1_18[61],stage1_17[116],stage1_16[169]}
   );
   gpc606_5 gpc682 (
      {stage0_16[248], stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[36],stage1_18[62],stage1_17[117],stage1_16[170]}
   );
   gpc606_5 gpc683 (
      {stage0_16[254], stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[37],stage1_18[63],stage1_17[118],stage1_16[171]}
   );
   gpc606_5 gpc684 (
      {stage0_16[260], stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[38],stage1_18[64],stage1_17[119],stage1_16[172]}
   );
   gpc606_5 gpc685 (
      {stage0_16[266], stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[39],stage1_18[65],stage1_17[120],stage1_16[173]}
   );
   gpc606_5 gpc686 (
      {stage0_16[272], stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[40],stage1_18[66],stage1_17[121],stage1_16[174]}
   );
   gpc606_5 gpc687 (
      {stage0_16[278], stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[41],stage1_18[67],stage1_17[122],stage1_16[175]}
   );
   gpc606_5 gpc688 (
      {stage0_16[284], stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[42],stage1_18[68],stage1_17[123],stage1_16[176]}
   );
   gpc606_5 gpc689 (
      {stage0_16[290], stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[43],stage1_18[69],stage1_17[124],stage1_16[177]}
   );
   gpc606_5 gpc690 (
      {stage0_16[296], stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[44],stage1_18[70],stage1_17[125],stage1_16[178]}
   );
   gpc606_5 gpc691 (
      {stage0_16[302], stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[45],stage1_18[71],stage1_17[126],stage1_16[179]}
   );
   gpc606_5 gpc692 (
      {stage0_16[308], stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[46],stage1_18[72],stage1_17[127],stage1_16[180]}
   );
   gpc606_5 gpc693 (
      {stage0_16[314], stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[47],stage1_18[73],stage1_17[128],stage1_16[181]}
   );
   gpc606_5 gpc694 (
      {stage0_16[320], stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[48],stage1_18[74],stage1_17[129],stage1_16[182]}
   );
   gpc606_5 gpc695 (
      {stage0_16[326], stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[49],stage1_18[75],stage1_17[130],stage1_16[183]}
   );
   gpc606_5 gpc696 (
      {stage0_16[332], stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[50],stage1_18[76],stage1_17[131],stage1_16[184]}
   );
   gpc606_5 gpc697 (
      {stage0_16[338], stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[51],stage1_18[77],stage1_17[132],stage1_16[185]}
   );
   gpc606_5 gpc698 (
      {stage0_16[344], stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[52],stage1_18[78],stage1_17[133],stage1_16[186]}
   );
   gpc606_5 gpc699 (
      {stage0_16[350], stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[53],stage1_18[79],stage1_17[134],stage1_16[187]}
   );
   gpc606_5 gpc700 (
      {stage0_16[356], stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[54],stage1_18[80],stage1_17[135],stage1_16[188]}
   );
   gpc606_5 gpc701 (
      {stage0_16[362], stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[55],stage1_18[81],stage1_17[136],stage1_16[189]}
   );
   gpc606_5 gpc702 (
      {stage0_16[368], stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[56],stage1_18[82],stage1_17[137],stage1_16[190]}
   );
   gpc606_5 gpc703 (
      {stage0_16[374], stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[57],stage1_18[83],stage1_17[138],stage1_16[191]}
   );
   gpc606_5 gpc704 (
      {stage0_16[380], stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[58],stage1_18[84],stage1_17[139],stage1_16[192]}
   );
   gpc606_5 gpc705 (
      {stage0_16[386], stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[59],stage1_18[85],stage1_17[140],stage1_16[193]}
   );
   gpc606_5 gpc706 (
      {stage0_16[392], stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[60],stage1_18[86],stage1_17[141],stage1_16[194]}
   );
   gpc606_5 gpc707 (
      {stage0_16[398], stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[61],stage1_18[87],stage1_17[142],stage1_16[195]}
   );
   gpc606_5 gpc708 (
      {stage0_16[404], stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[62],stage1_18[88],stage1_17[143],stage1_16[196]}
   );
   gpc606_5 gpc709 (
      {stage0_16[410], stage0_16[411], stage0_16[412], stage0_16[413], stage0_16[414], stage0_16[415]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[63],stage1_18[89],stage1_17[144],stage1_16[197]}
   );
   gpc606_5 gpc710 (
      {stage0_16[416], stage0_16[417], stage0_16[418], stage0_16[419], stage0_16[420], stage0_16[421]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[64],stage1_18[90],stage1_17[145],stage1_16[198]}
   );
   gpc606_5 gpc711 (
      {stage0_16[422], stage0_16[423], stage0_16[424], stage0_16[425], stage0_16[426], stage0_16[427]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[65],stage1_18[91],stage1_17[146],stage1_16[199]}
   );
   gpc606_5 gpc712 (
      {stage0_16[428], stage0_16[429], stage0_16[430], stage0_16[431], stage0_16[432], stage0_16[433]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[66],stage1_18[92],stage1_17[147],stage1_16[200]}
   );
   gpc606_5 gpc713 (
      {stage0_16[434], stage0_16[435], stage0_16[436], stage0_16[437], stage0_16[438], stage0_16[439]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[67],stage1_18[93],stage1_17[148],stage1_16[201]}
   );
   gpc606_5 gpc714 (
      {stage0_16[440], stage0_16[441], stage0_16[442], stage0_16[443], stage0_16[444], stage0_16[445]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[68],stage1_18[94],stage1_17[149],stage1_16[202]}
   );
   gpc606_5 gpc715 (
      {stage0_16[446], stage0_16[447], stage0_16[448], stage0_16[449], stage0_16[450], stage0_16[451]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[69],stage1_18[95],stage1_17[150],stage1_16[203]}
   );
   gpc606_5 gpc716 (
      {stage0_16[452], stage0_16[453], stage0_16[454], stage0_16[455], stage0_16[456], stage0_16[457]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[70],stage1_18[96],stage1_17[151],stage1_16[204]}
   );
   gpc606_5 gpc717 (
      {stage0_16[458], stage0_16[459], stage0_16[460], stage0_16[461], stage0_16[462], stage0_16[463]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[71],stage1_18[97],stage1_17[152],stage1_16[205]}
   );
   gpc606_5 gpc718 (
      {stage0_16[464], stage0_16[465], stage0_16[466], stage0_16[467], stage0_16[468], stage0_16[469]},
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage1_20[48],stage1_19[72],stage1_18[98],stage1_17[153],stage1_16[206]}
   );
   gpc606_5 gpc719 (
      {stage0_16[470], stage0_16[471], stage0_16[472], stage0_16[473], stage0_16[474], stage0_16[475]},
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage1_20[49],stage1_19[73],stage1_18[99],stage1_17[154],stage1_16[207]}
   );
   gpc606_5 gpc720 (
      {stage0_16[476], stage0_16[477], stage0_16[478], stage0_16[479], stage0_16[480], stage0_16[481]},
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage1_20[50],stage1_19[74],stage1_18[100],stage1_17[155],stage1_16[208]}
   );
   gpc606_5 gpc721 (
      {stage0_16[482], stage0_16[483], stage0_16[484], stage0_16[485], stage0_16[486], stage0_16[487]},
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage1_20[51],stage1_19[75],stage1_18[101],stage1_17[156],stage1_16[209]}
   );
   gpc606_5 gpc722 (
      {stage0_16[488], stage0_16[489], stage0_16[490], stage0_16[491], stage0_16[492], stage0_16[493]},
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316], stage0_18[317]},
      {stage1_20[52],stage1_19[76],stage1_18[102],stage1_17[157],stage1_16[210]}
   );
   gpc606_5 gpc723 (
      {stage0_16[494], stage0_16[495], stage0_16[496], stage0_16[497], stage0_16[498], stage0_16[499]},
      {stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321], stage0_18[322], stage0_18[323]},
      {stage1_20[53],stage1_19[77],stage1_18[103],stage1_17[158],stage1_16[211]}
   );
   gpc606_5 gpc724 (
      {stage0_16[500], stage0_16[501], stage0_16[502], stage0_16[503], stage0_16[504], stage0_16[505]},
      {stage0_18[324], stage0_18[325], stage0_18[326], stage0_18[327], stage0_18[328], stage0_18[329]},
      {stage1_20[54],stage1_19[78],stage1_18[104],stage1_17[159],stage1_16[212]}
   );
   gpc606_5 gpc725 (
      {stage0_16[506], stage0_16[507], stage0_16[508], stage0_16[509], stage0_16[510], stage0_16[511]},
      {stage0_18[330], stage0_18[331], stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335]},
      {stage1_20[55],stage1_19[79],stage1_18[105],stage1_17[160],stage1_16[213]}
   );
   gpc606_5 gpc726 (
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[56],stage1_19[80],stage1_18[106],stage1_17[161]}
   );
   gpc606_5 gpc727 (
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[57],stage1_19[81],stage1_18[107],stage1_17[162]}
   );
   gpc606_5 gpc728 (
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[58],stage1_19[82],stage1_18[108],stage1_17[163]}
   );
   gpc606_5 gpc729 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[59],stage1_19[83],stage1_18[109],stage1_17[164]}
   );
   gpc606_5 gpc730 (
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[60],stage1_19[84],stage1_18[110],stage1_17[165]}
   );
   gpc606_5 gpc731 (
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[61],stage1_19[85],stage1_18[111],stage1_17[166]}
   );
   gpc606_5 gpc732 (
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[62],stage1_19[86],stage1_18[112],stage1_17[167]}
   );
   gpc606_5 gpc733 (
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[63],stage1_19[87],stage1_18[113],stage1_17[168]}
   );
   gpc606_5 gpc734 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[64],stage1_19[88],stage1_18[114],stage1_17[169]}
   );
   gpc606_5 gpc735 (
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[65],stage1_19[89],stage1_18[115],stage1_17[170]}
   );
   gpc606_5 gpc736 (
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[66],stage1_19[90],stage1_18[116],stage1_17[171]}
   );
   gpc606_5 gpc737 (
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[67],stage1_19[91],stage1_18[117],stage1_17[172]}
   );
   gpc606_5 gpc738 (
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[68],stage1_19[92],stage1_18[118],stage1_17[173]}
   );
   gpc606_5 gpc739 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[69],stage1_19[93],stage1_18[119],stage1_17[174]}
   );
   gpc606_5 gpc740 (
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[70],stage1_19[94],stage1_18[120],stage1_17[175]}
   );
   gpc606_5 gpc741 (
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[71],stage1_19[95],stage1_18[121],stage1_17[176]}
   );
   gpc606_5 gpc742 (
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[72],stage1_19[96],stage1_18[122],stage1_17[177]}
   );
   gpc606_5 gpc743 (
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[73],stage1_19[97],stage1_18[123],stage1_17[178]}
   );
   gpc606_5 gpc744 (
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[74],stage1_19[98],stage1_18[124],stage1_17[179]}
   );
   gpc606_5 gpc745 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[75],stage1_19[99],stage1_18[125],stage1_17[180]}
   );
   gpc606_5 gpc746 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[76],stage1_19[100],stage1_18[126],stage1_17[181]}
   );
   gpc606_5 gpc747 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[77],stage1_19[101],stage1_18[127],stage1_17[182]}
   );
   gpc606_5 gpc748 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[78],stage1_19[102],stage1_18[128],stage1_17[183]}
   );
   gpc606_5 gpc749 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[79],stage1_19[103],stage1_18[129],stage1_17[184]}
   );
   gpc606_5 gpc750 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[80],stage1_19[104],stage1_18[130],stage1_17[185]}
   );
   gpc606_5 gpc751 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[81],stage1_19[105],stage1_18[131],stage1_17[186]}
   );
   gpc606_5 gpc752 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[82],stage1_19[106],stage1_18[132],stage1_17[187]}
   );
   gpc606_5 gpc753 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[83],stage1_19[107],stage1_18[133],stage1_17[188]}
   );
   gpc606_5 gpc754 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[84],stage1_19[108],stage1_18[134],stage1_17[189]}
   );
   gpc606_5 gpc755 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[85],stage1_19[109],stage1_18[135],stage1_17[190]}
   );
   gpc606_5 gpc756 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[86],stage1_19[110],stage1_18[136],stage1_17[191]}
   );
   gpc606_5 gpc757 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[87],stage1_19[111],stage1_18[137],stage1_17[192]}
   );
   gpc606_5 gpc758 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[88],stage1_19[112],stage1_18[138],stage1_17[193]}
   );
   gpc606_5 gpc759 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[89],stage1_19[113],stage1_18[139],stage1_17[194]}
   );
   gpc606_5 gpc760 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[90],stage1_19[114],stage1_18[140],stage1_17[195]}
   );
   gpc606_5 gpc761 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[91],stage1_19[115],stage1_18[141],stage1_17[196]}
   );
   gpc606_5 gpc762 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[92],stage1_19[116],stage1_18[142],stage1_17[197]}
   );
   gpc606_5 gpc763 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[93],stage1_19[117],stage1_18[143],stage1_17[198]}
   );
   gpc606_5 gpc764 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage1_21[38],stage1_20[94],stage1_19[118],stage1_18[144],stage1_17[199]}
   );
   gpc606_5 gpc765 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage1_21[39],stage1_20[95],stage1_19[119],stage1_18[145],stage1_17[200]}
   );
   gpc606_5 gpc766 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[240], stage0_19[241], stage0_19[242], stage0_19[243], stage0_19[244], stage0_19[245]},
      {stage1_21[40],stage1_20[96],stage1_19[120],stage1_18[146],stage1_17[201]}
   );
   gpc606_5 gpc767 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[246], stage0_19[247], stage0_19[248], stage0_19[249], stage0_19[250], stage0_19[251]},
      {stage1_21[41],stage1_20[97],stage1_19[121],stage1_18[147],stage1_17[202]}
   );
   gpc606_5 gpc768 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[252], stage0_19[253], stage0_19[254], stage0_19[255], stage0_19[256], stage0_19[257]},
      {stage1_21[42],stage1_20[98],stage1_19[122],stage1_18[148],stage1_17[203]}
   );
   gpc606_5 gpc769 (
      {stage0_17[402], stage0_17[403], stage0_17[404], stage0_17[405], stage0_17[406], stage0_17[407]},
      {stage0_19[258], stage0_19[259], stage0_19[260], stage0_19[261], stage0_19[262], stage0_19[263]},
      {stage1_21[43],stage1_20[99],stage1_19[123],stage1_18[149],stage1_17[204]}
   );
   gpc606_5 gpc770 (
      {stage0_17[408], stage0_17[409], stage0_17[410], stage0_17[411], stage0_17[412], stage0_17[413]},
      {stage0_19[264], stage0_19[265], stage0_19[266], stage0_19[267], stage0_19[268], stage0_19[269]},
      {stage1_21[44],stage1_20[100],stage1_19[124],stage1_18[150],stage1_17[205]}
   );
   gpc606_5 gpc771 (
      {stage0_17[414], stage0_17[415], stage0_17[416], stage0_17[417], stage0_17[418], stage0_17[419]},
      {stage0_19[270], stage0_19[271], stage0_19[272], stage0_19[273], stage0_19[274], stage0_19[275]},
      {stage1_21[45],stage1_20[101],stage1_19[125],stage1_18[151],stage1_17[206]}
   );
   gpc606_5 gpc772 (
      {stage0_17[420], stage0_17[421], stage0_17[422], stage0_17[423], stage0_17[424], stage0_17[425]},
      {stage0_19[276], stage0_19[277], stage0_19[278], stage0_19[279], stage0_19[280], stage0_19[281]},
      {stage1_21[46],stage1_20[102],stage1_19[126],stage1_18[152],stage1_17[207]}
   );
   gpc606_5 gpc773 (
      {stage0_17[426], stage0_17[427], stage0_17[428], stage0_17[429], stage0_17[430], stage0_17[431]},
      {stage0_19[282], stage0_19[283], stage0_19[284], stage0_19[285], stage0_19[286], stage0_19[287]},
      {stage1_21[47],stage1_20[103],stage1_19[127],stage1_18[153],stage1_17[208]}
   );
   gpc606_5 gpc774 (
      {stage0_17[432], stage0_17[433], stage0_17[434], stage0_17[435], stage0_17[436], stage0_17[437]},
      {stage0_19[288], stage0_19[289], stage0_19[290], stage0_19[291], stage0_19[292], stage0_19[293]},
      {stage1_21[48],stage1_20[104],stage1_19[128],stage1_18[154],stage1_17[209]}
   );
   gpc606_5 gpc775 (
      {stage0_17[438], stage0_17[439], stage0_17[440], stage0_17[441], stage0_17[442], stage0_17[443]},
      {stage0_19[294], stage0_19[295], stage0_19[296], stage0_19[297], stage0_19[298], stage0_19[299]},
      {stage1_21[49],stage1_20[105],stage1_19[129],stage1_18[155],stage1_17[210]}
   );
   gpc606_5 gpc776 (
      {stage0_17[444], stage0_17[445], stage0_17[446], stage0_17[447], stage0_17[448], stage0_17[449]},
      {stage0_19[300], stage0_19[301], stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305]},
      {stage1_21[50],stage1_20[106],stage1_19[130],stage1_18[156],stage1_17[211]}
   );
   gpc606_5 gpc777 (
      {stage0_17[450], stage0_17[451], stage0_17[452], stage0_17[453], stage0_17[454], stage0_17[455]},
      {stage0_19[306], stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage1_21[51],stage1_20[107],stage1_19[131],stage1_18[157],stage1_17[212]}
   );
   gpc606_5 gpc778 (
      {stage0_17[456], stage0_17[457], stage0_17[458], stage0_17[459], stage0_17[460], stage0_17[461]},
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316], stage0_19[317]},
      {stage1_21[52],stage1_20[108],stage1_19[132],stage1_18[158],stage1_17[213]}
   );
   gpc606_5 gpc779 (
      {stage0_17[462], stage0_17[463], stage0_17[464], stage0_17[465], stage0_17[466], stage0_17[467]},
      {stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321], stage0_19[322], stage0_19[323]},
      {stage1_21[53],stage1_20[109],stage1_19[133],stage1_18[159],stage1_17[214]}
   );
   gpc606_5 gpc780 (
      {stage0_17[468], stage0_17[469], stage0_17[470], stage0_17[471], stage0_17[472], stage0_17[473]},
      {stage0_19[324], stage0_19[325], stage0_19[326], stage0_19[327], stage0_19[328], stage0_19[329]},
      {stage1_21[54],stage1_20[110],stage1_19[134],stage1_18[160],stage1_17[215]}
   );
   gpc606_5 gpc781 (
      {stage0_17[474], stage0_17[475], stage0_17[476], stage0_17[477], stage0_17[478], stage0_17[479]},
      {stage0_19[330], stage0_19[331], stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335]},
      {stage1_21[55],stage1_20[111],stage1_19[135],stage1_18[161],stage1_17[216]}
   );
   gpc606_5 gpc782 (
      {stage0_17[480], stage0_17[481], stage0_17[482], stage0_17[483], stage0_17[484], stage0_17[485]},
      {stage0_19[336], stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage1_21[56],stage1_20[112],stage1_19[136],stage1_18[162],stage1_17[217]}
   );
   gpc606_5 gpc783 (
      {stage0_17[486], stage0_17[487], stage0_17[488], stage0_17[489], stage0_17[490], stage0_17[491]},
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346], stage0_19[347]},
      {stage1_21[57],stage1_20[113],stage1_19[137],stage1_18[163],stage1_17[218]}
   );
   gpc606_5 gpc784 (
      {stage0_17[492], stage0_17[493], stage0_17[494], stage0_17[495], stage0_17[496], stage0_17[497]},
      {stage0_19[348], stage0_19[349], stage0_19[350], stage0_19[351], stage0_19[352], stage0_19[353]},
      {stage1_21[58],stage1_20[114],stage1_19[138],stage1_18[164],stage1_17[219]}
   );
   gpc606_5 gpc785 (
      {stage0_17[498], stage0_17[499], stage0_17[500], stage0_17[501], stage0_17[502], stage0_17[503]},
      {stage0_19[354], stage0_19[355], stage0_19[356], stage0_19[357], stage0_19[358], stage0_19[359]},
      {stage1_21[59],stage1_20[115],stage1_19[139],stage1_18[165],stage1_17[220]}
   );
   gpc606_5 gpc786 (
      {stage0_17[504], stage0_17[505], stage0_17[506], stage0_17[507], stage0_17[508], stage0_17[509]},
      {stage0_19[360], stage0_19[361], stage0_19[362], stage0_19[363], stage0_19[364], stage0_19[365]},
      {stage1_21[60],stage1_20[116],stage1_19[140],stage1_18[166],stage1_17[221]}
   );
   gpc615_5 gpc787 (
      {stage0_18[336], stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340]},
      {stage0_19[366]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[61],stage1_20[117],stage1_19[141],stage1_18[167]}
   );
   gpc615_5 gpc788 (
      {stage0_18[341], stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345]},
      {stage0_19[367]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[62],stage1_20[118],stage1_19[142],stage1_18[168]}
   );
   gpc615_5 gpc789 (
      {stage0_18[346], stage0_18[347], stage0_18[348], stage0_18[349], stage0_18[350]},
      {stage0_19[368]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[63],stage1_20[119],stage1_19[143],stage1_18[169]}
   );
   gpc615_5 gpc790 (
      {stage0_18[351], stage0_18[352], stage0_18[353], stage0_18[354], stage0_18[355]},
      {stage0_19[369]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[64],stage1_20[120],stage1_19[144],stage1_18[170]}
   );
   gpc615_5 gpc791 (
      {stage0_18[356], stage0_18[357], stage0_18[358], stage0_18[359], stage0_18[360]},
      {stage0_19[370]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[65],stage1_20[121],stage1_19[145],stage1_18[171]}
   );
   gpc615_5 gpc792 (
      {stage0_18[361], stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365]},
      {stage0_19[371]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[66],stage1_20[122],stage1_19[146],stage1_18[172]}
   );
   gpc615_5 gpc793 (
      {stage0_18[366], stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370]},
      {stage0_19[372]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[67],stage1_20[123],stage1_19[147],stage1_18[173]}
   );
   gpc615_5 gpc794 (
      {stage0_18[371], stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375]},
      {stage0_19[373]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[68],stage1_20[124],stage1_19[148],stage1_18[174]}
   );
   gpc615_5 gpc795 (
      {stage0_18[376], stage0_18[377], stage0_18[378], stage0_18[379], stage0_18[380]},
      {stage0_19[374]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[69],stage1_20[125],stage1_19[149],stage1_18[175]}
   );
   gpc615_5 gpc796 (
      {stage0_18[381], stage0_18[382], stage0_18[383], stage0_18[384], stage0_18[385]},
      {stage0_19[375]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[70],stage1_20[126],stage1_19[150],stage1_18[176]}
   );
   gpc615_5 gpc797 (
      {stage0_18[386], stage0_18[387], stage0_18[388], stage0_18[389], stage0_18[390]},
      {stage0_19[376]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[71],stage1_20[127],stage1_19[151],stage1_18[177]}
   );
   gpc615_5 gpc798 (
      {stage0_18[391], stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395]},
      {stage0_19[377]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[72],stage1_20[128],stage1_19[152],stage1_18[178]}
   );
   gpc615_5 gpc799 (
      {stage0_18[396], stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400]},
      {stage0_19[378]},
      {stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77]},
      {stage1_22[12],stage1_21[73],stage1_20[129],stage1_19[153],stage1_18[179]}
   );
   gpc615_5 gpc800 (
      {stage0_18[401], stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405]},
      {stage0_19[379]},
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage1_22[13],stage1_21[74],stage1_20[130],stage1_19[154],stage1_18[180]}
   );
   gpc615_5 gpc801 (
      {stage0_18[406], stage0_18[407], stage0_18[408], stage0_18[409], stage0_18[410]},
      {stage0_19[380]},
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage1_22[14],stage1_21[75],stage1_20[131],stage1_19[155],stage1_18[181]}
   );
   gpc615_5 gpc802 (
      {stage0_18[411], stage0_18[412], stage0_18[413], stage0_18[414], stage0_18[415]},
      {stage0_19[381]},
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage1_22[15],stage1_21[76],stage1_20[132],stage1_19[156],stage1_18[182]}
   );
   gpc615_5 gpc803 (
      {stage0_18[416], stage0_18[417], stage0_18[418], stage0_18[419], stage0_18[420]},
      {stage0_19[382]},
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage1_22[16],stage1_21[77],stage1_20[133],stage1_19[157],stage1_18[183]}
   );
   gpc615_5 gpc804 (
      {stage0_18[421], stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425]},
      {stage0_19[383]},
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage1_22[17],stage1_21[78],stage1_20[134],stage1_19[158],stage1_18[184]}
   );
   gpc615_5 gpc805 (
      {stage0_18[426], stage0_18[427], stage0_18[428], stage0_18[429], stage0_18[430]},
      {stage0_19[384]},
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage1_22[18],stage1_21[79],stage1_20[135],stage1_19[159],stage1_18[185]}
   );
   gpc615_5 gpc806 (
      {stage0_18[431], stage0_18[432], stage0_18[433], stage0_18[434], stage0_18[435]},
      {stage0_19[385]},
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage1_22[19],stage1_21[80],stage1_20[136],stage1_19[160],stage1_18[186]}
   );
   gpc615_5 gpc807 (
      {stage0_18[436], stage0_18[437], stage0_18[438], stage0_18[439], stage0_18[440]},
      {stage0_19[386]},
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage1_22[20],stage1_21[81],stage1_20[137],stage1_19[161],stage1_18[187]}
   );
   gpc615_5 gpc808 (
      {stage0_18[441], stage0_18[442], stage0_18[443], stage0_18[444], stage0_18[445]},
      {stage0_19[387]},
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage1_22[21],stage1_21[82],stage1_20[138],stage1_19[162],stage1_18[188]}
   );
   gpc615_5 gpc809 (
      {stage0_18[446], stage0_18[447], stage0_18[448], stage0_18[449], stage0_18[450]},
      {stage0_19[388]},
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage1_22[22],stage1_21[83],stage1_20[139],stage1_19[163],stage1_18[189]}
   );
   gpc615_5 gpc810 (
      {stage0_18[451], stage0_18[452], stage0_18[453], stage0_18[454], stage0_18[455]},
      {stage0_19[389]},
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage1_22[23],stage1_21[84],stage1_20[140],stage1_19[164],stage1_18[190]}
   );
   gpc615_5 gpc811 (
      {stage0_18[456], stage0_18[457], stage0_18[458], stage0_18[459], stage0_18[460]},
      {stage0_19[390]},
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage1_22[24],stage1_21[85],stage1_20[141],stage1_19[165],stage1_18[191]}
   );
   gpc615_5 gpc812 (
      {stage0_18[461], stage0_18[462], stage0_18[463], stage0_18[464], stage0_18[465]},
      {stage0_19[391]},
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage1_22[25],stage1_21[86],stage1_20[142],stage1_19[166],stage1_18[192]}
   );
   gpc615_5 gpc813 (
      {stage0_18[466], stage0_18[467], stage0_18[468], stage0_18[469], stage0_18[470]},
      {stage0_19[392]},
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage1_22[26],stage1_21[87],stage1_20[143],stage1_19[167],stage1_18[193]}
   );
   gpc615_5 gpc814 (
      {stage0_18[471], stage0_18[472], stage0_18[473], stage0_18[474], stage0_18[475]},
      {stage0_19[393]},
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage1_22[27],stage1_21[88],stage1_20[144],stage1_19[168],stage1_18[194]}
   );
   gpc615_5 gpc815 (
      {stage0_18[476], stage0_18[477], stage0_18[478], stage0_18[479], stage0_18[480]},
      {stage0_19[394]},
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage1_22[28],stage1_21[89],stage1_20[145],stage1_19[169],stage1_18[195]}
   );
   gpc615_5 gpc816 (
      {stage0_18[481], stage0_18[482], stage0_18[483], stage0_18[484], stage0_18[485]},
      {stage0_19[395]},
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage1_22[29],stage1_21[90],stage1_20[146],stage1_19[170],stage1_18[196]}
   );
   gpc615_5 gpc817 (
      {stage0_18[486], stage0_18[487], stage0_18[488], stage0_18[489], stage0_18[490]},
      {stage0_19[396]},
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage1_22[30],stage1_21[91],stage1_20[147],stage1_19[171],stage1_18[197]}
   );
   gpc615_5 gpc818 (
      {stage0_18[491], stage0_18[492], stage0_18[493], stage0_18[494], stage0_18[495]},
      {stage0_19[397]},
      {stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190], stage0_20[191]},
      {stage1_22[31],stage1_21[92],stage1_20[148],stage1_19[172],stage1_18[198]}
   );
   gpc615_5 gpc819 (
      {stage0_18[496], stage0_18[497], stage0_18[498], stage0_18[499], stage0_18[500]},
      {stage0_19[398]},
      {stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196], stage0_20[197]},
      {stage1_22[32],stage1_21[93],stage1_20[149],stage1_19[173],stage1_18[199]}
   );
   gpc615_5 gpc820 (
      {stage0_18[501], stage0_18[502], stage0_18[503], stage0_18[504], stage0_18[505]},
      {stage0_19[399]},
      {stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202], stage0_20[203]},
      {stage1_22[33],stage1_21[94],stage1_20[150],stage1_19[174],stage1_18[200]}
   );
   gpc615_5 gpc821 (
      {stage0_18[506], stage0_18[507], stage0_18[508], stage0_18[509], stage0_18[510]},
      {stage0_19[400]},
      {stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208], stage0_20[209]},
      {stage1_22[34],stage1_21[95],stage1_20[151],stage1_19[175],stage1_18[201]}
   );
   gpc615_5 gpc822 (
      {stage0_19[401], stage0_19[402], stage0_19[403], stage0_19[404], stage0_19[405]},
      {stage0_20[210]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[35],stage1_21[96],stage1_20[152],stage1_19[176]}
   );
   gpc615_5 gpc823 (
      {stage0_19[406], stage0_19[407], stage0_19[408], stage0_19[409], stage0_19[410]},
      {stage0_20[211]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[36],stage1_21[97],stage1_20[153],stage1_19[177]}
   );
   gpc615_5 gpc824 (
      {stage0_19[411], stage0_19[412], stage0_19[413], stage0_19[414], stage0_19[415]},
      {stage0_20[212]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[37],stage1_21[98],stage1_20[154],stage1_19[178]}
   );
   gpc615_5 gpc825 (
      {stage0_19[416], stage0_19[417], stage0_19[418], stage0_19[419], stage0_19[420]},
      {stage0_20[213]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[38],stage1_21[99],stage1_20[155],stage1_19[179]}
   );
   gpc615_5 gpc826 (
      {stage0_19[421], stage0_19[422], stage0_19[423], stage0_19[424], stage0_19[425]},
      {stage0_20[214]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[39],stage1_21[100],stage1_20[156],stage1_19[180]}
   );
   gpc615_5 gpc827 (
      {stage0_19[426], stage0_19[427], stage0_19[428], stage0_19[429], stage0_19[430]},
      {stage0_20[215]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[40],stage1_21[101],stage1_20[157],stage1_19[181]}
   );
   gpc606_5 gpc828 (
      {stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220], stage0_20[221]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[6],stage1_22[41],stage1_21[102],stage1_20[158]}
   );
   gpc606_5 gpc829 (
      {stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226], stage0_20[227]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[7],stage1_22[42],stage1_21[103],stage1_20[159]}
   );
   gpc606_5 gpc830 (
      {stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232], stage0_20[233]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[8],stage1_22[43],stage1_21[104],stage1_20[160]}
   );
   gpc606_5 gpc831 (
      {stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238], stage0_20[239]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[9],stage1_22[44],stage1_21[105],stage1_20[161]}
   );
   gpc606_5 gpc832 (
      {stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244], stage0_20[245]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[10],stage1_22[45],stage1_21[106],stage1_20[162]}
   );
   gpc606_5 gpc833 (
      {stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249], stage0_20[250], stage0_20[251]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[11],stage1_22[46],stage1_21[107],stage1_20[163]}
   );
   gpc606_5 gpc834 (
      {stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255], stage0_20[256], stage0_20[257]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[12],stage1_22[47],stage1_21[108],stage1_20[164]}
   );
   gpc606_5 gpc835 (
      {stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261], stage0_20[262], stage0_20[263]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[13],stage1_22[48],stage1_21[109],stage1_20[165]}
   );
   gpc606_5 gpc836 (
      {stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267], stage0_20[268], stage0_20[269]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[14],stage1_22[49],stage1_21[110],stage1_20[166]}
   );
   gpc606_5 gpc837 (
      {stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273], stage0_20[274], stage0_20[275]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[15],stage1_22[50],stage1_21[111],stage1_20[167]}
   );
   gpc606_5 gpc838 (
      {stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279], stage0_20[280], stage0_20[281]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[16],stage1_22[51],stage1_21[112],stage1_20[168]}
   );
   gpc606_5 gpc839 (
      {stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285], stage0_20[286], stage0_20[287]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[17],stage1_22[52],stage1_21[113],stage1_20[169]}
   );
   gpc606_5 gpc840 (
      {stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291], stage0_20[292], stage0_20[293]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[18],stage1_22[53],stage1_21[114],stage1_20[170]}
   );
   gpc606_5 gpc841 (
      {stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297], stage0_20[298], stage0_20[299]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[19],stage1_22[54],stage1_21[115],stage1_20[171]}
   );
   gpc606_5 gpc842 (
      {stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303], stage0_20[304], stage0_20[305]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[20],stage1_22[55],stage1_21[116],stage1_20[172]}
   );
   gpc606_5 gpc843 (
      {stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309], stage0_20[310], stage0_20[311]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[21],stage1_22[56],stage1_21[117],stage1_20[173]}
   );
   gpc606_5 gpc844 (
      {stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315], stage0_20[316], stage0_20[317]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[22],stage1_22[57],stage1_21[118],stage1_20[174]}
   );
   gpc606_5 gpc845 (
      {stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321], stage0_20[322], stage0_20[323]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[23],stage1_22[58],stage1_21[119],stage1_20[175]}
   );
   gpc606_5 gpc846 (
      {stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327], stage0_20[328], stage0_20[329]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[24],stage1_22[59],stage1_21[120],stage1_20[176]}
   );
   gpc606_5 gpc847 (
      {stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333], stage0_20[334], stage0_20[335]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[25],stage1_22[60],stage1_21[121],stage1_20[177]}
   );
   gpc606_5 gpc848 (
      {stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339], stage0_20[340], stage0_20[341]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[26],stage1_22[61],stage1_21[122],stage1_20[178]}
   );
   gpc606_5 gpc849 (
      {stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345], stage0_20[346], stage0_20[347]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[27],stage1_22[62],stage1_21[123],stage1_20[179]}
   );
   gpc606_5 gpc850 (
      {stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351], stage0_20[352], stage0_20[353]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[28],stage1_22[63],stage1_21[124],stage1_20[180]}
   );
   gpc606_5 gpc851 (
      {stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357], stage0_20[358], stage0_20[359]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[29],stage1_22[64],stage1_21[125],stage1_20[181]}
   );
   gpc606_5 gpc852 (
      {stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363], stage0_20[364], stage0_20[365]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[30],stage1_22[65],stage1_21[126],stage1_20[182]}
   );
   gpc606_5 gpc853 (
      {stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369], stage0_20[370], stage0_20[371]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[31],stage1_22[66],stage1_21[127],stage1_20[183]}
   );
   gpc606_5 gpc854 (
      {stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375], stage0_20[376], stage0_20[377]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[32],stage1_22[67],stage1_21[128],stage1_20[184]}
   );
   gpc606_5 gpc855 (
      {stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381], stage0_20[382], stage0_20[383]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[33],stage1_22[68],stage1_21[129],stage1_20[185]}
   );
   gpc606_5 gpc856 (
      {stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387], stage0_20[388], stage0_20[389]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[34],stage1_22[69],stage1_21[130],stage1_20[186]}
   );
   gpc606_5 gpc857 (
      {stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393], stage0_20[394], stage0_20[395]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[35],stage1_22[70],stage1_21[131],stage1_20[187]}
   );
   gpc606_5 gpc858 (
      {stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399], stage0_20[400], stage0_20[401]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[36],stage1_22[71],stage1_21[132],stage1_20[188]}
   );
   gpc606_5 gpc859 (
      {stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405], stage0_20[406], stage0_20[407]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[37],stage1_22[72],stage1_21[133],stage1_20[189]}
   );
   gpc606_5 gpc860 (
      {stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411], stage0_20[412], stage0_20[413]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[38],stage1_22[73],stage1_21[134],stage1_20[190]}
   );
   gpc606_5 gpc861 (
      {stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417], stage0_20[418], stage0_20[419]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[39],stage1_22[74],stage1_21[135],stage1_20[191]}
   );
   gpc606_5 gpc862 (
      {stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423], stage0_20[424], stage0_20[425]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[40],stage1_22[75],stage1_21[136],stage1_20[192]}
   );
   gpc606_5 gpc863 (
      {stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429], stage0_20[430], stage0_20[431]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[41],stage1_22[76],stage1_21[137],stage1_20[193]}
   );
   gpc606_5 gpc864 (
      {stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435], stage0_20[436], stage0_20[437]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[42],stage1_22[77],stage1_21[138],stage1_20[194]}
   );
   gpc606_5 gpc865 (
      {stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441], stage0_20[442], stage0_20[443]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[43],stage1_22[78],stage1_21[139],stage1_20[195]}
   );
   gpc606_5 gpc866 (
      {stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447], stage0_20[448], stage0_20[449]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[44],stage1_22[79],stage1_21[140],stage1_20[196]}
   );
   gpc606_5 gpc867 (
      {stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453], stage0_20[454], stage0_20[455]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[45],stage1_22[80],stage1_21[141],stage1_20[197]}
   );
   gpc606_5 gpc868 (
      {stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459], stage0_20[460], stage0_20[461]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[46],stage1_22[81],stage1_21[142],stage1_20[198]}
   );
   gpc606_5 gpc869 (
      {stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465], stage0_20[466], stage0_20[467]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[47],stage1_22[82],stage1_21[143],stage1_20[199]}
   );
   gpc606_5 gpc870 (
      {stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471], stage0_20[472], stage0_20[473]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[48],stage1_22[83],stage1_21[144],stage1_20[200]}
   );
   gpc606_5 gpc871 (
      {stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477], stage0_20[478], stage0_20[479]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[49],stage1_22[84],stage1_21[145],stage1_20[201]}
   );
   gpc606_5 gpc872 (
      {stage0_20[480], stage0_20[481], stage0_20[482], stage0_20[483], stage0_20[484], stage0_20[485]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[50],stage1_22[85],stage1_21[146],stage1_20[202]}
   );
   gpc606_5 gpc873 (
      {stage0_20[486], stage0_20[487], stage0_20[488], stage0_20[489], stage0_20[490], stage0_20[491]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[51],stage1_22[86],stage1_21[147],stage1_20[203]}
   );
   gpc606_5 gpc874 (
      {stage0_20[492], stage0_20[493], stage0_20[494], stage0_20[495], stage0_20[496], stage0_20[497]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[52],stage1_22[87],stage1_21[148],stage1_20[204]}
   );
   gpc606_5 gpc875 (
      {stage0_20[498], stage0_20[499], stage0_20[500], stage0_20[501], stage0_20[502], stage0_20[503]},
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286], stage0_22[287]},
      {stage1_24[47],stage1_23[53],stage1_22[88],stage1_21[149],stage1_20[205]}
   );
   gpc606_5 gpc876 (
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[48],stage1_23[54],stage1_22[89],stage1_21[150]}
   );
   gpc606_5 gpc877 (
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[49],stage1_23[55],stage1_22[90],stage1_21[151]}
   );
   gpc606_5 gpc878 (
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[50],stage1_23[56],stage1_22[91],stage1_21[152]}
   );
   gpc606_5 gpc879 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[51],stage1_23[57],stage1_22[92],stage1_21[153]}
   );
   gpc606_5 gpc880 (
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[52],stage1_23[58],stage1_22[93],stage1_21[154]}
   );
   gpc606_5 gpc881 (
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[53],stage1_23[59],stage1_22[94],stage1_21[155]}
   );
   gpc606_5 gpc882 (
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[54],stage1_23[60],stage1_22[95],stage1_21[156]}
   );
   gpc606_5 gpc883 (
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[55],stage1_23[61],stage1_22[96],stage1_21[157]}
   );
   gpc606_5 gpc884 (
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[56],stage1_23[62],stage1_22[97],stage1_21[158]}
   );
   gpc606_5 gpc885 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[57],stage1_23[63],stage1_22[98],stage1_21[159]}
   );
   gpc606_5 gpc886 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[58],stage1_23[64],stage1_22[99],stage1_21[160]}
   );
   gpc606_5 gpc887 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[59],stage1_23[65],stage1_22[100],stage1_21[161]}
   );
   gpc606_5 gpc888 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[60],stage1_23[66],stage1_22[101],stage1_21[162]}
   );
   gpc606_5 gpc889 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[61],stage1_23[67],stage1_22[102],stage1_21[163]}
   );
   gpc606_5 gpc890 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[62],stage1_23[68],stage1_22[103],stage1_21[164]}
   );
   gpc606_5 gpc891 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[63],stage1_23[69],stage1_22[104],stage1_21[165]}
   );
   gpc606_5 gpc892 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[64],stage1_23[70],stage1_22[105],stage1_21[166]}
   );
   gpc606_5 gpc893 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[65],stage1_23[71],stage1_22[106],stage1_21[167]}
   );
   gpc606_5 gpc894 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[66],stage1_23[72],stage1_22[107],stage1_21[168]}
   );
   gpc606_5 gpc895 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[67],stage1_23[73],stage1_22[108],stage1_21[169]}
   );
   gpc606_5 gpc896 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[68],stage1_23[74],stage1_22[109],stage1_21[170]}
   );
   gpc606_5 gpc897 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[69],stage1_23[75],stage1_22[110],stage1_21[171]}
   );
   gpc606_5 gpc898 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[70],stage1_23[76],stage1_22[111],stage1_21[172]}
   );
   gpc606_5 gpc899 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[71],stage1_23[77],stage1_22[112],stage1_21[173]}
   );
   gpc606_5 gpc900 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[72],stage1_23[78],stage1_22[113],stage1_21[174]}
   );
   gpc606_5 gpc901 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[73],stage1_23[79],stage1_22[114],stage1_21[175]}
   );
   gpc606_5 gpc902 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[74],stage1_23[80],stage1_22[115],stage1_21[176]}
   );
   gpc606_5 gpc903 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[75],stage1_23[81],stage1_22[116],stage1_21[177]}
   );
   gpc606_5 gpc904 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[76],stage1_23[82],stage1_22[117],stage1_21[178]}
   );
   gpc606_5 gpc905 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[77],stage1_23[83],stage1_22[118],stage1_21[179]}
   );
   gpc606_5 gpc906 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[78],stage1_23[84],stage1_22[119],stage1_21[180]}
   );
   gpc606_5 gpc907 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage1_25[31],stage1_24[79],stage1_23[85],stage1_22[120],stage1_21[181]}
   );
   gpc606_5 gpc908 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage1_25[32],stage1_24[80],stage1_23[86],stage1_22[121],stage1_21[182]}
   );
   gpc606_5 gpc909 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage1_25[33],stage1_24[81],stage1_23[87],stage1_22[122],stage1_21[183]}
   );
   gpc606_5 gpc910 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage1_25[34],stage1_24[82],stage1_23[88],stage1_22[123],stage1_21[184]}
   );
   gpc606_5 gpc911 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage1_25[35],stage1_24[83],stage1_23[89],stage1_22[124],stage1_21[185]}
   );
   gpc606_5 gpc912 (
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage1_25[36],stage1_24[84],stage1_23[90],stage1_22[125],stage1_21[186]}
   );
   gpc606_5 gpc913 (
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage1_25[37],stage1_24[85],stage1_23[91],stage1_22[126],stage1_21[187]}
   );
   gpc606_5 gpc914 (
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage1_25[38],stage1_24[86],stage1_23[92],stage1_22[127],stage1_21[188]}
   );
   gpc606_5 gpc915 (
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage1_25[39],stage1_24[87],stage1_23[93],stage1_22[128],stage1_21[189]}
   );
   gpc615_5 gpc916 (
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280]},
      {stage0_22[288]},
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage1_25[40],stage1_24[88],stage1_23[94],stage1_22[129],stage1_21[190]}
   );
   gpc615_5 gpc917 (
      {stage0_21[281], stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285]},
      {stage0_22[289]},
      {stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251]},
      {stage1_25[41],stage1_24[89],stage1_23[95],stage1_22[130],stage1_21[191]}
   );
   gpc615_5 gpc918 (
      {stage0_21[286], stage0_21[287], stage0_21[288], stage0_21[289], stage0_21[290]},
      {stage0_22[290]},
      {stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage1_25[42],stage1_24[90],stage1_23[96],stage1_22[131],stage1_21[192]}
   );
   gpc615_5 gpc919 (
      {stage0_21[291], stage0_21[292], stage0_21[293], stage0_21[294], stage0_21[295]},
      {stage0_22[291]},
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262], stage0_23[263]},
      {stage1_25[43],stage1_24[91],stage1_23[97],stage1_22[132],stage1_21[193]}
   );
   gpc615_5 gpc920 (
      {stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299], stage0_21[300]},
      {stage0_22[292]},
      {stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268], stage0_23[269]},
      {stage1_25[44],stage1_24[92],stage1_23[98],stage1_22[133],stage1_21[194]}
   );
   gpc615_5 gpc921 (
      {stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_22[293]},
      {stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274], stage0_23[275]},
      {stage1_25[45],stage1_24[93],stage1_23[99],stage1_22[134],stage1_21[195]}
   );
   gpc615_5 gpc922 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310]},
      {stage0_22[294]},
      {stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281]},
      {stage1_25[46],stage1_24[94],stage1_23[100],stage1_22[135],stage1_21[196]}
   );
   gpc615_5 gpc923 (
      {stage0_21[311], stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315]},
      {stage0_22[295]},
      {stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage1_25[47],stage1_24[95],stage1_23[101],stage1_22[136],stage1_21[197]}
   );
   gpc615_5 gpc924 (
      {stage0_21[316], stage0_21[317], stage0_21[318], stage0_21[319], stage0_21[320]},
      {stage0_22[296]},
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292], stage0_23[293]},
      {stage1_25[48],stage1_24[96],stage1_23[102],stage1_22[137],stage1_21[198]}
   );
   gpc615_5 gpc925 (
      {stage0_21[321], stage0_21[322], stage0_21[323], stage0_21[324], stage0_21[325]},
      {stage0_22[297]},
      {stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298], stage0_23[299]},
      {stage1_25[49],stage1_24[97],stage1_23[103],stage1_22[138],stage1_21[199]}
   );
   gpc615_5 gpc926 (
      {stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329], stage0_21[330]},
      {stage0_22[298]},
      {stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304], stage0_23[305]},
      {stage1_25[50],stage1_24[98],stage1_23[104],stage1_22[139],stage1_21[200]}
   );
   gpc615_5 gpc927 (
      {stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_22[299]},
      {stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311]},
      {stage1_25[51],stage1_24[99],stage1_23[105],stage1_22[140],stage1_21[201]}
   );
   gpc615_5 gpc928 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340]},
      {stage0_22[300]},
      {stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage1_25[52],stage1_24[100],stage1_23[106],stage1_22[141],stage1_21[202]}
   );
   gpc615_5 gpc929 (
      {stage0_21[341], stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345]},
      {stage0_22[301]},
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322], stage0_23[323]},
      {stage1_25[53],stage1_24[101],stage1_23[107],stage1_22[142],stage1_21[203]}
   );
   gpc615_5 gpc930 (
      {stage0_21[346], stage0_21[347], stage0_21[348], stage0_21[349], stage0_21[350]},
      {stage0_22[302]},
      {stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328], stage0_23[329]},
      {stage1_25[54],stage1_24[102],stage1_23[108],stage1_22[143],stage1_21[204]}
   );
   gpc615_5 gpc931 (
      {stage0_21[351], stage0_21[352], stage0_21[353], stage0_21[354], stage0_21[355]},
      {stage0_22[303]},
      {stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334], stage0_23[335]},
      {stage1_25[55],stage1_24[103],stage1_23[109],stage1_22[144],stage1_21[205]}
   );
   gpc615_5 gpc932 (
      {stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359], stage0_21[360]},
      {stage0_22[304]},
      {stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341]},
      {stage1_25[56],stage1_24[104],stage1_23[110],stage1_22[145],stage1_21[206]}
   );
   gpc615_5 gpc933 (
      {stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_22[305]},
      {stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage1_25[57],stage1_24[105],stage1_23[111],stage1_22[146],stage1_21[207]}
   );
   gpc615_5 gpc934 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370]},
      {stage0_22[306]},
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352], stage0_23[353]},
      {stage1_25[58],stage1_24[106],stage1_23[112],stage1_22[147],stage1_21[208]}
   );
   gpc615_5 gpc935 (
      {stage0_21[371], stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375]},
      {stage0_22[307]},
      {stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358], stage0_23[359]},
      {stage1_25[59],stage1_24[107],stage1_23[113],stage1_22[148],stage1_21[209]}
   );
   gpc615_5 gpc936 (
      {stage0_21[376], stage0_21[377], stage0_21[378], stage0_21[379], stage0_21[380]},
      {stage0_22[308]},
      {stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364], stage0_23[365]},
      {stage1_25[60],stage1_24[108],stage1_23[114],stage1_22[149],stage1_21[210]}
   );
   gpc615_5 gpc937 (
      {stage0_21[381], stage0_21[382], stage0_21[383], stage0_21[384], stage0_21[385]},
      {stage0_22[309]},
      {stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371]},
      {stage1_25[61],stage1_24[109],stage1_23[115],stage1_22[150],stage1_21[211]}
   );
   gpc615_5 gpc938 (
      {stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389], stage0_21[390]},
      {stage0_22[310]},
      {stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage1_25[62],stage1_24[110],stage1_23[116],stage1_22[151],stage1_21[212]}
   );
   gpc615_5 gpc939 (
      {stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_22[311]},
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382], stage0_23[383]},
      {stage1_25[63],stage1_24[111],stage1_23[117],stage1_22[152],stage1_21[213]}
   );
   gpc615_5 gpc940 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400]},
      {stage0_22[312]},
      {stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387], stage0_23[388], stage0_23[389]},
      {stage1_25[64],stage1_24[112],stage1_23[118],stage1_22[153],stage1_21[214]}
   );
   gpc615_5 gpc941 (
      {stage0_21[401], stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405]},
      {stage0_22[313]},
      {stage0_23[390], stage0_23[391], stage0_23[392], stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage1_25[65],stage1_24[113],stage1_23[119],stage1_22[154],stage1_21[215]}
   );
   gpc615_5 gpc942 (
      {stage0_21[406], stage0_21[407], stage0_21[408], stage0_21[409], stage0_21[410]},
      {stage0_22[314]},
      {stage0_23[396], stage0_23[397], stage0_23[398], stage0_23[399], stage0_23[400], stage0_23[401]},
      {stage1_25[66],stage1_24[114],stage1_23[120],stage1_22[155],stage1_21[216]}
   );
   gpc615_5 gpc943 (
      {stage0_21[411], stage0_21[412], stage0_21[413], stage0_21[414], stage0_21[415]},
      {stage0_22[315]},
      {stage0_23[402], stage0_23[403], stage0_23[404], stage0_23[405], stage0_23[406], stage0_23[407]},
      {stage1_25[67],stage1_24[115],stage1_23[121],stage1_22[156],stage1_21[217]}
   );
   gpc615_5 gpc944 (
      {stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419], stage0_21[420]},
      {stage0_22[316]},
      {stage0_23[408], stage0_23[409], stage0_23[410], stage0_23[411], stage0_23[412], stage0_23[413]},
      {stage1_25[68],stage1_24[116],stage1_23[122],stage1_22[157],stage1_21[218]}
   );
   gpc615_5 gpc945 (
      {stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_22[317]},
      {stage0_23[414], stage0_23[415], stage0_23[416], stage0_23[417], stage0_23[418], stage0_23[419]},
      {stage1_25[69],stage1_24[117],stage1_23[123],stage1_22[158],stage1_21[219]}
   );
   gpc615_5 gpc946 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430]},
      {stage0_22[318]},
      {stage0_23[420], stage0_23[421], stage0_23[422], stage0_23[423], stage0_23[424], stage0_23[425]},
      {stage1_25[70],stage1_24[118],stage1_23[124],stage1_22[159],stage1_21[220]}
   );
   gpc615_5 gpc947 (
      {stage0_21[431], stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435]},
      {stage0_22[319]},
      {stage0_23[426], stage0_23[427], stage0_23[428], stage0_23[429], stage0_23[430], stage0_23[431]},
      {stage1_25[71],stage1_24[119],stage1_23[125],stage1_22[160],stage1_21[221]}
   );
   gpc615_5 gpc948 (
      {stage0_21[436], stage0_21[437], stage0_21[438], stage0_21[439], stage0_21[440]},
      {stage0_22[320]},
      {stage0_23[432], stage0_23[433], stage0_23[434], stage0_23[435], stage0_23[436], stage0_23[437]},
      {stage1_25[72],stage1_24[120],stage1_23[126],stage1_22[161],stage1_21[222]}
   );
   gpc615_5 gpc949 (
      {stage0_21[441], stage0_21[442], stage0_21[443], stage0_21[444], stage0_21[445]},
      {stage0_22[321]},
      {stage0_23[438], stage0_23[439], stage0_23[440], stage0_23[441], stage0_23[442], stage0_23[443]},
      {stage1_25[73],stage1_24[121],stage1_23[127],stage1_22[162],stage1_21[223]}
   );
   gpc615_5 gpc950 (
      {stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449], stage0_21[450]},
      {stage0_22[322]},
      {stage0_23[444], stage0_23[445], stage0_23[446], stage0_23[447], stage0_23[448], stage0_23[449]},
      {stage1_25[74],stage1_24[122],stage1_23[128],stage1_22[163],stage1_21[224]}
   );
   gpc615_5 gpc951 (
      {stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_22[323]},
      {stage0_23[450], stage0_23[451], stage0_23[452], stage0_23[453], stage0_23[454], stage0_23[455]},
      {stage1_25[75],stage1_24[123],stage1_23[129],stage1_22[164],stage1_21[225]}
   );
   gpc615_5 gpc952 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460]},
      {stage0_22[324]},
      {stage0_23[456], stage0_23[457], stage0_23[458], stage0_23[459], stage0_23[460], stage0_23[461]},
      {stage1_25[76],stage1_24[124],stage1_23[130],stage1_22[165],stage1_21[226]}
   );
   gpc615_5 gpc953 (
      {stage0_21[461], stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465]},
      {stage0_22[325]},
      {stage0_23[462], stage0_23[463], stage0_23[464], stage0_23[465], stage0_23[466], stage0_23[467]},
      {stage1_25[77],stage1_24[125],stage1_23[131],stage1_22[166],stage1_21[227]}
   );
   gpc615_5 gpc954 (
      {stage0_21[466], stage0_21[467], stage0_21[468], stage0_21[469], stage0_21[470]},
      {stage0_22[326]},
      {stage0_23[468], stage0_23[469], stage0_23[470], stage0_23[471], stage0_23[472], stage0_23[473]},
      {stage1_25[78],stage1_24[126],stage1_23[132],stage1_22[167],stage1_21[228]}
   );
   gpc606_5 gpc955 (
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331], stage0_22[332]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[79],stage1_24[127],stage1_23[133],stage1_22[168]}
   );
   gpc606_5 gpc956 (
      {stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336], stage0_22[337], stage0_22[338]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[80],stage1_24[128],stage1_23[134],stage1_22[169]}
   );
   gpc606_5 gpc957 (
      {stage0_22[339], stage0_22[340], stage0_22[341], stage0_22[342], stage0_22[343], stage0_22[344]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[81],stage1_24[129],stage1_23[135],stage1_22[170]}
   );
   gpc606_5 gpc958 (
      {stage0_22[345], stage0_22[346], stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[82],stage1_24[130],stage1_23[136],stage1_22[171]}
   );
   gpc606_5 gpc959 (
      {stage0_22[351], stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[83],stage1_24[131],stage1_23[137],stage1_22[172]}
   );
   gpc606_5 gpc960 (
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361], stage0_22[362]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[84],stage1_24[132],stage1_23[138],stage1_22[173]}
   );
   gpc606_5 gpc961 (
      {stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366], stage0_22[367], stage0_22[368]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[85],stage1_24[133],stage1_23[139],stage1_22[174]}
   );
   gpc606_5 gpc962 (
      {stage0_22[369], stage0_22[370], stage0_22[371], stage0_22[372], stage0_22[373], stage0_22[374]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[86],stage1_24[134],stage1_23[140],stage1_22[175]}
   );
   gpc606_5 gpc963 (
      {stage0_22[375], stage0_22[376], stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[87],stage1_24[135],stage1_23[141],stage1_22[176]}
   );
   gpc606_5 gpc964 (
      {stage0_22[381], stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[88],stage1_24[136],stage1_23[142],stage1_22[177]}
   );
   gpc606_5 gpc965 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391], stage0_22[392]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[89],stage1_24[137],stage1_23[143],stage1_22[178]}
   );
   gpc615_5 gpc966 (
      {stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396], stage0_22[397]},
      {stage0_23[474]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[90],stage1_24[138],stage1_23[144],stage1_22[179]}
   );
   gpc615_5 gpc967 (
      {stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401], stage0_22[402]},
      {stage0_23[475]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[91],stage1_24[139],stage1_23[145],stage1_22[180]}
   );
   gpc615_5 gpc968 (
      {stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406], stage0_22[407]},
      {stage0_23[476]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[92],stage1_24[140],stage1_23[146],stage1_22[181]}
   );
   gpc615_5 gpc969 (
      {stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411], stage0_22[412]},
      {stage0_23[477]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[93],stage1_24[141],stage1_23[147],stage1_22[182]}
   );
   gpc615_5 gpc970 (
      {stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416], stage0_22[417]},
      {stage0_23[478]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[94],stage1_24[142],stage1_23[148],stage1_22[183]}
   );
   gpc615_5 gpc971 (
      {stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421], stage0_22[422]},
      {stage0_23[479]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[95],stage1_24[143],stage1_23[149],stage1_22[184]}
   );
   gpc615_5 gpc972 (
      {stage0_23[480], stage0_23[481], stage0_23[482], stage0_23[483], stage0_23[484]},
      {stage0_24[102]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[17],stage1_25[96],stage1_24[144],stage1_23[150]}
   );
   gpc615_5 gpc973 (
      {stage0_23[485], stage0_23[486], stage0_23[487], stage0_23[488], stage0_23[489]},
      {stage0_24[103]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[18],stage1_25[97],stage1_24[145],stage1_23[151]}
   );
   gpc615_5 gpc974 (
      {stage0_23[490], stage0_23[491], stage0_23[492], stage0_23[493], stage0_23[494]},
      {stage0_24[104]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[19],stage1_25[98],stage1_24[146],stage1_23[152]}
   );
   gpc615_5 gpc975 (
      {stage0_23[495], stage0_23[496], stage0_23[497], stage0_23[498], stage0_23[499]},
      {stage0_24[105]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[20],stage1_25[99],stage1_24[147],stage1_23[153]}
   );
   gpc606_5 gpc976 (
      {stage0_24[106], stage0_24[107], stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[4],stage1_26[21],stage1_25[100],stage1_24[148]}
   );
   gpc606_5 gpc977 (
      {stage0_24[112], stage0_24[113], stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[5],stage1_26[22],stage1_25[101],stage1_24[149]}
   );
   gpc606_5 gpc978 (
      {stage0_24[118], stage0_24[119], stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[6],stage1_26[23],stage1_25[102],stage1_24[150]}
   );
   gpc606_5 gpc979 (
      {stage0_24[124], stage0_24[125], stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[7],stage1_26[24],stage1_25[103],stage1_24[151]}
   );
   gpc606_5 gpc980 (
      {stage0_24[130], stage0_24[131], stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[8],stage1_26[25],stage1_25[104],stage1_24[152]}
   );
   gpc606_5 gpc981 (
      {stage0_24[136], stage0_24[137], stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[9],stage1_26[26],stage1_25[105],stage1_24[153]}
   );
   gpc606_5 gpc982 (
      {stage0_24[142], stage0_24[143], stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[10],stage1_26[27],stage1_25[106],stage1_24[154]}
   );
   gpc606_5 gpc983 (
      {stage0_24[148], stage0_24[149], stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[11],stage1_26[28],stage1_25[107],stage1_24[155]}
   );
   gpc606_5 gpc984 (
      {stage0_24[154], stage0_24[155], stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[12],stage1_26[29],stage1_25[108],stage1_24[156]}
   );
   gpc606_5 gpc985 (
      {stage0_24[160], stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[13],stage1_26[30],stage1_25[109],stage1_24[157]}
   );
   gpc606_5 gpc986 (
      {stage0_24[166], stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170], stage0_24[171]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[14],stage1_26[31],stage1_25[110],stage1_24[158]}
   );
   gpc606_5 gpc987 (
      {stage0_24[172], stage0_24[173], stage0_24[174], stage0_24[175], stage0_24[176], stage0_24[177]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[15],stage1_26[32],stage1_25[111],stage1_24[159]}
   );
   gpc606_5 gpc988 (
      {stage0_24[178], stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[16],stage1_26[33],stage1_25[112],stage1_24[160]}
   );
   gpc606_5 gpc989 (
      {stage0_24[184], stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[17],stage1_26[34],stage1_25[113],stage1_24[161]}
   );
   gpc606_5 gpc990 (
      {stage0_24[190], stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[18],stage1_26[35],stage1_25[114],stage1_24[162]}
   );
   gpc606_5 gpc991 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200], stage0_24[201]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[19],stage1_26[36],stage1_25[115],stage1_24[163]}
   );
   gpc606_5 gpc992 (
      {stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205], stage0_24[206], stage0_24[207]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[20],stage1_26[37],stage1_25[116],stage1_24[164]}
   );
   gpc606_5 gpc993 (
      {stage0_24[208], stage0_24[209], stage0_24[210], stage0_24[211], stage0_24[212], stage0_24[213]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[21],stage1_26[38],stage1_25[117],stage1_24[165]}
   );
   gpc606_5 gpc994 (
      {stage0_24[214], stage0_24[215], stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[22],stage1_26[39],stage1_25[118],stage1_24[166]}
   );
   gpc606_5 gpc995 (
      {stage0_24[220], stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[23],stage1_26[40],stage1_25[119],stage1_24[167]}
   );
   gpc606_5 gpc996 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230], stage0_24[231]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[24],stage1_26[41],stage1_25[120],stage1_24[168]}
   );
   gpc606_5 gpc997 (
      {stage0_24[232], stage0_24[233], stage0_24[234], stage0_24[235], stage0_24[236], stage0_24[237]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[25],stage1_26[42],stage1_25[121],stage1_24[169]}
   );
   gpc606_5 gpc998 (
      {stage0_24[238], stage0_24[239], stage0_24[240], stage0_24[241], stage0_24[242], stage0_24[243]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[26],stage1_26[43],stage1_25[122],stage1_24[170]}
   );
   gpc606_5 gpc999 (
      {stage0_24[244], stage0_24[245], stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[27],stage1_26[44],stage1_25[123],stage1_24[171]}
   );
   gpc606_5 gpc1000 (
      {stage0_24[250], stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[28],stage1_26[45],stage1_25[124],stage1_24[172]}
   );
   gpc606_5 gpc1001 (
      {stage0_24[256], stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260], stage0_24[261]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[29],stage1_26[46],stage1_25[125],stage1_24[173]}
   );
   gpc606_5 gpc1002 (
      {stage0_24[262], stage0_24[263], stage0_24[264], stage0_24[265], stage0_24[266], stage0_24[267]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[30],stage1_26[47],stage1_25[126],stage1_24[174]}
   );
   gpc606_5 gpc1003 (
      {stage0_24[268], stage0_24[269], stage0_24[270], stage0_24[271], stage0_24[272], stage0_24[273]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[31],stage1_26[48],stage1_25[127],stage1_24[175]}
   );
   gpc606_5 gpc1004 (
      {stage0_24[274], stage0_24[275], stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[32],stage1_26[49],stage1_25[128],stage1_24[176]}
   );
   gpc606_5 gpc1005 (
      {stage0_24[280], stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[33],stage1_26[50],stage1_25[129],stage1_24[177]}
   );
   gpc606_5 gpc1006 (
      {stage0_24[286], stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290], stage0_24[291]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[34],stage1_26[51],stage1_25[130],stage1_24[178]}
   );
   gpc606_5 gpc1007 (
      {stage0_24[292], stage0_24[293], stage0_24[294], stage0_24[295], stage0_24[296], stage0_24[297]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[35],stage1_26[52],stage1_25[131],stage1_24[179]}
   );
   gpc606_5 gpc1008 (
      {stage0_24[298], stage0_24[299], stage0_24[300], stage0_24[301], stage0_24[302], stage0_24[303]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[36],stage1_26[53],stage1_25[132],stage1_24[180]}
   );
   gpc606_5 gpc1009 (
      {stage0_24[304], stage0_24[305], stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[37],stage1_26[54],stage1_25[133],stage1_24[181]}
   );
   gpc606_5 gpc1010 (
      {stage0_24[310], stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[38],stage1_26[55],stage1_25[134],stage1_24[182]}
   );
   gpc606_5 gpc1011 (
      {stage0_24[316], stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320], stage0_24[321]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[39],stage1_26[56],stage1_25[135],stage1_24[183]}
   );
   gpc606_5 gpc1012 (
      {stage0_24[322], stage0_24[323], stage0_24[324], stage0_24[325], stage0_24[326], stage0_24[327]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[40],stage1_26[57],stage1_25[136],stage1_24[184]}
   );
   gpc606_5 gpc1013 (
      {stage0_24[328], stage0_24[329], stage0_24[330], stage0_24[331], stage0_24[332], stage0_24[333]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[41],stage1_26[58],stage1_25[137],stage1_24[185]}
   );
   gpc606_5 gpc1014 (
      {stage0_24[334], stage0_24[335], stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[42],stage1_26[59],stage1_25[138],stage1_24[186]}
   );
   gpc606_5 gpc1015 (
      {stage0_24[340], stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[43],stage1_26[60],stage1_25[139],stage1_24[187]}
   );
   gpc606_5 gpc1016 (
      {stage0_24[346], stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350], stage0_24[351]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[44],stage1_26[61],stage1_25[140],stage1_24[188]}
   );
   gpc615_5 gpc1017 (
      {stage0_24[352], stage0_24[353], stage0_24[354], stage0_24[355], stage0_24[356]},
      {stage0_25[24]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[45],stage1_26[62],stage1_25[141],stage1_24[189]}
   );
   gpc615_5 gpc1018 (
      {stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360], stage0_24[361]},
      {stage0_25[25]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[46],stage1_26[63],stage1_25[142],stage1_24[190]}
   );
   gpc615_5 gpc1019 (
      {stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365], stage0_24[366]},
      {stage0_25[26]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[47],stage1_26[64],stage1_25[143],stage1_24[191]}
   );
   gpc615_5 gpc1020 (
      {stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370], stage0_24[371]},
      {stage0_25[27]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[48],stage1_26[65],stage1_25[144],stage1_24[192]}
   );
   gpc615_5 gpc1021 (
      {stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375], stage0_24[376]},
      {stage0_25[28]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[49],stage1_26[66],stage1_25[145],stage1_24[193]}
   );
   gpc615_5 gpc1022 (
      {stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380], stage0_24[381]},
      {stage0_25[29]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[50],stage1_26[67],stage1_25[146],stage1_24[194]}
   );
   gpc615_5 gpc1023 (
      {stage0_24[382], stage0_24[383], stage0_24[384], stage0_24[385], stage0_24[386]},
      {stage0_25[30]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[51],stage1_26[68],stage1_25[147],stage1_24[195]}
   );
   gpc615_5 gpc1024 (
      {stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390], stage0_24[391]},
      {stage0_25[31]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[52],stage1_26[69],stage1_25[148],stage1_24[196]}
   );
   gpc615_5 gpc1025 (
      {stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395], stage0_24[396]},
      {stage0_25[32]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[53],stage1_26[70],stage1_25[149],stage1_24[197]}
   );
   gpc615_5 gpc1026 (
      {stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400], stage0_24[401]},
      {stage0_25[33]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[54],stage1_26[71],stage1_25[150],stage1_24[198]}
   );
   gpc615_5 gpc1027 (
      {stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405], stage0_24[406]},
      {stage0_25[34]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[55],stage1_26[72],stage1_25[151],stage1_24[199]}
   );
   gpc615_5 gpc1028 (
      {stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410], stage0_24[411]},
      {stage0_25[35]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[56],stage1_26[73],stage1_25[152],stage1_24[200]}
   );
   gpc615_5 gpc1029 (
      {stage0_24[412], stage0_24[413], stage0_24[414], stage0_24[415], stage0_24[416]},
      {stage0_25[36]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[57],stage1_26[74],stage1_25[153],stage1_24[201]}
   );
   gpc615_5 gpc1030 (
      {stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420], stage0_24[421]},
      {stage0_25[37]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[58],stage1_26[75],stage1_25[154],stage1_24[202]}
   );
   gpc615_5 gpc1031 (
      {stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425], stage0_24[426]},
      {stage0_25[38]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[59],stage1_26[76],stage1_25[155],stage1_24[203]}
   );
   gpc615_5 gpc1032 (
      {stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430], stage0_24[431]},
      {stage0_25[39]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[60],stage1_26[77],stage1_25[156],stage1_24[204]}
   );
   gpc615_5 gpc1033 (
      {stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435], stage0_24[436]},
      {stage0_25[40]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[61],stage1_26[78],stage1_25[157],stage1_24[205]}
   );
   gpc615_5 gpc1034 (
      {stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440], stage0_24[441]},
      {stage0_25[41]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[62],stage1_26[79],stage1_25[158],stage1_24[206]}
   );
   gpc615_5 gpc1035 (
      {stage0_24[442], stage0_24[443], stage0_24[444], stage0_24[445], stage0_24[446]},
      {stage0_25[42]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[63],stage1_26[80],stage1_25[159],stage1_24[207]}
   );
   gpc615_5 gpc1036 (
      {stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450], stage0_24[451]},
      {stage0_25[43]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[64],stage1_26[81],stage1_25[160],stage1_24[208]}
   );
   gpc615_5 gpc1037 (
      {stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455], stage0_24[456]},
      {stage0_25[44]},
      {stage0_26[366], stage0_26[367], stage0_26[368], stage0_26[369], stage0_26[370], stage0_26[371]},
      {stage1_28[61],stage1_27[65],stage1_26[82],stage1_25[161],stage1_24[209]}
   );
   gpc615_5 gpc1038 (
      {stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460], stage0_24[461]},
      {stage0_25[45]},
      {stage0_26[372], stage0_26[373], stage0_26[374], stage0_26[375], stage0_26[376], stage0_26[377]},
      {stage1_28[62],stage1_27[66],stage1_26[83],stage1_25[162],stage1_24[210]}
   );
   gpc615_5 gpc1039 (
      {stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465], stage0_24[466]},
      {stage0_25[46]},
      {stage0_26[378], stage0_26[379], stage0_26[380], stage0_26[381], stage0_26[382], stage0_26[383]},
      {stage1_28[63],stage1_27[67],stage1_26[84],stage1_25[163],stage1_24[211]}
   );
   gpc615_5 gpc1040 (
      {stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470], stage0_24[471]},
      {stage0_25[47]},
      {stage0_26[384], stage0_26[385], stage0_26[386], stage0_26[387], stage0_26[388], stage0_26[389]},
      {stage1_28[64],stage1_27[68],stage1_26[85],stage1_25[164],stage1_24[212]}
   );
   gpc615_5 gpc1041 (
      {stage0_24[472], stage0_24[473], stage0_24[474], stage0_24[475], stage0_24[476]},
      {stage0_25[48]},
      {stage0_26[390], stage0_26[391], stage0_26[392], stage0_26[393], stage0_26[394], stage0_26[395]},
      {stage1_28[65],stage1_27[69],stage1_26[86],stage1_25[165],stage1_24[213]}
   );
   gpc615_5 gpc1042 (
      {stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480], stage0_24[481]},
      {stage0_25[49]},
      {stage0_26[396], stage0_26[397], stage0_26[398], stage0_26[399], stage0_26[400], stage0_26[401]},
      {stage1_28[66],stage1_27[70],stage1_26[87],stage1_25[166],stage1_24[214]}
   );
   gpc615_5 gpc1043 (
      {stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485], stage0_24[486]},
      {stage0_25[50]},
      {stage0_26[402], stage0_26[403], stage0_26[404], stage0_26[405], stage0_26[406], stage0_26[407]},
      {stage1_28[67],stage1_27[71],stage1_26[88],stage1_25[167],stage1_24[215]}
   );
   gpc615_5 gpc1044 (
      {stage0_24[487], stage0_24[488], stage0_24[489], stage0_24[490], stage0_24[491]},
      {stage0_25[51]},
      {stage0_26[408], stage0_26[409], stage0_26[410], stage0_26[411], stage0_26[412], stage0_26[413]},
      {stage1_28[68],stage1_27[72],stage1_26[89],stage1_25[168],stage1_24[216]}
   );
   gpc615_5 gpc1045 (
      {stage0_24[492], stage0_24[493], stage0_24[494], stage0_24[495], stage0_24[496]},
      {stage0_25[52]},
      {stage0_26[414], stage0_26[415], stage0_26[416], stage0_26[417], stage0_26[418], stage0_26[419]},
      {stage1_28[69],stage1_27[73],stage1_26[90],stage1_25[169],stage1_24[217]}
   );
   gpc615_5 gpc1046 (
      {stage0_24[497], stage0_24[498], stage0_24[499], stage0_24[500], stage0_24[501]},
      {stage0_25[53]},
      {stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423], stage0_26[424], stage0_26[425]},
      {stage1_28[70],stage1_27[74],stage1_26[91],stage1_25[170],stage1_24[218]}
   );
   gpc615_5 gpc1047 (
      {stage0_24[502], stage0_24[503], stage0_24[504], stage0_24[505], stage0_24[506]},
      {stage0_25[54]},
      {stage0_26[426], stage0_26[427], stage0_26[428], stage0_26[429], stage0_26[430], stage0_26[431]},
      {stage1_28[71],stage1_27[75],stage1_26[92],stage1_25[171],stage1_24[219]}
   );
   gpc615_5 gpc1048 (
      {stage0_24[507], stage0_24[508], stage0_24[509], stage0_24[510], stage0_24[511]},
      {stage0_25[55]},
      {stage0_26[432], stage0_26[433], stage0_26[434], stage0_26[435], stage0_26[436], stage0_26[437]},
      {stage1_28[72],stage1_27[76],stage1_26[93],stage1_25[172],stage1_24[220]}
   );
   gpc606_5 gpc1049 (
      {stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59], stage0_25[60], stage0_25[61]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[73],stage1_27[77],stage1_26[94],stage1_25[173]}
   );
   gpc606_5 gpc1050 (
      {stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65], stage0_25[66], stage0_25[67]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[74],stage1_27[78],stage1_26[95],stage1_25[174]}
   );
   gpc606_5 gpc1051 (
      {stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71], stage0_25[72], stage0_25[73]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[75],stage1_27[79],stage1_26[96],stage1_25[175]}
   );
   gpc606_5 gpc1052 (
      {stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77], stage0_25[78], stage0_25[79]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[76],stage1_27[80],stage1_26[97],stage1_25[176]}
   );
   gpc606_5 gpc1053 (
      {stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83], stage0_25[84], stage0_25[85]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[77],stage1_27[81],stage1_26[98],stage1_25[177]}
   );
   gpc606_5 gpc1054 (
      {stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89], stage0_25[90], stage0_25[91]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[78],stage1_27[82],stage1_26[99],stage1_25[178]}
   );
   gpc606_5 gpc1055 (
      {stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95], stage0_25[96], stage0_25[97]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[79],stage1_27[83],stage1_26[100],stage1_25[179]}
   );
   gpc606_5 gpc1056 (
      {stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101], stage0_25[102], stage0_25[103]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[80],stage1_27[84],stage1_26[101],stage1_25[180]}
   );
   gpc606_5 gpc1057 (
      {stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107], stage0_25[108], stage0_25[109]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[81],stage1_27[85],stage1_26[102],stage1_25[181]}
   );
   gpc606_5 gpc1058 (
      {stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113], stage0_25[114], stage0_25[115]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[82],stage1_27[86],stage1_26[103],stage1_25[182]}
   );
   gpc606_5 gpc1059 (
      {stage0_25[116], stage0_25[117], stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[83],stage1_27[87],stage1_26[104],stage1_25[183]}
   );
   gpc606_5 gpc1060 (
      {stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[84],stage1_27[88],stage1_26[105],stage1_25[184]}
   );
   gpc606_5 gpc1061 (
      {stage0_25[128], stage0_25[129], stage0_25[130], stage0_25[131], stage0_25[132], stage0_25[133]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[85],stage1_27[89],stage1_26[106],stage1_25[185]}
   );
   gpc606_5 gpc1062 (
      {stage0_25[134], stage0_25[135], stage0_25[136], stage0_25[137], stage0_25[138], stage0_25[139]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[86],stage1_27[90],stage1_26[107],stage1_25[186]}
   );
   gpc606_5 gpc1063 (
      {stage0_25[140], stage0_25[141], stage0_25[142], stage0_25[143], stage0_25[144], stage0_25[145]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[87],stage1_27[91],stage1_26[108],stage1_25[187]}
   );
   gpc606_5 gpc1064 (
      {stage0_25[146], stage0_25[147], stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[88],stage1_27[92],stage1_26[109],stage1_25[188]}
   );
   gpc606_5 gpc1065 (
      {stage0_25[152], stage0_25[153], stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[89],stage1_27[93],stage1_26[110],stage1_25[189]}
   );
   gpc606_5 gpc1066 (
      {stage0_25[158], stage0_25[159], stage0_25[160], stage0_25[161], stage0_25[162], stage0_25[163]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[90],stage1_27[94],stage1_26[111],stage1_25[190]}
   );
   gpc606_5 gpc1067 (
      {stage0_25[164], stage0_25[165], stage0_25[166], stage0_25[167], stage0_25[168], stage0_25[169]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[91],stage1_27[95],stage1_26[112],stage1_25[191]}
   );
   gpc606_5 gpc1068 (
      {stage0_25[170], stage0_25[171], stage0_25[172], stage0_25[173], stage0_25[174], stage0_25[175]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[92],stage1_27[96],stage1_26[113],stage1_25[192]}
   );
   gpc606_5 gpc1069 (
      {stage0_25[176], stage0_25[177], stage0_25[178], stage0_25[179], stage0_25[180], stage0_25[181]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[93],stage1_27[97],stage1_26[114],stage1_25[193]}
   );
   gpc606_5 gpc1070 (
      {stage0_25[182], stage0_25[183], stage0_25[184], stage0_25[185], stage0_25[186], stage0_25[187]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[94],stage1_27[98],stage1_26[115],stage1_25[194]}
   );
   gpc606_5 gpc1071 (
      {stage0_25[188], stage0_25[189], stage0_25[190], stage0_25[191], stage0_25[192], stage0_25[193]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[95],stage1_27[99],stage1_26[116],stage1_25[195]}
   );
   gpc606_5 gpc1072 (
      {stage0_25[194], stage0_25[195], stage0_25[196], stage0_25[197], stage0_25[198], stage0_25[199]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[96],stage1_27[100],stage1_26[117],stage1_25[196]}
   );
   gpc606_5 gpc1073 (
      {stage0_25[200], stage0_25[201], stage0_25[202], stage0_25[203], stage0_25[204], stage0_25[205]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[97],stage1_27[101],stage1_26[118],stage1_25[197]}
   );
   gpc606_5 gpc1074 (
      {stage0_25[206], stage0_25[207], stage0_25[208], stage0_25[209], stage0_25[210], stage0_25[211]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[98],stage1_27[102],stage1_26[119],stage1_25[198]}
   );
   gpc606_5 gpc1075 (
      {stage0_25[212], stage0_25[213], stage0_25[214], stage0_25[215], stage0_25[216], stage0_25[217]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[99],stage1_27[103],stage1_26[120],stage1_25[199]}
   );
   gpc606_5 gpc1076 (
      {stage0_25[218], stage0_25[219], stage0_25[220], stage0_25[221], stage0_25[222], stage0_25[223]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[100],stage1_27[104],stage1_26[121],stage1_25[200]}
   );
   gpc606_5 gpc1077 (
      {stage0_25[224], stage0_25[225], stage0_25[226], stage0_25[227], stage0_25[228], stage0_25[229]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[101],stage1_27[105],stage1_26[122],stage1_25[201]}
   );
   gpc606_5 gpc1078 (
      {stage0_25[230], stage0_25[231], stage0_25[232], stage0_25[233], stage0_25[234], stage0_25[235]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[102],stage1_27[106],stage1_26[123],stage1_25[202]}
   );
   gpc606_5 gpc1079 (
      {stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239], stage0_25[240], stage0_25[241]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[103],stage1_27[107],stage1_26[124],stage1_25[203]}
   );
   gpc606_5 gpc1080 (
      {stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245], stage0_25[246], stage0_25[247]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[104],stage1_27[108],stage1_26[125],stage1_25[204]}
   );
   gpc606_5 gpc1081 (
      {stage0_25[248], stage0_25[249], stage0_25[250], stage0_25[251], stage0_25[252], stage0_25[253]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[105],stage1_27[109],stage1_26[126],stage1_25[205]}
   );
   gpc606_5 gpc1082 (
      {stage0_25[254], stage0_25[255], stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[106],stage1_27[110],stage1_26[127],stage1_25[206]}
   );
   gpc606_5 gpc1083 (
      {stage0_25[260], stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[107],stage1_27[111],stage1_26[128],stage1_25[207]}
   );
   gpc606_5 gpc1084 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270], stage0_25[271]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[108],stage1_27[112],stage1_26[129],stage1_25[208]}
   );
   gpc606_5 gpc1085 (
      {stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275], stage0_25[276], stage0_25[277]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[109],stage1_27[113],stage1_26[130],stage1_25[209]}
   );
   gpc606_5 gpc1086 (
      {stage0_25[278], stage0_25[279], stage0_25[280], stage0_25[281], stage0_25[282], stage0_25[283]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[110],stage1_27[114],stage1_26[131],stage1_25[210]}
   );
   gpc606_5 gpc1087 (
      {stage0_25[284], stage0_25[285], stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[111],stage1_27[115],stage1_26[132],stage1_25[211]}
   );
   gpc606_5 gpc1088 (
      {stage0_25[290], stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[112],stage1_27[116],stage1_26[133],stage1_25[212]}
   );
   gpc606_5 gpc1089 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300], stage0_25[301]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[113],stage1_27[117],stage1_26[134],stage1_25[213]}
   );
   gpc606_5 gpc1090 (
      {stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305], stage0_25[306], stage0_25[307]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[114],stage1_27[118],stage1_26[135],stage1_25[214]}
   );
   gpc606_5 gpc1091 (
      {stage0_25[308], stage0_25[309], stage0_25[310], stage0_25[311], stage0_25[312], stage0_25[313]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[115],stage1_27[119],stage1_26[136],stage1_25[215]}
   );
   gpc606_5 gpc1092 (
      {stage0_25[314], stage0_25[315], stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[116],stage1_27[120],stage1_26[137],stage1_25[216]}
   );
   gpc606_5 gpc1093 (
      {stage0_25[320], stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[117],stage1_27[121],stage1_26[138],stage1_25[217]}
   );
   gpc606_5 gpc1094 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330], stage0_25[331]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[118],stage1_27[122],stage1_26[139],stage1_25[218]}
   );
   gpc606_5 gpc1095 (
      {stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335], stage0_25[336], stage0_25[337]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[119],stage1_27[123],stage1_26[140],stage1_25[219]}
   );
   gpc606_5 gpc1096 (
      {stage0_25[338], stage0_25[339], stage0_25[340], stage0_25[341], stage0_25[342], stage0_25[343]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[120],stage1_27[124],stage1_26[141],stage1_25[220]}
   );
   gpc606_5 gpc1097 (
      {stage0_25[344], stage0_25[345], stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[121],stage1_27[125],stage1_26[142],stage1_25[221]}
   );
   gpc606_5 gpc1098 (
      {stage0_25[350], stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[122],stage1_27[126],stage1_26[143],stage1_25[222]}
   );
   gpc606_5 gpc1099 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360], stage0_25[361]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[123],stage1_27[127],stage1_26[144],stage1_25[223]}
   );
   gpc606_5 gpc1100 (
      {stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365], stage0_25[366], stage0_25[367]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[124],stage1_27[128],stage1_26[145],stage1_25[224]}
   );
   gpc606_5 gpc1101 (
      {stage0_25[368], stage0_25[369], stage0_25[370], stage0_25[371], stage0_25[372], stage0_25[373]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[125],stage1_27[129],stage1_26[146],stage1_25[225]}
   );
   gpc606_5 gpc1102 (
      {stage0_25[374], stage0_25[375], stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[126],stage1_27[130],stage1_26[147],stage1_25[226]}
   );
   gpc606_5 gpc1103 (
      {stage0_25[380], stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327], stage0_27[328], stage0_27[329]},
      {stage1_29[54],stage1_28[127],stage1_27[131],stage1_26[148],stage1_25[227]}
   );
   gpc606_5 gpc1104 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390], stage0_25[391]},
      {stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[55],stage1_28[128],stage1_27[132],stage1_26[149],stage1_25[228]}
   );
   gpc606_5 gpc1105 (
      {stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395], stage0_25[396], stage0_25[397]},
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341]},
      {stage1_29[56],stage1_28[129],stage1_27[133],stage1_26[150],stage1_25[229]}
   );
   gpc606_5 gpc1106 (
      {stage0_25[398], stage0_25[399], stage0_25[400], stage0_25[401], stage0_25[402], stage0_25[403]},
      {stage0_27[342], stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage1_29[57],stage1_28[130],stage1_27[134],stage1_26[151],stage1_25[230]}
   );
   gpc606_5 gpc1107 (
      {stage0_25[404], stage0_25[405], stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409]},
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352], stage0_27[353]},
      {stage1_29[58],stage1_28[131],stage1_27[135],stage1_26[152],stage1_25[231]}
   );
   gpc606_5 gpc1108 (
      {stage0_25[410], stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357], stage0_27[358], stage0_27[359]},
      {stage1_29[59],stage1_28[132],stage1_27[136],stage1_26[153],stage1_25[232]}
   );
   gpc606_5 gpc1109 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420], stage0_25[421]},
      {stage0_27[360], stage0_27[361], stage0_27[362], stage0_27[363], stage0_27[364], stage0_27[365]},
      {stage1_29[60],stage1_28[133],stage1_27[137],stage1_26[154],stage1_25[233]}
   );
   gpc606_5 gpc1110 (
      {stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425], stage0_25[426], stage0_25[427]},
      {stage0_27[366], stage0_27[367], stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371]},
      {stage1_29[61],stage1_28[134],stage1_27[138],stage1_26[155],stage1_25[234]}
   );
   gpc606_5 gpc1111 (
      {stage0_25[428], stage0_25[429], stage0_25[430], stage0_25[431], stage0_25[432], stage0_25[433]},
      {stage0_27[372], stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage1_29[62],stage1_28[135],stage1_27[139],stage1_26[156],stage1_25[235]}
   );
   gpc606_5 gpc1112 (
      {stage0_25[434], stage0_25[435], stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439]},
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382], stage0_27[383]},
      {stage1_29[63],stage1_28[136],stage1_27[140],stage1_26[157],stage1_25[236]}
   );
   gpc606_5 gpc1113 (
      {stage0_25[440], stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387], stage0_27[388], stage0_27[389]},
      {stage1_29[64],stage1_28[137],stage1_27[141],stage1_26[158],stage1_25[237]}
   );
   gpc606_5 gpc1114 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450], stage0_25[451]},
      {stage0_27[390], stage0_27[391], stage0_27[392], stage0_27[393], stage0_27[394], stage0_27[395]},
      {stage1_29[65],stage1_28[138],stage1_27[142],stage1_26[159],stage1_25[238]}
   );
   gpc606_5 gpc1115 (
      {stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455], stage0_25[456], stage0_25[457]},
      {stage0_27[396], stage0_27[397], stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401]},
      {stage1_29[66],stage1_28[139],stage1_27[143],stage1_26[160],stage1_25[239]}
   );
   gpc606_5 gpc1116 (
      {stage0_25[458], stage0_25[459], stage0_25[460], stage0_25[461], stage0_25[462], stage0_25[463]},
      {stage0_27[402], stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage1_29[67],stage1_28[140],stage1_27[144],stage1_26[161],stage1_25[240]}
   );
   gpc606_5 gpc1117 (
      {stage0_25[464], stage0_25[465], stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469]},
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412], stage0_27[413]},
      {stage1_29[68],stage1_28[141],stage1_27[145],stage1_26[162],stage1_25[241]}
   );
   gpc606_5 gpc1118 (
      {stage0_25[470], stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417], stage0_27[418], stage0_27[419]},
      {stage1_29[69],stage1_28[142],stage1_27[146],stage1_26[163],stage1_25[242]}
   );
   gpc606_5 gpc1119 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480], stage0_25[481]},
      {stage0_27[420], stage0_27[421], stage0_27[422], stage0_27[423], stage0_27[424], stage0_27[425]},
      {stage1_29[70],stage1_28[143],stage1_27[147],stage1_26[164],stage1_25[243]}
   );
   gpc615_5 gpc1120 (
      {stage0_26[438], stage0_26[439], stage0_26[440], stage0_26[441], stage0_26[442]},
      {stage0_27[426]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[71],stage1_28[144],stage1_27[148],stage1_26[165]}
   );
   gpc615_5 gpc1121 (
      {stage0_26[443], stage0_26[444], stage0_26[445], stage0_26[446], stage0_26[447]},
      {stage0_27[427]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[72],stage1_28[145],stage1_27[149],stage1_26[166]}
   );
   gpc615_5 gpc1122 (
      {stage0_26[448], stage0_26[449], stage0_26[450], stage0_26[451], stage0_26[452]},
      {stage0_27[428]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[73],stage1_28[146],stage1_27[150],stage1_26[167]}
   );
   gpc615_5 gpc1123 (
      {stage0_26[453], stage0_26[454], stage0_26[455], stage0_26[456], stage0_26[457]},
      {stage0_27[429]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[74],stage1_28[147],stage1_27[151],stage1_26[168]}
   );
   gpc615_5 gpc1124 (
      {stage0_26[458], stage0_26[459], stage0_26[460], stage0_26[461], stage0_26[462]},
      {stage0_27[430]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[75],stage1_28[148],stage1_27[152],stage1_26[169]}
   );
   gpc615_5 gpc1125 (
      {stage0_26[463], stage0_26[464], stage0_26[465], stage0_26[466], stage0_26[467]},
      {stage0_27[431]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[76],stage1_28[149],stage1_27[153],stage1_26[170]}
   );
   gpc615_5 gpc1126 (
      {stage0_26[468], stage0_26[469], stage0_26[470], stage0_26[471], stage0_26[472]},
      {stage0_27[432]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[77],stage1_28[150],stage1_27[154],stage1_26[171]}
   );
   gpc615_5 gpc1127 (
      {stage0_26[473], stage0_26[474], stage0_26[475], stage0_26[476], stage0_26[477]},
      {stage0_27[433]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[78],stage1_28[151],stage1_27[155],stage1_26[172]}
   );
   gpc615_5 gpc1128 (
      {stage0_26[478], stage0_26[479], stage0_26[480], stage0_26[481], stage0_26[482]},
      {stage0_27[434]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[79],stage1_28[152],stage1_27[156],stage1_26[173]}
   );
   gpc615_5 gpc1129 (
      {stage0_26[483], stage0_26[484], stage0_26[485], stage0_26[486], stage0_26[487]},
      {stage0_27[435]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[80],stage1_28[153],stage1_27[157],stage1_26[174]}
   );
   gpc615_5 gpc1130 (
      {stage0_26[488], stage0_26[489], stage0_26[490], stage0_26[491], stage0_26[492]},
      {stage0_27[436]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[81],stage1_28[154],stage1_27[158],stage1_26[175]}
   );
   gpc615_5 gpc1131 (
      {stage0_26[493], stage0_26[494], stage0_26[495], stage0_26[496], stage0_26[497]},
      {stage0_27[437]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[82],stage1_28[155],stage1_27[159],stage1_26[176]}
   );
   gpc606_5 gpc1132 (
      {stage0_27[438], stage0_27[439], stage0_27[440], stage0_27[441], stage0_27[442], stage0_27[443]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[12],stage1_29[83],stage1_28[156],stage1_27[160]}
   );
   gpc606_5 gpc1133 (
      {stage0_27[444], stage0_27[445], stage0_27[446], stage0_27[447], stage0_27[448], stage0_27[449]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[13],stage1_29[84],stage1_28[157],stage1_27[161]}
   );
   gpc606_5 gpc1134 (
      {stage0_27[450], stage0_27[451], stage0_27[452], stage0_27[453], stage0_27[454], stage0_27[455]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[14],stage1_29[85],stage1_28[158],stage1_27[162]}
   );
   gpc606_5 gpc1135 (
      {stage0_27[456], stage0_27[457], stage0_27[458], stage0_27[459], stage0_27[460], stage0_27[461]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[15],stage1_29[86],stage1_28[159],stage1_27[163]}
   );
   gpc606_5 gpc1136 (
      {stage0_27[462], stage0_27[463], stage0_27[464], stage0_27[465], stage0_27[466], stage0_27[467]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[16],stage1_29[87],stage1_28[160],stage1_27[164]}
   );
   gpc606_5 gpc1137 (
      {stage0_27[468], stage0_27[469], stage0_27[470], stage0_27[471], stage0_27[472], stage0_27[473]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[17],stage1_29[88],stage1_28[161],stage1_27[165]}
   );
   gpc615_5 gpc1138 (
      {stage0_27[474], stage0_27[475], stage0_27[476], stage0_27[477], stage0_27[478]},
      {stage0_28[72]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[18],stage1_29[89],stage1_28[162],stage1_27[166]}
   );
   gpc606_5 gpc1139 (
      {stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[7],stage1_30[19],stage1_29[90],stage1_28[163]}
   );
   gpc606_5 gpc1140 (
      {stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[8],stage1_30[20],stage1_29[91],stage1_28[164]}
   );
   gpc606_5 gpc1141 (
      {stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[9],stage1_30[21],stage1_29[92],stage1_28[165]}
   );
   gpc606_5 gpc1142 (
      {stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[10],stage1_30[22],stage1_29[93],stage1_28[166]}
   );
   gpc606_5 gpc1143 (
      {stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[11],stage1_30[23],stage1_29[94],stage1_28[167]}
   );
   gpc606_5 gpc1144 (
      {stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[12],stage1_30[24],stage1_29[95],stage1_28[168]}
   );
   gpc606_5 gpc1145 (
      {stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[13],stage1_30[25],stage1_29[96],stage1_28[169]}
   );
   gpc606_5 gpc1146 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[14],stage1_30[26],stage1_29[97],stage1_28[170]}
   );
   gpc606_5 gpc1147 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[15],stage1_30[27],stage1_29[98],stage1_28[171]}
   );
   gpc606_5 gpc1148 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[16],stage1_30[28],stage1_29[99],stage1_28[172]}
   );
   gpc606_5 gpc1149 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[17],stage1_30[29],stage1_29[100],stage1_28[173]}
   );
   gpc606_5 gpc1150 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[18],stage1_30[30],stage1_29[101],stage1_28[174]}
   );
   gpc606_5 gpc1151 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[19],stage1_30[31],stage1_29[102],stage1_28[175]}
   );
   gpc606_5 gpc1152 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[20],stage1_30[32],stage1_29[103],stage1_28[176]}
   );
   gpc606_5 gpc1153 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[21],stage1_30[33],stage1_29[104],stage1_28[177]}
   );
   gpc606_5 gpc1154 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[22],stage1_30[34],stage1_29[105],stage1_28[178]}
   );
   gpc606_5 gpc1155 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[23],stage1_30[35],stage1_29[106],stage1_28[179]}
   );
   gpc606_5 gpc1156 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[24],stage1_30[36],stage1_29[107],stage1_28[180]}
   );
   gpc606_5 gpc1157 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[25],stage1_30[37],stage1_29[108],stage1_28[181]}
   );
   gpc606_5 gpc1158 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[26],stage1_30[38],stage1_29[109],stage1_28[182]}
   );
   gpc606_5 gpc1159 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[27],stage1_30[39],stage1_29[110],stage1_28[183]}
   );
   gpc606_5 gpc1160 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[28],stage1_30[40],stage1_29[111],stage1_28[184]}
   );
   gpc606_5 gpc1161 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[29],stage1_30[41],stage1_29[112],stage1_28[185]}
   );
   gpc606_5 gpc1162 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[30],stage1_30[42],stage1_29[113],stage1_28[186]}
   );
   gpc606_5 gpc1163 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[31],stage1_30[43],stage1_29[114],stage1_28[187]}
   );
   gpc606_5 gpc1164 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[32],stage1_30[44],stage1_29[115],stage1_28[188]}
   );
   gpc606_5 gpc1165 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[33],stage1_30[45],stage1_29[116],stage1_28[189]}
   );
   gpc606_5 gpc1166 (
      {stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239], stage0_28[240]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[34],stage1_30[46],stage1_29[117],stage1_28[190]}
   );
   gpc606_5 gpc1167 (
      {stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245], stage0_28[246]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[35],stage1_30[47],stage1_29[118],stage1_28[191]}
   );
   gpc606_5 gpc1168 (
      {stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251], stage0_28[252]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[36],stage1_30[48],stage1_29[119],stage1_28[192]}
   );
   gpc606_5 gpc1169 (
      {stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257], stage0_28[258]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[37],stage1_30[49],stage1_29[120],stage1_28[193]}
   );
   gpc606_5 gpc1170 (
      {stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263], stage0_28[264]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[38],stage1_30[50],stage1_29[121],stage1_28[194]}
   );
   gpc606_5 gpc1171 (
      {stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269], stage0_28[270]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[39],stage1_30[51],stage1_29[122],stage1_28[195]}
   );
   gpc606_5 gpc1172 (
      {stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275], stage0_28[276]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[40],stage1_30[52],stage1_29[123],stage1_28[196]}
   );
   gpc606_5 gpc1173 (
      {stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281], stage0_28[282]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[41],stage1_30[53],stage1_29[124],stage1_28[197]}
   );
   gpc606_5 gpc1174 (
      {stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287], stage0_28[288]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[42],stage1_30[54],stage1_29[125],stage1_28[198]}
   );
   gpc606_5 gpc1175 (
      {stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293], stage0_28[294]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[43],stage1_30[55],stage1_29[126],stage1_28[199]}
   );
   gpc606_5 gpc1176 (
      {stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299], stage0_28[300]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[44],stage1_30[56],stage1_29[127],stage1_28[200]}
   );
   gpc615_5 gpc1177 (
      {stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305]},
      {stage0_29[42]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[45],stage1_30[57],stage1_29[128],stage1_28[201]}
   );
   gpc615_5 gpc1178 (
      {stage0_28[306], stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310]},
      {stage0_29[43]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[46],stage1_30[58],stage1_29[129],stage1_28[202]}
   );
   gpc615_5 gpc1179 (
      {stage0_28[311], stage0_28[312], stage0_28[313], stage0_28[314], stage0_28[315]},
      {stage0_29[44]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[47],stage1_30[59],stage1_29[130],stage1_28[203]}
   );
   gpc615_5 gpc1180 (
      {stage0_28[316], stage0_28[317], stage0_28[318], stage0_28[319], stage0_28[320]},
      {stage0_29[45]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[48],stage1_30[60],stage1_29[131],stage1_28[204]}
   );
   gpc615_5 gpc1181 (
      {stage0_28[321], stage0_28[322], stage0_28[323], stage0_28[324], stage0_28[325]},
      {stage0_29[46]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[49],stage1_30[61],stage1_29[132],stage1_28[205]}
   );
   gpc615_5 gpc1182 (
      {stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329], stage0_28[330]},
      {stage0_29[47]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[50],stage1_30[62],stage1_29[133],stage1_28[206]}
   );
   gpc615_5 gpc1183 (
      {stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335]},
      {stage0_29[48]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[51],stage1_30[63],stage1_29[134],stage1_28[207]}
   );
   gpc615_5 gpc1184 (
      {stage0_28[336], stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340]},
      {stage0_29[49]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[52],stage1_30[64],stage1_29[135],stage1_28[208]}
   );
   gpc615_5 gpc1185 (
      {stage0_28[341], stage0_28[342], stage0_28[343], stage0_28[344], stage0_28[345]},
      {stage0_29[50]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[53],stage1_30[65],stage1_29[136],stage1_28[209]}
   );
   gpc615_5 gpc1186 (
      {stage0_28[346], stage0_28[347], stage0_28[348], stage0_28[349], stage0_28[350]},
      {stage0_29[51]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[54],stage1_30[66],stage1_29[137],stage1_28[210]}
   );
   gpc615_5 gpc1187 (
      {stage0_28[351], stage0_28[352], stage0_28[353], stage0_28[354], stage0_28[355]},
      {stage0_29[52]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[55],stage1_30[67],stage1_29[138],stage1_28[211]}
   );
   gpc615_5 gpc1188 (
      {stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359], stage0_28[360]},
      {stage0_29[53]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[56],stage1_30[68],stage1_29[139],stage1_28[212]}
   );
   gpc615_5 gpc1189 (
      {stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365]},
      {stage0_29[54]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[57],stage1_30[69],stage1_29[140],stage1_28[213]}
   );
   gpc615_5 gpc1190 (
      {stage0_28[366], stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370]},
      {stage0_29[55]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[58],stage1_30[70],stage1_29[141],stage1_28[214]}
   );
   gpc615_5 gpc1191 (
      {stage0_28[371], stage0_28[372], stage0_28[373], stage0_28[374], stage0_28[375]},
      {stage0_29[56]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[59],stage1_30[71],stage1_29[142],stage1_28[215]}
   );
   gpc615_5 gpc1192 (
      {stage0_28[376], stage0_28[377], stage0_28[378], stage0_28[379], stage0_28[380]},
      {stage0_29[57]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[60],stage1_30[72],stage1_29[143],stage1_28[216]}
   );
   gpc615_5 gpc1193 (
      {stage0_28[381], stage0_28[382], stage0_28[383], stage0_28[384], stage0_28[385]},
      {stage0_29[58]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[61],stage1_30[73],stage1_29[144],stage1_28[217]}
   );
   gpc615_5 gpc1194 (
      {stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389], stage0_28[390]},
      {stage0_29[59]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[62],stage1_30[74],stage1_29[145],stage1_28[218]}
   );
   gpc615_5 gpc1195 (
      {stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395]},
      {stage0_29[60]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[63],stage1_30[75],stage1_29[146],stage1_28[219]}
   );
   gpc615_5 gpc1196 (
      {stage0_28[396], stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400]},
      {stage0_29[61]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[64],stage1_30[76],stage1_29[147],stage1_28[220]}
   );
   gpc615_5 gpc1197 (
      {stage0_28[401], stage0_28[402], stage0_28[403], stage0_28[404], stage0_28[405]},
      {stage0_29[62]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[65],stage1_30[77],stage1_29[148],stage1_28[221]}
   );
   gpc615_5 gpc1198 (
      {stage0_28[406], stage0_28[407], stage0_28[408], stage0_28[409], stage0_28[410]},
      {stage0_29[63]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[66],stage1_30[78],stage1_29[149],stage1_28[222]}
   );
   gpc615_5 gpc1199 (
      {stage0_28[411], stage0_28[412], stage0_28[413], stage0_28[414], stage0_28[415]},
      {stage0_29[64]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[67],stage1_30[79],stage1_29[150],stage1_28[223]}
   );
   gpc615_5 gpc1200 (
      {stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419], stage0_28[420]},
      {stage0_29[65]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[68],stage1_30[80],stage1_29[151],stage1_28[224]}
   );
   gpc615_5 gpc1201 (
      {stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425]},
      {stage0_29[66]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[69],stage1_30[81],stage1_29[152],stage1_28[225]}
   );
   gpc615_5 gpc1202 (
      {stage0_28[426], stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430]},
      {stage0_29[67]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[70],stage1_30[82],stage1_29[153],stage1_28[226]}
   );
   gpc615_5 gpc1203 (
      {stage0_28[431], stage0_28[432], stage0_28[433], stage0_28[434], stage0_28[435]},
      {stage0_29[68]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[71],stage1_30[83],stage1_29[154],stage1_28[227]}
   );
   gpc615_5 gpc1204 (
      {stage0_28[436], stage0_28[437], stage0_28[438], stage0_28[439], stage0_28[440]},
      {stage0_29[69]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[72],stage1_30[84],stage1_29[155],stage1_28[228]}
   );
   gpc615_5 gpc1205 (
      {stage0_28[441], stage0_28[442], stage0_28[443], stage0_28[444], stage0_28[445]},
      {stage0_29[70]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[73],stage1_30[85],stage1_29[156],stage1_28[229]}
   );
   gpc615_5 gpc1206 (
      {stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449], stage0_28[450]},
      {stage0_29[71]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[74],stage1_30[86],stage1_29[157],stage1_28[230]}
   );
   gpc615_5 gpc1207 (
      {stage0_28[451], stage0_28[452], stage0_28[453], stage0_28[454], stage0_28[455]},
      {stage0_29[72]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[75],stage1_30[87],stage1_29[158],stage1_28[231]}
   );
   gpc615_5 gpc1208 (
      {stage0_28[456], stage0_28[457], stage0_28[458], stage0_28[459], stage0_28[460]},
      {stage0_29[73]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[76],stage1_30[88],stage1_29[159],stage1_28[232]}
   );
   gpc615_5 gpc1209 (
      {stage0_28[461], stage0_28[462], stage0_28[463], stage0_28[464], stage0_28[465]},
      {stage0_29[74]},
      {stage0_30[420], stage0_30[421], stage0_30[422], stage0_30[423], stage0_30[424], stage0_30[425]},
      {stage1_32[70],stage1_31[77],stage1_30[89],stage1_29[160],stage1_28[233]}
   );
   gpc615_5 gpc1210 (
      {stage0_28[466], stage0_28[467], stage0_28[468], stage0_28[469], stage0_28[470]},
      {stage0_29[75]},
      {stage0_30[426], stage0_30[427], stage0_30[428], stage0_30[429], stage0_30[430], stage0_30[431]},
      {stage1_32[71],stage1_31[78],stage1_30[90],stage1_29[161],stage1_28[234]}
   );
   gpc615_5 gpc1211 (
      {stage0_28[471], stage0_28[472], stage0_28[473], stage0_28[474], stage0_28[475]},
      {stage0_29[76]},
      {stage0_30[432], stage0_30[433], stage0_30[434], stage0_30[435], stage0_30[436], stage0_30[437]},
      {stage1_32[72],stage1_31[79],stage1_30[91],stage1_29[162],stage1_28[235]}
   );
   gpc615_5 gpc1212 (
      {stage0_28[476], stage0_28[477], stage0_28[478], stage0_28[479], stage0_28[480]},
      {stage0_29[77]},
      {stage0_30[438], stage0_30[439], stage0_30[440], stage0_30[441], stage0_30[442], stage0_30[443]},
      {stage1_32[73],stage1_31[80],stage1_30[92],stage1_29[163],stage1_28[236]}
   );
   gpc615_5 gpc1213 (
      {stage0_28[481], stage0_28[482], stage0_28[483], stage0_28[484], stage0_28[485]},
      {stage0_29[78]},
      {stage0_30[444], stage0_30[445], stage0_30[446], stage0_30[447], stage0_30[448], stage0_30[449]},
      {stage1_32[74],stage1_31[81],stage1_30[93],stage1_29[164],stage1_28[237]}
   );
   gpc615_5 gpc1214 (
      {stage0_28[486], stage0_28[487], stage0_28[488], stage0_28[489], stage0_28[490]},
      {stage0_29[79]},
      {stage0_30[450], stage0_30[451], stage0_30[452], stage0_30[453], stage0_30[454], stage0_30[455]},
      {stage1_32[75],stage1_31[82],stage1_30[94],stage1_29[165],stage1_28[238]}
   );
   gpc615_5 gpc1215 (
      {stage0_28[491], stage0_28[492], stage0_28[493], stage0_28[494], stage0_28[495]},
      {stage0_29[80]},
      {stage0_30[456], stage0_30[457], stage0_30[458], stage0_30[459], stage0_30[460], stage0_30[461]},
      {stage1_32[76],stage1_31[83],stage1_30[95],stage1_29[166],stage1_28[239]}
   );
   gpc615_5 gpc1216 (
      {stage0_28[496], stage0_28[497], stage0_28[498], stage0_28[499], stage0_28[500]},
      {stage0_29[81]},
      {stage0_30[462], stage0_30[463], stage0_30[464], stage0_30[465], stage0_30[466], stage0_30[467]},
      {stage1_32[77],stage1_31[84],stage1_30[96],stage1_29[167],stage1_28[240]}
   );
   gpc615_5 gpc1217 (
      {stage0_28[501], stage0_28[502], stage0_28[503], stage0_28[504], stage0_28[505]},
      {stage0_29[82]},
      {stage0_30[468], stage0_30[469], stage0_30[470], stage0_30[471], stage0_30[472], stage0_30[473]},
      {stage1_32[78],stage1_31[85],stage1_30[97],stage1_29[168],stage1_28[241]}
   );
   gpc606_5 gpc1218 (
      {stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[79],stage1_31[86],stage1_30[98],stage1_29[169]}
   );
   gpc606_5 gpc1219 (
      {stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[80],stage1_31[87],stage1_30[99],stage1_29[170]}
   );
   gpc606_5 gpc1220 (
      {stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[81],stage1_31[88],stage1_30[100],stage1_29[171]}
   );
   gpc606_5 gpc1221 (
      {stage0_29[101], stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[82],stage1_31[89],stage1_30[101],stage1_29[172]}
   );
   gpc606_5 gpc1222 (
      {stage0_29[107], stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[83],stage1_31[90],stage1_30[102],stage1_29[173]}
   );
   gpc606_5 gpc1223 (
      {stage0_29[113], stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[84],stage1_31[91],stage1_30[103],stage1_29[174]}
   );
   gpc606_5 gpc1224 (
      {stage0_29[119], stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[85],stage1_31[92],stage1_30[104],stage1_29[175]}
   );
   gpc606_5 gpc1225 (
      {stage0_29[125], stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[86],stage1_31[93],stage1_30[105],stage1_29[176]}
   );
   gpc606_5 gpc1226 (
      {stage0_29[131], stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[87],stage1_31[94],stage1_30[106],stage1_29[177]}
   );
   gpc606_5 gpc1227 (
      {stage0_29[137], stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[88],stage1_31[95],stage1_30[107],stage1_29[178]}
   );
   gpc606_5 gpc1228 (
      {stage0_29[143], stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[89],stage1_31[96],stage1_30[108],stage1_29[179]}
   );
   gpc606_5 gpc1229 (
      {stage0_29[149], stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[90],stage1_31[97],stage1_30[109],stage1_29[180]}
   );
   gpc606_5 gpc1230 (
      {stage0_29[155], stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[91],stage1_31[98],stage1_30[110],stage1_29[181]}
   );
   gpc606_5 gpc1231 (
      {stage0_29[161], stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[92],stage1_31[99],stage1_30[111],stage1_29[182]}
   );
   gpc606_5 gpc1232 (
      {stage0_29[167], stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[93],stage1_31[100],stage1_30[112],stage1_29[183]}
   );
   gpc606_5 gpc1233 (
      {stage0_29[173], stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[94],stage1_31[101],stage1_30[113],stage1_29[184]}
   );
   gpc606_5 gpc1234 (
      {stage0_29[179], stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[95],stage1_31[102],stage1_30[114],stage1_29[185]}
   );
   gpc606_5 gpc1235 (
      {stage0_29[185], stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[96],stage1_31[103],stage1_30[115],stage1_29[186]}
   );
   gpc606_5 gpc1236 (
      {stage0_29[191], stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[97],stage1_31[104],stage1_30[116],stage1_29[187]}
   );
   gpc606_5 gpc1237 (
      {stage0_29[197], stage0_29[198], stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[98],stage1_31[105],stage1_30[117],stage1_29[188]}
   );
   gpc606_5 gpc1238 (
      {stage0_29[203], stage0_29[204], stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[99],stage1_31[106],stage1_30[118],stage1_29[189]}
   );
   gpc606_5 gpc1239 (
      {stage0_29[209], stage0_29[210], stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[100],stage1_31[107],stage1_30[119],stage1_29[190]}
   );
   gpc606_5 gpc1240 (
      {stage0_29[215], stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[101],stage1_31[108],stage1_30[120],stage1_29[191]}
   );
   gpc606_5 gpc1241 (
      {stage0_29[221], stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[102],stage1_31[109],stage1_30[121],stage1_29[192]}
   );
   gpc606_5 gpc1242 (
      {stage0_29[227], stage0_29[228], stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[103],stage1_31[110],stage1_30[122],stage1_29[193]}
   );
   gpc606_5 gpc1243 (
      {stage0_29[233], stage0_29[234], stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[104],stage1_31[111],stage1_30[123],stage1_29[194]}
   );
   gpc606_5 gpc1244 (
      {stage0_29[239], stage0_29[240], stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[105],stage1_31[112],stage1_30[124],stage1_29[195]}
   );
   gpc606_5 gpc1245 (
      {stage0_29[245], stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[106],stage1_31[113],stage1_30[125],stage1_29[196]}
   );
   gpc606_5 gpc1246 (
      {stage0_29[251], stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255], stage0_29[256]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[107],stage1_31[114],stage1_30[126],stage1_29[197]}
   );
   gpc606_5 gpc1247 (
      {stage0_29[257], stage0_29[258], stage0_29[259], stage0_29[260], stage0_29[261], stage0_29[262]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[108],stage1_31[115],stage1_30[127],stage1_29[198]}
   );
   gpc606_5 gpc1248 (
      {stage0_29[263], stage0_29[264], stage0_29[265], stage0_29[266], stage0_29[267], stage0_29[268]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[109],stage1_31[116],stage1_30[128],stage1_29[199]}
   );
   gpc606_5 gpc1249 (
      {stage0_29[269], stage0_29[270], stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[110],stage1_31[117],stage1_30[129],stage1_29[200]}
   );
   gpc606_5 gpc1250 (
      {stage0_29[275], stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[111],stage1_31[118],stage1_30[130],stage1_29[201]}
   );
   gpc606_5 gpc1251 (
      {stage0_29[281], stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285], stage0_29[286]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[112],stage1_31[119],stage1_30[131],stage1_29[202]}
   );
   gpc606_5 gpc1252 (
      {stage0_29[287], stage0_29[288], stage0_29[289], stage0_29[290], stage0_29[291], stage0_29[292]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[113],stage1_31[120],stage1_30[132],stage1_29[203]}
   );
   gpc606_5 gpc1253 (
      {stage0_29[293], stage0_29[294], stage0_29[295], stage0_29[296], stage0_29[297], stage0_29[298]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[114],stage1_31[121],stage1_30[133],stage1_29[204]}
   );
   gpc606_5 gpc1254 (
      {stage0_29[299], stage0_29[300], stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[115],stage1_31[122],stage1_30[134],stage1_29[205]}
   );
   gpc606_5 gpc1255 (
      {stage0_29[305], stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[116],stage1_31[123],stage1_30[135],stage1_29[206]}
   );
   gpc606_5 gpc1256 (
      {stage0_29[311], stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315], stage0_29[316]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[117],stage1_31[124],stage1_30[136],stage1_29[207]}
   );
   gpc606_5 gpc1257 (
      {stage0_29[317], stage0_29[318], stage0_29[319], stage0_29[320], stage0_29[321], stage0_29[322]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[118],stage1_31[125],stage1_30[137],stage1_29[208]}
   );
   gpc606_5 gpc1258 (
      {stage0_29[323], stage0_29[324], stage0_29[325], stage0_29[326], stage0_29[327], stage0_29[328]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[119],stage1_31[126],stage1_30[138],stage1_29[209]}
   );
   gpc606_5 gpc1259 (
      {stage0_29[329], stage0_29[330], stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[120],stage1_31[127],stage1_30[139],stage1_29[210]}
   );
   gpc606_5 gpc1260 (
      {stage0_29[335], stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[121],stage1_31[128],stage1_30[140],stage1_29[211]}
   );
   gpc606_5 gpc1261 (
      {stage0_29[341], stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345], stage0_29[346]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[122],stage1_31[129],stage1_30[141],stage1_29[212]}
   );
   gpc606_5 gpc1262 (
      {stage0_29[347], stage0_29[348], stage0_29[349], stage0_29[350], stage0_29[351], stage0_29[352]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[123],stage1_31[130],stage1_30[142],stage1_29[213]}
   );
   gpc606_5 gpc1263 (
      {stage0_29[353], stage0_29[354], stage0_29[355], stage0_29[356], stage0_29[357], stage0_29[358]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[124],stage1_31[131],stage1_30[143],stage1_29[214]}
   );
   gpc606_5 gpc1264 (
      {stage0_29[359], stage0_29[360], stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[125],stage1_31[132],stage1_30[144],stage1_29[215]}
   );
   gpc606_5 gpc1265 (
      {stage0_29[365], stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[126],stage1_31[133],stage1_30[145],stage1_29[216]}
   );
   gpc606_5 gpc1266 (
      {stage0_29[371], stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375], stage0_29[376]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[127],stage1_31[134],stage1_30[146],stage1_29[217]}
   );
   gpc606_5 gpc1267 (
      {stage0_29[377], stage0_29[378], stage0_29[379], stage0_29[380], stage0_29[381], stage0_29[382]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[128],stage1_31[135],stage1_30[147],stage1_29[218]}
   );
   gpc606_5 gpc1268 (
      {stage0_29[383], stage0_29[384], stage0_29[385], stage0_29[386], stage0_29[387], stage0_29[388]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[129],stage1_31[136],stage1_30[148],stage1_29[219]}
   );
   gpc606_5 gpc1269 (
      {stage0_29[389], stage0_29[390], stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[130],stage1_31[137],stage1_30[149],stage1_29[220]}
   );
   gpc606_5 gpc1270 (
      {stage0_29[395], stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[131],stage1_31[138],stage1_30[150],stage1_29[221]}
   );
   gpc606_5 gpc1271 (
      {stage0_29[401], stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405], stage0_29[406]},
      {stage0_31[318], stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage1_33[53],stage1_32[132],stage1_31[139],stage1_30[151],stage1_29[222]}
   );
   gpc606_5 gpc1272 (
      {stage0_29[407], stage0_29[408], stage0_29[409], stage0_29[410], stage0_29[411], stage0_29[412]},
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329]},
      {stage1_33[54],stage1_32[133],stage1_31[140],stage1_30[152],stage1_29[223]}
   );
   gpc606_5 gpc1273 (
      {stage0_29[413], stage0_29[414], stage0_29[415], stage0_29[416], stage0_29[417], stage0_29[418]},
      {stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage1_33[55],stage1_32[134],stage1_31[141],stage1_30[153],stage1_29[224]}
   );
   gpc606_5 gpc1274 (
      {stage0_29[419], stage0_29[420], stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424]},
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340], stage0_31[341]},
      {stage1_33[56],stage1_32[135],stage1_31[142],stage1_30[154],stage1_29[225]}
   );
   gpc606_5 gpc1275 (
      {stage0_29[425], stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430]},
      {stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347]},
      {stage1_33[57],stage1_32[136],stage1_31[143],stage1_30[155],stage1_29[226]}
   );
   gpc606_5 gpc1276 (
      {stage0_29[431], stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435], stage0_29[436]},
      {stage0_31[348], stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage1_33[58],stage1_32[137],stage1_31[144],stage1_30[156],stage1_29[227]}
   );
   gpc606_5 gpc1277 (
      {stage0_29[437], stage0_29[438], stage0_29[439], stage0_29[440], stage0_29[441], stage0_29[442]},
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359]},
      {stage1_33[59],stage1_32[138],stage1_31[145],stage1_30[157],stage1_29[228]}
   );
   gpc606_5 gpc1278 (
      {stage0_29[443], stage0_29[444], stage0_29[445], stage0_29[446], stage0_29[447], stage0_29[448]},
      {stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage1_33[60],stage1_32[139],stage1_31[146],stage1_30[158],stage1_29[229]}
   );
   gpc606_5 gpc1279 (
      {stage0_29[449], stage0_29[450], stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454]},
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370], stage0_31[371]},
      {stage1_33[61],stage1_32[140],stage1_31[147],stage1_30[159],stage1_29[230]}
   );
   gpc606_5 gpc1280 (
      {stage0_29[455], stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460]},
      {stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377]},
      {stage1_33[62],stage1_32[141],stage1_31[148],stage1_30[160],stage1_29[231]}
   );
   gpc606_5 gpc1281 (
      {stage0_29[461], stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465], stage0_29[466]},
      {stage0_31[378], stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage1_33[63],stage1_32[142],stage1_31[149],stage1_30[161],stage1_29[232]}
   );
   gpc606_5 gpc1282 (
      {stage0_29[467], stage0_29[468], stage0_29[469], stage0_29[470], stage0_29[471], stage0_29[472]},
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389]},
      {stage1_33[64],stage1_32[143],stage1_31[150],stage1_30[162],stage1_29[233]}
   );
   gpc606_5 gpc1283 (
      {stage0_29[473], stage0_29[474], stage0_29[475], stage0_29[476], stage0_29[477], stage0_29[478]},
      {stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage1_33[65],stage1_32[144],stage1_31[151],stage1_30[163],stage1_29[234]}
   );
   gpc606_5 gpc1284 (
      {stage0_29[479], stage0_29[480], stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484]},
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400], stage0_31[401]},
      {stage1_33[66],stage1_32[145],stage1_31[152],stage1_30[164],stage1_29[235]}
   );
   gpc606_5 gpc1285 (
      {stage0_29[485], stage0_29[486], stage0_29[487], stage0_29[488], stage0_29[489], stage0_29[490]},
      {stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407]},
      {stage1_33[67],stage1_32[146],stage1_31[153],stage1_30[165],stage1_29[236]}
   );
   gpc606_5 gpc1286 (
      {stage0_29[491], stage0_29[492], stage0_29[493], stage0_29[494], stage0_29[495], stage0_29[496]},
      {stage0_31[408], stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage1_33[68],stage1_32[147],stage1_31[154],stage1_30[166],stage1_29[237]}
   );
   gpc606_5 gpc1287 (
      {stage0_29[497], stage0_29[498], stage0_29[499], stage0_29[500], stage0_29[501], stage0_29[502]},
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419]},
      {stage1_33[69],stage1_32[148],stage1_31[155],stage1_30[167],stage1_29[238]}
   );
   gpc606_5 gpc1288 (
      {stage0_29[503], stage0_29[504], stage0_29[505], stage0_29[506], stage0_29[507], stage0_29[508]},
      {stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage1_33[70],stage1_32[149],stage1_31[156],stage1_30[168],stage1_29[239]}
   );
   gpc1_1 gpc1289 (
      {stage0_0[502]},
      {stage1_0[101]}
   );
   gpc1_1 gpc1290 (
      {stage0_0[503]},
      {stage1_0[102]}
   );
   gpc1_1 gpc1291 (
      {stage0_0[504]},
      {stage1_0[103]}
   );
   gpc1_1 gpc1292 (
      {stage0_0[505]},
      {stage1_0[104]}
   );
   gpc1_1 gpc1293 (
      {stage0_0[506]},
      {stage1_0[105]}
   );
   gpc1_1 gpc1294 (
      {stage0_0[507]},
      {stage1_0[106]}
   );
   gpc1_1 gpc1295 (
      {stage0_0[508]},
      {stage1_0[107]}
   );
   gpc1_1 gpc1296 (
      {stage0_0[509]},
      {stage1_0[108]}
   );
   gpc1_1 gpc1297 (
      {stage0_0[510]},
      {stage1_0[109]}
   );
   gpc1_1 gpc1298 (
      {stage0_0[511]},
      {stage1_0[110]}
   );
   gpc1_1 gpc1299 (
      {stage0_1[453]},
      {stage1_1[140]}
   );
   gpc1_1 gpc1300 (
      {stage0_1[454]},
      {stage1_1[141]}
   );
   gpc1_1 gpc1301 (
      {stage0_1[455]},
      {stage1_1[142]}
   );
   gpc1_1 gpc1302 (
      {stage0_1[456]},
      {stage1_1[143]}
   );
   gpc1_1 gpc1303 (
      {stage0_1[457]},
      {stage1_1[144]}
   );
   gpc1_1 gpc1304 (
      {stage0_1[458]},
      {stage1_1[145]}
   );
   gpc1_1 gpc1305 (
      {stage0_1[459]},
      {stage1_1[146]}
   );
   gpc1_1 gpc1306 (
      {stage0_1[460]},
      {stage1_1[147]}
   );
   gpc1_1 gpc1307 (
      {stage0_1[461]},
      {stage1_1[148]}
   );
   gpc1_1 gpc1308 (
      {stage0_1[462]},
      {stage1_1[149]}
   );
   gpc1_1 gpc1309 (
      {stage0_1[463]},
      {stage1_1[150]}
   );
   gpc1_1 gpc1310 (
      {stage0_1[464]},
      {stage1_1[151]}
   );
   gpc1_1 gpc1311 (
      {stage0_1[465]},
      {stage1_1[152]}
   );
   gpc1_1 gpc1312 (
      {stage0_1[466]},
      {stage1_1[153]}
   );
   gpc1_1 gpc1313 (
      {stage0_1[467]},
      {stage1_1[154]}
   );
   gpc1_1 gpc1314 (
      {stage0_1[468]},
      {stage1_1[155]}
   );
   gpc1_1 gpc1315 (
      {stage0_1[469]},
      {stage1_1[156]}
   );
   gpc1_1 gpc1316 (
      {stage0_1[470]},
      {stage1_1[157]}
   );
   gpc1_1 gpc1317 (
      {stage0_1[471]},
      {stage1_1[158]}
   );
   gpc1_1 gpc1318 (
      {stage0_1[472]},
      {stage1_1[159]}
   );
   gpc1_1 gpc1319 (
      {stage0_1[473]},
      {stage1_1[160]}
   );
   gpc1_1 gpc1320 (
      {stage0_1[474]},
      {stage1_1[161]}
   );
   gpc1_1 gpc1321 (
      {stage0_1[475]},
      {stage1_1[162]}
   );
   gpc1_1 gpc1322 (
      {stage0_1[476]},
      {stage1_1[163]}
   );
   gpc1_1 gpc1323 (
      {stage0_1[477]},
      {stage1_1[164]}
   );
   gpc1_1 gpc1324 (
      {stage0_1[478]},
      {stage1_1[165]}
   );
   gpc1_1 gpc1325 (
      {stage0_1[479]},
      {stage1_1[166]}
   );
   gpc1_1 gpc1326 (
      {stage0_1[480]},
      {stage1_1[167]}
   );
   gpc1_1 gpc1327 (
      {stage0_1[481]},
      {stage1_1[168]}
   );
   gpc1_1 gpc1328 (
      {stage0_1[482]},
      {stage1_1[169]}
   );
   gpc1_1 gpc1329 (
      {stage0_1[483]},
      {stage1_1[170]}
   );
   gpc1_1 gpc1330 (
      {stage0_1[484]},
      {stage1_1[171]}
   );
   gpc1_1 gpc1331 (
      {stage0_1[485]},
      {stage1_1[172]}
   );
   gpc1_1 gpc1332 (
      {stage0_1[486]},
      {stage1_1[173]}
   );
   gpc1_1 gpc1333 (
      {stage0_1[487]},
      {stage1_1[174]}
   );
   gpc1_1 gpc1334 (
      {stage0_1[488]},
      {stage1_1[175]}
   );
   gpc1_1 gpc1335 (
      {stage0_1[489]},
      {stage1_1[176]}
   );
   gpc1_1 gpc1336 (
      {stage0_1[490]},
      {stage1_1[177]}
   );
   gpc1_1 gpc1337 (
      {stage0_1[491]},
      {stage1_1[178]}
   );
   gpc1_1 gpc1338 (
      {stage0_1[492]},
      {stage1_1[179]}
   );
   gpc1_1 gpc1339 (
      {stage0_1[493]},
      {stage1_1[180]}
   );
   gpc1_1 gpc1340 (
      {stage0_1[494]},
      {stage1_1[181]}
   );
   gpc1_1 gpc1341 (
      {stage0_1[495]},
      {stage1_1[182]}
   );
   gpc1_1 gpc1342 (
      {stage0_1[496]},
      {stage1_1[183]}
   );
   gpc1_1 gpc1343 (
      {stage0_1[497]},
      {stage1_1[184]}
   );
   gpc1_1 gpc1344 (
      {stage0_1[498]},
      {stage1_1[185]}
   );
   gpc1_1 gpc1345 (
      {stage0_1[499]},
      {stage1_1[186]}
   );
   gpc1_1 gpc1346 (
      {stage0_1[500]},
      {stage1_1[187]}
   );
   gpc1_1 gpc1347 (
      {stage0_1[501]},
      {stage1_1[188]}
   );
   gpc1_1 gpc1348 (
      {stage0_1[502]},
      {stage1_1[189]}
   );
   gpc1_1 gpc1349 (
      {stage0_1[503]},
      {stage1_1[190]}
   );
   gpc1_1 gpc1350 (
      {stage0_1[504]},
      {stage1_1[191]}
   );
   gpc1_1 gpc1351 (
      {stage0_1[505]},
      {stage1_1[192]}
   );
   gpc1_1 gpc1352 (
      {stage0_1[506]},
      {stage1_1[193]}
   );
   gpc1_1 gpc1353 (
      {stage0_1[507]},
      {stage1_1[194]}
   );
   gpc1_1 gpc1354 (
      {stage0_1[508]},
      {stage1_1[195]}
   );
   gpc1_1 gpc1355 (
      {stage0_1[509]},
      {stage1_1[196]}
   );
   gpc1_1 gpc1356 (
      {stage0_1[510]},
      {stage1_1[197]}
   );
   gpc1_1 gpc1357 (
      {stage0_1[511]},
      {stage1_1[198]}
   );
   gpc1_1 gpc1358 (
      {stage0_2[481]},
      {stage1_2[157]}
   );
   gpc1_1 gpc1359 (
      {stage0_2[482]},
      {stage1_2[158]}
   );
   gpc1_1 gpc1360 (
      {stage0_2[483]},
      {stage1_2[159]}
   );
   gpc1_1 gpc1361 (
      {stage0_2[484]},
      {stage1_2[160]}
   );
   gpc1_1 gpc1362 (
      {stage0_2[485]},
      {stage1_2[161]}
   );
   gpc1_1 gpc1363 (
      {stage0_2[486]},
      {stage1_2[162]}
   );
   gpc1_1 gpc1364 (
      {stage0_2[487]},
      {stage1_2[163]}
   );
   gpc1_1 gpc1365 (
      {stage0_2[488]},
      {stage1_2[164]}
   );
   gpc1_1 gpc1366 (
      {stage0_2[489]},
      {stage1_2[165]}
   );
   gpc1_1 gpc1367 (
      {stage0_2[490]},
      {stage1_2[166]}
   );
   gpc1_1 gpc1368 (
      {stage0_2[491]},
      {stage1_2[167]}
   );
   gpc1_1 gpc1369 (
      {stage0_2[492]},
      {stage1_2[168]}
   );
   gpc1_1 gpc1370 (
      {stage0_2[493]},
      {stage1_2[169]}
   );
   gpc1_1 gpc1371 (
      {stage0_2[494]},
      {stage1_2[170]}
   );
   gpc1_1 gpc1372 (
      {stage0_2[495]},
      {stage1_2[171]}
   );
   gpc1_1 gpc1373 (
      {stage0_2[496]},
      {stage1_2[172]}
   );
   gpc1_1 gpc1374 (
      {stage0_2[497]},
      {stage1_2[173]}
   );
   gpc1_1 gpc1375 (
      {stage0_2[498]},
      {stage1_2[174]}
   );
   gpc1_1 gpc1376 (
      {stage0_2[499]},
      {stage1_2[175]}
   );
   gpc1_1 gpc1377 (
      {stage0_2[500]},
      {stage1_2[176]}
   );
   gpc1_1 gpc1378 (
      {stage0_2[501]},
      {stage1_2[177]}
   );
   gpc1_1 gpc1379 (
      {stage0_2[502]},
      {stage1_2[178]}
   );
   gpc1_1 gpc1380 (
      {stage0_2[503]},
      {stage1_2[179]}
   );
   gpc1_1 gpc1381 (
      {stage0_2[504]},
      {stage1_2[180]}
   );
   gpc1_1 gpc1382 (
      {stage0_2[505]},
      {stage1_2[181]}
   );
   gpc1_1 gpc1383 (
      {stage0_2[506]},
      {stage1_2[182]}
   );
   gpc1_1 gpc1384 (
      {stage0_2[507]},
      {stage1_2[183]}
   );
   gpc1_1 gpc1385 (
      {stage0_2[508]},
      {stage1_2[184]}
   );
   gpc1_1 gpc1386 (
      {stage0_2[509]},
      {stage1_2[185]}
   );
   gpc1_1 gpc1387 (
      {stage0_2[510]},
      {stage1_2[186]}
   );
   gpc1_1 gpc1388 (
      {stage0_2[511]},
      {stage1_2[187]}
   );
   gpc1_1 gpc1389 (
      {stage0_3[414]},
      {stage1_3[179]}
   );
   gpc1_1 gpc1390 (
      {stage0_3[415]},
      {stage1_3[180]}
   );
   gpc1_1 gpc1391 (
      {stage0_3[416]},
      {stage1_3[181]}
   );
   gpc1_1 gpc1392 (
      {stage0_3[417]},
      {stage1_3[182]}
   );
   gpc1_1 gpc1393 (
      {stage0_3[418]},
      {stage1_3[183]}
   );
   gpc1_1 gpc1394 (
      {stage0_3[419]},
      {stage1_3[184]}
   );
   gpc1_1 gpc1395 (
      {stage0_3[420]},
      {stage1_3[185]}
   );
   gpc1_1 gpc1396 (
      {stage0_3[421]},
      {stage1_3[186]}
   );
   gpc1_1 gpc1397 (
      {stage0_3[422]},
      {stage1_3[187]}
   );
   gpc1_1 gpc1398 (
      {stage0_3[423]},
      {stage1_3[188]}
   );
   gpc1_1 gpc1399 (
      {stage0_3[424]},
      {stage1_3[189]}
   );
   gpc1_1 gpc1400 (
      {stage0_3[425]},
      {stage1_3[190]}
   );
   gpc1_1 gpc1401 (
      {stage0_3[426]},
      {stage1_3[191]}
   );
   gpc1_1 gpc1402 (
      {stage0_3[427]},
      {stage1_3[192]}
   );
   gpc1_1 gpc1403 (
      {stage0_3[428]},
      {stage1_3[193]}
   );
   gpc1_1 gpc1404 (
      {stage0_3[429]},
      {stage1_3[194]}
   );
   gpc1_1 gpc1405 (
      {stage0_3[430]},
      {stage1_3[195]}
   );
   gpc1_1 gpc1406 (
      {stage0_3[431]},
      {stage1_3[196]}
   );
   gpc1_1 gpc1407 (
      {stage0_3[432]},
      {stage1_3[197]}
   );
   gpc1_1 gpc1408 (
      {stage0_3[433]},
      {stage1_3[198]}
   );
   gpc1_1 gpc1409 (
      {stage0_3[434]},
      {stage1_3[199]}
   );
   gpc1_1 gpc1410 (
      {stage0_3[435]},
      {stage1_3[200]}
   );
   gpc1_1 gpc1411 (
      {stage0_3[436]},
      {stage1_3[201]}
   );
   gpc1_1 gpc1412 (
      {stage0_3[437]},
      {stage1_3[202]}
   );
   gpc1_1 gpc1413 (
      {stage0_3[438]},
      {stage1_3[203]}
   );
   gpc1_1 gpc1414 (
      {stage0_3[439]},
      {stage1_3[204]}
   );
   gpc1_1 gpc1415 (
      {stage0_3[440]},
      {stage1_3[205]}
   );
   gpc1_1 gpc1416 (
      {stage0_3[441]},
      {stage1_3[206]}
   );
   gpc1_1 gpc1417 (
      {stage0_3[442]},
      {stage1_3[207]}
   );
   gpc1_1 gpc1418 (
      {stage0_3[443]},
      {stage1_3[208]}
   );
   gpc1_1 gpc1419 (
      {stage0_3[444]},
      {stage1_3[209]}
   );
   gpc1_1 gpc1420 (
      {stage0_3[445]},
      {stage1_3[210]}
   );
   gpc1_1 gpc1421 (
      {stage0_3[446]},
      {stage1_3[211]}
   );
   gpc1_1 gpc1422 (
      {stage0_3[447]},
      {stage1_3[212]}
   );
   gpc1_1 gpc1423 (
      {stage0_3[448]},
      {stage1_3[213]}
   );
   gpc1_1 gpc1424 (
      {stage0_3[449]},
      {stage1_3[214]}
   );
   gpc1_1 gpc1425 (
      {stage0_3[450]},
      {stage1_3[215]}
   );
   gpc1_1 gpc1426 (
      {stage0_3[451]},
      {stage1_3[216]}
   );
   gpc1_1 gpc1427 (
      {stage0_3[452]},
      {stage1_3[217]}
   );
   gpc1_1 gpc1428 (
      {stage0_3[453]},
      {stage1_3[218]}
   );
   gpc1_1 gpc1429 (
      {stage0_3[454]},
      {stage1_3[219]}
   );
   gpc1_1 gpc1430 (
      {stage0_3[455]},
      {stage1_3[220]}
   );
   gpc1_1 gpc1431 (
      {stage0_3[456]},
      {stage1_3[221]}
   );
   gpc1_1 gpc1432 (
      {stage0_3[457]},
      {stage1_3[222]}
   );
   gpc1_1 gpc1433 (
      {stage0_3[458]},
      {stage1_3[223]}
   );
   gpc1_1 gpc1434 (
      {stage0_3[459]},
      {stage1_3[224]}
   );
   gpc1_1 gpc1435 (
      {stage0_3[460]},
      {stage1_3[225]}
   );
   gpc1_1 gpc1436 (
      {stage0_3[461]},
      {stage1_3[226]}
   );
   gpc1_1 gpc1437 (
      {stage0_3[462]},
      {stage1_3[227]}
   );
   gpc1_1 gpc1438 (
      {stage0_3[463]},
      {stage1_3[228]}
   );
   gpc1_1 gpc1439 (
      {stage0_3[464]},
      {stage1_3[229]}
   );
   gpc1_1 gpc1440 (
      {stage0_3[465]},
      {stage1_3[230]}
   );
   gpc1_1 gpc1441 (
      {stage0_3[466]},
      {stage1_3[231]}
   );
   gpc1_1 gpc1442 (
      {stage0_3[467]},
      {stage1_3[232]}
   );
   gpc1_1 gpc1443 (
      {stage0_3[468]},
      {stage1_3[233]}
   );
   gpc1_1 gpc1444 (
      {stage0_3[469]},
      {stage1_3[234]}
   );
   gpc1_1 gpc1445 (
      {stage0_3[470]},
      {stage1_3[235]}
   );
   gpc1_1 gpc1446 (
      {stage0_3[471]},
      {stage1_3[236]}
   );
   gpc1_1 gpc1447 (
      {stage0_3[472]},
      {stage1_3[237]}
   );
   gpc1_1 gpc1448 (
      {stage0_3[473]},
      {stage1_3[238]}
   );
   gpc1_1 gpc1449 (
      {stage0_3[474]},
      {stage1_3[239]}
   );
   gpc1_1 gpc1450 (
      {stage0_3[475]},
      {stage1_3[240]}
   );
   gpc1_1 gpc1451 (
      {stage0_3[476]},
      {stage1_3[241]}
   );
   gpc1_1 gpc1452 (
      {stage0_3[477]},
      {stage1_3[242]}
   );
   gpc1_1 gpc1453 (
      {stage0_3[478]},
      {stage1_3[243]}
   );
   gpc1_1 gpc1454 (
      {stage0_3[479]},
      {stage1_3[244]}
   );
   gpc1_1 gpc1455 (
      {stage0_3[480]},
      {stage1_3[245]}
   );
   gpc1_1 gpc1456 (
      {stage0_3[481]},
      {stage1_3[246]}
   );
   gpc1_1 gpc1457 (
      {stage0_3[482]},
      {stage1_3[247]}
   );
   gpc1_1 gpc1458 (
      {stage0_3[483]},
      {stage1_3[248]}
   );
   gpc1_1 gpc1459 (
      {stage0_3[484]},
      {stage1_3[249]}
   );
   gpc1_1 gpc1460 (
      {stage0_3[485]},
      {stage1_3[250]}
   );
   gpc1_1 gpc1461 (
      {stage0_3[486]},
      {stage1_3[251]}
   );
   gpc1_1 gpc1462 (
      {stage0_3[487]},
      {stage1_3[252]}
   );
   gpc1_1 gpc1463 (
      {stage0_3[488]},
      {stage1_3[253]}
   );
   gpc1_1 gpc1464 (
      {stage0_3[489]},
      {stage1_3[254]}
   );
   gpc1_1 gpc1465 (
      {stage0_3[490]},
      {stage1_3[255]}
   );
   gpc1_1 gpc1466 (
      {stage0_3[491]},
      {stage1_3[256]}
   );
   gpc1_1 gpc1467 (
      {stage0_3[492]},
      {stage1_3[257]}
   );
   gpc1_1 gpc1468 (
      {stage0_3[493]},
      {stage1_3[258]}
   );
   gpc1_1 gpc1469 (
      {stage0_3[494]},
      {stage1_3[259]}
   );
   gpc1_1 gpc1470 (
      {stage0_3[495]},
      {stage1_3[260]}
   );
   gpc1_1 gpc1471 (
      {stage0_3[496]},
      {stage1_3[261]}
   );
   gpc1_1 gpc1472 (
      {stage0_3[497]},
      {stage1_3[262]}
   );
   gpc1_1 gpc1473 (
      {stage0_3[498]},
      {stage1_3[263]}
   );
   gpc1_1 gpc1474 (
      {stage0_3[499]},
      {stage1_3[264]}
   );
   gpc1_1 gpc1475 (
      {stage0_3[500]},
      {stage1_3[265]}
   );
   gpc1_1 gpc1476 (
      {stage0_3[501]},
      {stage1_3[266]}
   );
   gpc1_1 gpc1477 (
      {stage0_3[502]},
      {stage1_3[267]}
   );
   gpc1_1 gpc1478 (
      {stage0_3[503]},
      {stage1_3[268]}
   );
   gpc1_1 gpc1479 (
      {stage0_3[504]},
      {stage1_3[269]}
   );
   gpc1_1 gpc1480 (
      {stage0_3[505]},
      {stage1_3[270]}
   );
   gpc1_1 gpc1481 (
      {stage0_3[506]},
      {stage1_3[271]}
   );
   gpc1_1 gpc1482 (
      {stage0_3[507]},
      {stage1_3[272]}
   );
   gpc1_1 gpc1483 (
      {stage0_3[508]},
      {stage1_3[273]}
   );
   gpc1_1 gpc1484 (
      {stage0_3[509]},
      {stage1_3[274]}
   );
   gpc1_1 gpc1485 (
      {stage0_3[510]},
      {stage1_3[275]}
   );
   gpc1_1 gpc1486 (
      {stage0_3[511]},
      {stage1_3[276]}
   );
   gpc1_1 gpc1487 (
      {stage0_6[446]},
      {stage1_6[177]}
   );
   gpc1_1 gpc1488 (
      {stage0_6[447]},
      {stage1_6[178]}
   );
   gpc1_1 gpc1489 (
      {stage0_6[448]},
      {stage1_6[179]}
   );
   gpc1_1 gpc1490 (
      {stage0_6[449]},
      {stage1_6[180]}
   );
   gpc1_1 gpc1491 (
      {stage0_6[450]},
      {stage1_6[181]}
   );
   gpc1_1 gpc1492 (
      {stage0_6[451]},
      {stage1_6[182]}
   );
   gpc1_1 gpc1493 (
      {stage0_6[452]},
      {stage1_6[183]}
   );
   gpc1_1 gpc1494 (
      {stage0_6[453]},
      {stage1_6[184]}
   );
   gpc1_1 gpc1495 (
      {stage0_6[454]},
      {stage1_6[185]}
   );
   gpc1_1 gpc1496 (
      {stage0_6[455]},
      {stage1_6[186]}
   );
   gpc1_1 gpc1497 (
      {stage0_6[456]},
      {stage1_6[187]}
   );
   gpc1_1 gpc1498 (
      {stage0_6[457]},
      {stage1_6[188]}
   );
   gpc1_1 gpc1499 (
      {stage0_6[458]},
      {stage1_6[189]}
   );
   gpc1_1 gpc1500 (
      {stage0_6[459]},
      {stage1_6[190]}
   );
   gpc1_1 gpc1501 (
      {stage0_6[460]},
      {stage1_6[191]}
   );
   gpc1_1 gpc1502 (
      {stage0_6[461]},
      {stage1_6[192]}
   );
   gpc1_1 gpc1503 (
      {stage0_6[462]},
      {stage1_6[193]}
   );
   gpc1_1 gpc1504 (
      {stage0_6[463]},
      {stage1_6[194]}
   );
   gpc1_1 gpc1505 (
      {stage0_6[464]},
      {stage1_6[195]}
   );
   gpc1_1 gpc1506 (
      {stage0_6[465]},
      {stage1_6[196]}
   );
   gpc1_1 gpc1507 (
      {stage0_6[466]},
      {stage1_6[197]}
   );
   gpc1_1 gpc1508 (
      {stage0_6[467]},
      {stage1_6[198]}
   );
   gpc1_1 gpc1509 (
      {stage0_6[468]},
      {stage1_6[199]}
   );
   gpc1_1 gpc1510 (
      {stage0_6[469]},
      {stage1_6[200]}
   );
   gpc1_1 gpc1511 (
      {stage0_6[470]},
      {stage1_6[201]}
   );
   gpc1_1 gpc1512 (
      {stage0_6[471]},
      {stage1_6[202]}
   );
   gpc1_1 gpc1513 (
      {stage0_6[472]},
      {stage1_6[203]}
   );
   gpc1_1 gpc1514 (
      {stage0_6[473]},
      {stage1_6[204]}
   );
   gpc1_1 gpc1515 (
      {stage0_6[474]},
      {stage1_6[205]}
   );
   gpc1_1 gpc1516 (
      {stage0_6[475]},
      {stage1_6[206]}
   );
   gpc1_1 gpc1517 (
      {stage0_6[476]},
      {stage1_6[207]}
   );
   gpc1_1 gpc1518 (
      {stage0_6[477]},
      {stage1_6[208]}
   );
   gpc1_1 gpc1519 (
      {stage0_6[478]},
      {stage1_6[209]}
   );
   gpc1_1 gpc1520 (
      {stage0_6[479]},
      {stage1_6[210]}
   );
   gpc1_1 gpc1521 (
      {stage0_6[480]},
      {stage1_6[211]}
   );
   gpc1_1 gpc1522 (
      {stage0_6[481]},
      {stage1_6[212]}
   );
   gpc1_1 gpc1523 (
      {stage0_6[482]},
      {stage1_6[213]}
   );
   gpc1_1 gpc1524 (
      {stage0_6[483]},
      {stage1_6[214]}
   );
   gpc1_1 gpc1525 (
      {stage0_6[484]},
      {stage1_6[215]}
   );
   gpc1_1 gpc1526 (
      {stage0_6[485]},
      {stage1_6[216]}
   );
   gpc1_1 gpc1527 (
      {stage0_6[486]},
      {stage1_6[217]}
   );
   gpc1_1 gpc1528 (
      {stage0_6[487]},
      {stage1_6[218]}
   );
   gpc1_1 gpc1529 (
      {stage0_6[488]},
      {stage1_6[219]}
   );
   gpc1_1 gpc1530 (
      {stage0_6[489]},
      {stage1_6[220]}
   );
   gpc1_1 gpc1531 (
      {stage0_6[490]},
      {stage1_6[221]}
   );
   gpc1_1 gpc1532 (
      {stage0_6[491]},
      {stage1_6[222]}
   );
   gpc1_1 gpc1533 (
      {stage0_6[492]},
      {stage1_6[223]}
   );
   gpc1_1 gpc1534 (
      {stage0_6[493]},
      {stage1_6[224]}
   );
   gpc1_1 gpc1535 (
      {stage0_6[494]},
      {stage1_6[225]}
   );
   gpc1_1 gpc1536 (
      {stage0_6[495]},
      {stage1_6[226]}
   );
   gpc1_1 gpc1537 (
      {stage0_6[496]},
      {stage1_6[227]}
   );
   gpc1_1 gpc1538 (
      {stage0_6[497]},
      {stage1_6[228]}
   );
   gpc1_1 gpc1539 (
      {stage0_6[498]},
      {stage1_6[229]}
   );
   gpc1_1 gpc1540 (
      {stage0_6[499]},
      {stage1_6[230]}
   );
   gpc1_1 gpc1541 (
      {stage0_6[500]},
      {stage1_6[231]}
   );
   gpc1_1 gpc1542 (
      {stage0_6[501]},
      {stage1_6[232]}
   );
   gpc1_1 gpc1543 (
      {stage0_6[502]},
      {stage1_6[233]}
   );
   gpc1_1 gpc1544 (
      {stage0_6[503]},
      {stage1_6[234]}
   );
   gpc1_1 gpc1545 (
      {stage0_6[504]},
      {stage1_6[235]}
   );
   gpc1_1 gpc1546 (
      {stage0_6[505]},
      {stage1_6[236]}
   );
   gpc1_1 gpc1547 (
      {stage0_6[506]},
      {stage1_6[237]}
   );
   gpc1_1 gpc1548 (
      {stage0_6[507]},
      {stage1_6[238]}
   );
   gpc1_1 gpc1549 (
      {stage0_6[508]},
      {stage1_6[239]}
   );
   gpc1_1 gpc1550 (
      {stage0_6[509]},
      {stage1_6[240]}
   );
   gpc1_1 gpc1551 (
      {stage0_6[510]},
      {stage1_6[241]}
   );
   gpc1_1 gpc1552 (
      {stage0_6[511]},
      {stage1_6[242]}
   );
   gpc1_1 gpc1553 (
      {stage0_8[377]},
      {stage1_8[214]}
   );
   gpc1_1 gpc1554 (
      {stage0_8[378]},
      {stage1_8[215]}
   );
   gpc1_1 gpc1555 (
      {stage0_8[379]},
      {stage1_8[216]}
   );
   gpc1_1 gpc1556 (
      {stage0_8[380]},
      {stage1_8[217]}
   );
   gpc1_1 gpc1557 (
      {stage0_8[381]},
      {stage1_8[218]}
   );
   gpc1_1 gpc1558 (
      {stage0_8[382]},
      {stage1_8[219]}
   );
   gpc1_1 gpc1559 (
      {stage0_8[383]},
      {stage1_8[220]}
   );
   gpc1_1 gpc1560 (
      {stage0_8[384]},
      {stage1_8[221]}
   );
   gpc1_1 gpc1561 (
      {stage0_8[385]},
      {stage1_8[222]}
   );
   gpc1_1 gpc1562 (
      {stage0_8[386]},
      {stage1_8[223]}
   );
   gpc1_1 gpc1563 (
      {stage0_8[387]},
      {stage1_8[224]}
   );
   gpc1_1 gpc1564 (
      {stage0_8[388]},
      {stage1_8[225]}
   );
   gpc1_1 gpc1565 (
      {stage0_8[389]},
      {stage1_8[226]}
   );
   gpc1_1 gpc1566 (
      {stage0_8[390]},
      {stage1_8[227]}
   );
   gpc1_1 gpc1567 (
      {stage0_8[391]},
      {stage1_8[228]}
   );
   gpc1_1 gpc1568 (
      {stage0_8[392]},
      {stage1_8[229]}
   );
   gpc1_1 gpc1569 (
      {stage0_8[393]},
      {stage1_8[230]}
   );
   gpc1_1 gpc1570 (
      {stage0_8[394]},
      {stage1_8[231]}
   );
   gpc1_1 gpc1571 (
      {stage0_8[395]},
      {stage1_8[232]}
   );
   gpc1_1 gpc1572 (
      {stage0_8[396]},
      {stage1_8[233]}
   );
   gpc1_1 gpc1573 (
      {stage0_8[397]},
      {stage1_8[234]}
   );
   gpc1_1 gpc1574 (
      {stage0_8[398]},
      {stage1_8[235]}
   );
   gpc1_1 gpc1575 (
      {stage0_8[399]},
      {stage1_8[236]}
   );
   gpc1_1 gpc1576 (
      {stage0_8[400]},
      {stage1_8[237]}
   );
   gpc1_1 gpc1577 (
      {stage0_8[401]},
      {stage1_8[238]}
   );
   gpc1_1 gpc1578 (
      {stage0_8[402]},
      {stage1_8[239]}
   );
   gpc1_1 gpc1579 (
      {stage0_8[403]},
      {stage1_8[240]}
   );
   gpc1_1 gpc1580 (
      {stage0_8[404]},
      {stage1_8[241]}
   );
   gpc1_1 gpc1581 (
      {stage0_8[405]},
      {stage1_8[242]}
   );
   gpc1_1 gpc1582 (
      {stage0_8[406]},
      {stage1_8[243]}
   );
   gpc1_1 gpc1583 (
      {stage0_8[407]},
      {stage1_8[244]}
   );
   gpc1_1 gpc1584 (
      {stage0_8[408]},
      {stage1_8[245]}
   );
   gpc1_1 gpc1585 (
      {stage0_8[409]},
      {stage1_8[246]}
   );
   gpc1_1 gpc1586 (
      {stage0_8[410]},
      {stage1_8[247]}
   );
   gpc1_1 gpc1587 (
      {stage0_8[411]},
      {stage1_8[248]}
   );
   gpc1_1 gpc1588 (
      {stage0_8[412]},
      {stage1_8[249]}
   );
   gpc1_1 gpc1589 (
      {stage0_8[413]},
      {stage1_8[250]}
   );
   gpc1_1 gpc1590 (
      {stage0_8[414]},
      {stage1_8[251]}
   );
   gpc1_1 gpc1591 (
      {stage0_8[415]},
      {stage1_8[252]}
   );
   gpc1_1 gpc1592 (
      {stage0_8[416]},
      {stage1_8[253]}
   );
   gpc1_1 gpc1593 (
      {stage0_8[417]},
      {stage1_8[254]}
   );
   gpc1_1 gpc1594 (
      {stage0_8[418]},
      {stage1_8[255]}
   );
   gpc1_1 gpc1595 (
      {stage0_8[419]},
      {stage1_8[256]}
   );
   gpc1_1 gpc1596 (
      {stage0_8[420]},
      {stage1_8[257]}
   );
   gpc1_1 gpc1597 (
      {stage0_8[421]},
      {stage1_8[258]}
   );
   gpc1_1 gpc1598 (
      {stage0_8[422]},
      {stage1_8[259]}
   );
   gpc1_1 gpc1599 (
      {stage0_8[423]},
      {stage1_8[260]}
   );
   gpc1_1 gpc1600 (
      {stage0_8[424]},
      {stage1_8[261]}
   );
   gpc1_1 gpc1601 (
      {stage0_8[425]},
      {stage1_8[262]}
   );
   gpc1_1 gpc1602 (
      {stage0_8[426]},
      {stage1_8[263]}
   );
   gpc1_1 gpc1603 (
      {stage0_8[427]},
      {stage1_8[264]}
   );
   gpc1_1 gpc1604 (
      {stage0_8[428]},
      {stage1_8[265]}
   );
   gpc1_1 gpc1605 (
      {stage0_8[429]},
      {stage1_8[266]}
   );
   gpc1_1 gpc1606 (
      {stage0_8[430]},
      {stage1_8[267]}
   );
   gpc1_1 gpc1607 (
      {stage0_8[431]},
      {stage1_8[268]}
   );
   gpc1_1 gpc1608 (
      {stage0_8[432]},
      {stage1_8[269]}
   );
   gpc1_1 gpc1609 (
      {stage0_8[433]},
      {stage1_8[270]}
   );
   gpc1_1 gpc1610 (
      {stage0_8[434]},
      {stage1_8[271]}
   );
   gpc1_1 gpc1611 (
      {stage0_8[435]},
      {stage1_8[272]}
   );
   gpc1_1 gpc1612 (
      {stage0_8[436]},
      {stage1_8[273]}
   );
   gpc1_1 gpc1613 (
      {stage0_8[437]},
      {stage1_8[274]}
   );
   gpc1_1 gpc1614 (
      {stage0_8[438]},
      {stage1_8[275]}
   );
   gpc1_1 gpc1615 (
      {stage0_8[439]},
      {stage1_8[276]}
   );
   gpc1_1 gpc1616 (
      {stage0_8[440]},
      {stage1_8[277]}
   );
   gpc1_1 gpc1617 (
      {stage0_8[441]},
      {stage1_8[278]}
   );
   gpc1_1 gpc1618 (
      {stage0_8[442]},
      {stage1_8[279]}
   );
   gpc1_1 gpc1619 (
      {stage0_8[443]},
      {stage1_8[280]}
   );
   gpc1_1 gpc1620 (
      {stage0_8[444]},
      {stage1_8[281]}
   );
   gpc1_1 gpc1621 (
      {stage0_8[445]},
      {stage1_8[282]}
   );
   gpc1_1 gpc1622 (
      {stage0_8[446]},
      {stage1_8[283]}
   );
   gpc1_1 gpc1623 (
      {stage0_8[447]},
      {stage1_8[284]}
   );
   gpc1_1 gpc1624 (
      {stage0_8[448]},
      {stage1_8[285]}
   );
   gpc1_1 gpc1625 (
      {stage0_8[449]},
      {stage1_8[286]}
   );
   gpc1_1 gpc1626 (
      {stage0_8[450]},
      {stage1_8[287]}
   );
   gpc1_1 gpc1627 (
      {stage0_8[451]},
      {stage1_8[288]}
   );
   gpc1_1 gpc1628 (
      {stage0_8[452]},
      {stage1_8[289]}
   );
   gpc1_1 gpc1629 (
      {stage0_8[453]},
      {stage1_8[290]}
   );
   gpc1_1 gpc1630 (
      {stage0_8[454]},
      {stage1_8[291]}
   );
   gpc1_1 gpc1631 (
      {stage0_8[455]},
      {stage1_8[292]}
   );
   gpc1_1 gpc1632 (
      {stage0_8[456]},
      {stage1_8[293]}
   );
   gpc1_1 gpc1633 (
      {stage0_8[457]},
      {stage1_8[294]}
   );
   gpc1_1 gpc1634 (
      {stage0_8[458]},
      {stage1_8[295]}
   );
   gpc1_1 gpc1635 (
      {stage0_8[459]},
      {stage1_8[296]}
   );
   gpc1_1 gpc1636 (
      {stage0_8[460]},
      {stage1_8[297]}
   );
   gpc1_1 gpc1637 (
      {stage0_8[461]},
      {stage1_8[298]}
   );
   gpc1_1 gpc1638 (
      {stage0_8[462]},
      {stage1_8[299]}
   );
   gpc1_1 gpc1639 (
      {stage0_8[463]},
      {stage1_8[300]}
   );
   gpc1_1 gpc1640 (
      {stage0_8[464]},
      {stage1_8[301]}
   );
   gpc1_1 gpc1641 (
      {stage0_8[465]},
      {stage1_8[302]}
   );
   gpc1_1 gpc1642 (
      {stage0_8[466]},
      {stage1_8[303]}
   );
   gpc1_1 gpc1643 (
      {stage0_8[467]},
      {stage1_8[304]}
   );
   gpc1_1 gpc1644 (
      {stage0_8[468]},
      {stage1_8[305]}
   );
   gpc1_1 gpc1645 (
      {stage0_8[469]},
      {stage1_8[306]}
   );
   gpc1_1 gpc1646 (
      {stage0_8[470]},
      {stage1_8[307]}
   );
   gpc1_1 gpc1647 (
      {stage0_8[471]},
      {stage1_8[308]}
   );
   gpc1_1 gpc1648 (
      {stage0_8[472]},
      {stage1_8[309]}
   );
   gpc1_1 gpc1649 (
      {stage0_8[473]},
      {stage1_8[310]}
   );
   gpc1_1 gpc1650 (
      {stage0_8[474]},
      {stage1_8[311]}
   );
   gpc1_1 gpc1651 (
      {stage0_8[475]},
      {stage1_8[312]}
   );
   gpc1_1 gpc1652 (
      {stage0_8[476]},
      {stage1_8[313]}
   );
   gpc1_1 gpc1653 (
      {stage0_8[477]},
      {stage1_8[314]}
   );
   gpc1_1 gpc1654 (
      {stage0_8[478]},
      {stage1_8[315]}
   );
   gpc1_1 gpc1655 (
      {stage0_8[479]},
      {stage1_8[316]}
   );
   gpc1_1 gpc1656 (
      {stage0_8[480]},
      {stage1_8[317]}
   );
   gpc1_1 gpc1657 (
      {stage0_8[481]},
      {stage1_8[318]}
   );
   gpc1_1 gpc1658 (
      {stage0_8[482]},
      {stage1_8[319]}
   );
   gpc1_1 gpc1659 (
      {stage0_8[483]},
      {stage1_8[320]}
   );
   gpc1_1 gpc1660 (
      {stage0_8[484]},
      {stage1_8[321]}
   );
   gpc1_1 gpc1661 (
      {stage0_8[485]},
      {stage1_8[322]}
   );
   gpc1_1 gpc1662 (
      {stage0_8[486]},
      {stage1_8[323]}
   );
   gpc1_1 gpc1663 (
      {stage0_8[487]},
      {stage1_8[324]}
   );
   gpc1_1 gpc1664 (
      {stage0_8[488]},
      {stage1_8[325]}
   );
   gpc1_1 gpc1665 (
      {stage0_8[489]},
      {stage1_8[326]}
   );
   gpc1_1 gpc1666 (
      {stage0_8[490]},
      {stage1_8[327]}
   );
   gpc1_1 gpc1667 (
      {stage0_8[491]},
      {stage1_8[328]}
   );
   gpc1_1 gpc1668 (
      {stage0_8[492]},
      {stage1_8[329]}
   );
   gpc1_1 gpc1669 (
      {stage0_8[493]},
      {stage1_8[330]}
   );
   gpc1_1 gpc1670 (
      {stage0_8[494]},
      {stage1_8[331]}
   );
   gpc1_1 gpc1671 (
      {stage0_8[495]},
      {stage1_8[332]}
   );
   gpc1_1 gpc1672 (
      {stage0_8[496]},
      {stage1_8[333]}
   );
   gpc1_1 gpc1673 (
      {stage0_8[497]},
      {stage1_8[334]}
   );
   gpc1_1 gpc1674 (
      {stage0_8[498]},
      {stage1_8[335]}
   );
   gpc1_1 gpc1675 (
      {stage0_8[499]},
      {stage1_8[336]}
   );
   gpc1_1 gpc1676 (
      {stage0_8[500]},
      {stage1_8[337]}
   );
   gpc1_1 gpc1677 (
      {stage0_8[501]},
      {stage1_8[338]}
   );
   gpc1_1 gpc1678 (
      {stage0_8[502]},
      {stage1_8[339]}
   );
   gpc1_1 gpc1679 (
      {stage0_8[503]},
      {stage1_8[340]}
   );
   gpc1_1 gpc1680 (
      {stage0_8[504]},
      {stage1_8[341]}
   );
   gpc1_1 gpc1681 (
      {stage0_8[505]},
      {stage1_8[342]}
   );
   gpc1_1 gpc1682 (
      {stage0_8[506]},
      {stage1_8[343]}
   );
   gpc1_1 gpc1683 (
      {stage0_8[507]},
      {stage1_8[344]}
   );
   gpc1_1 gpc1684 (
      {stage0_8[508]},
      {stage1_8[345]}
   );
   gpc1_1 gpc1685 (
      {stage0_8[509]},
      {stage1_8[346]}
   );
   gpc1_1 gpc1686 (
      {stage0_8[510]},
      {stage1_8[347]}
   );
   gpc1_1 gpc1687 (
      {stage0_8[511]},
      {stage1_8[348]}
   );
   gpc1_1 gpc1688 (
      {stage0_9[509]},
      {stage1_9[209]}
   );
   gpc1_1 gpc1689 (
      {stage0_9[510]},
      {stage1_9[210]}
   );
   gpc1_1 gpc1690 (
      {stage0_9[511]},
      {stage1_9[211]}
   );
   gpc1_1 gpc1691 (
      {stage0_11[501]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1692 (
      {stage0_11[502]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1693 (
      {stage0_11[503]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1694 (
      {stage0_11[504]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1695 (
      {stage0_11[505]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1696 (
      {stage0_11[506]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1697 (
      {stage0_11[507]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1698 (
      {stage0_11[508]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1699 (
      {stage0_11[509]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1700 (
      {stage0_11[510]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1701 (
      {stage0_11[511]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1702 (
      {stage0_13[507]},
      {stage1_13[227]}
   );
   gpc1_1 gpc1703 (
      {stage0_13[508]},
      {stage1_13[228]}
   );
   gpc1_1 gpc1704 (
      {stage0_13[509]},
      {stage1_13[229]}
   );
   gpc1_1 gpc1705 (
      {stage0_13[510]},
      {stage1_13[230]}
   );
   gpc1_1 gpc1706 (
      {stage0_13[511]},
      {stage1_13[231]}
   );
   gpc1_1 gpc1707 (
      {stage0_14[472]},
      {stage1_14[192]}
   );
   gpc1_1 gpc1708 (
      {stage0_14[473]},
      {stage1_14[193]}
   );
   gpc1_1 gpc1709 (
      {stage0_14[474]},
      {stage1_14[194]}
   );
   gpc1_1 gpc1710 (
      {stage0_14[475]},
      {stage1_14[195]}
   );
   gpc1_1 gpc1711 (
      {stage0_14[476]},
      {stage1_14[196]}
   );
   gpc1_1 gpc1712 (
      {stage0_14[477]},
      {stage1_14[197]}
   );
   gpc1_1 gpc1713 (
      {stage0_14[478]},
      {stage1_14[198]}
   );
   gpc1_1 gpc1714 (
      {stage0_14[479]},
      {stage1_14[199]}
   );
   gpc1_1 gpc1715 (
      {stage0_14[480]},
      {stage1_14[200]}
   );
   gpc1_1 gpc1716 (
      {stage0_14[481]},
      {stage1_14[201]}
   );
   gpc1_1 gpc1717 (
      {stage0_14[482]},
      {stage1_14[202]}
   );
   gpc1_1 gpc1718 (
      {stage0_14[483]},
      {stage1_14[203]}
   );
   gpc1_1 gpc1719 (
      {stage0_14[484]},
      {stage1_14[204]}
   );
   gpc1_1 gpc1720 (
      {stage0_14[485]},
      {stage1_14[205]}
   );
   gpc1_1 gpc1721 (
      {stage0_14[486]},
      {stage1_14[206]}
   );
   gpc1_1 gpc1722 (
      {stage0_14[487]},
      {stage1_14[207]}
   );
   gpc1_1 gpc1723 (
      {stage0_14[488]},
      {stage1_14[208]}
   );
   gpc1_1 gpc1724 (
      {stage0_14[489]},
      {stage1_14[209]}
   );
   gpc1_1 gpc1725 (
      {stage0_14[490]},
      {stage1_14[210]}
   );
   gpc1_1 gpc1726 (
      {stage0_14[491]},
      {stage1_14[211]}
   );
   gpc1_1 gpc1727 (
      {stage0_14[492]},
      {stage1_14[212]}
   );
   gpc1_1 gpc1728 (
      {stage0_14[493]},
      {stage1_14[213]}
   );
   gpc1_1 gpc1729 (
      {stage0_14[494]},
      {stage1_14[214]}
   );
   gpc1_1 gpc1730 (
      {stage0_14[495]},
      {stage1_14[215]}
   );
   gpc1_1 gpc1731 (
      {stage0_14[496]},
      {stage1_14[216]}
   );
   gpc1_1 gpc1732 (
      {stage0_14[497]},
      {stage1_14[217]}
   );
   gpc1_1 gpc1733 (
      {stage0_14[498]},
      {stage1_14[218]}
   );
   gpc1_1 gpc1734 (
      {stage0_14[499]},
      {stage1_14[219]}
   );
   gpc1_1 gpc1735 (
      {stage0_14[500]},
      {stage1_14[220]}
   );
   gpc1_1 gpc1736 (
      {stage0_14[501]},
      {stage1_14[221]}
   );
   gpc1_1 gpc1737 (
      {stage0_14[502]},
      {stage1_14[222]}
   );
   gpc1_1 gpc1738 (
      {stage0_14[503]},
      {stage1_14[223]}
   );
   gpc1_1 gpc1739 (
      {stage0_14[504]},
      {stage1_14[224]}
   );
   gpc1_1 gpc1740 (
      {stage0_14[505]},
      {stage1_14[225]}
   );
   gpc1_1 gpc1741 (
      {stage0_14[506]},
      {stage1_14[226]}
   );
   gpc1_1 gpc1742 (
      {stage0_14[507]},
      {stage1_14[227]}
   );
   gpc1_1 gpc1743 (
      {stage0_14[508]},
      {stage1_14[228]}
   );
   gpc1_1 gpc1744 (
      {stage0_14[509]},
      {stage1_14[229]}
   );
   gpc1_1 gpc1745 (
      {stage0_14[510]},
      {stage1_14[230]}
   );
   gpc1_1 gpc1746 (
      {stage0_14[511]},
      {stage1_14[231]}
   );
   gpc1_1 gpc1747 (
      {stage0_15[456]},
      {stage1_15[181]}
   );
   gpc1_1 gpc1748 (
      {stage0_15[457]},
      {stage1_15[182]}
   );
   gpc1_1 gpc1749 (
      {stage0_15[458]},
      {stage1_15[183]}
   );
   gpc1_1 gpc1750 (
      {stage0_15[459]},
      {stage1_15[184]}
   );
   gpc1_1 gpc1751 (
      {stage0_15[460]},
      {stage1_15[185]}
   );
   gpc1_1 gpc1752 (
      {stage0_15[461]},
      {stage1_15[186]}
   );
   gpc1_1 gpc1753 (
      {stage0_15[462]},
      {stage1_15[187]}
   );
   gpc1_1 gpc1754 (
      {stage0_15[463]},
      {stage1_15[188]}
   );
   gpc1_1 gpc1755 (
      {stage0_15[464]},
      {stage1_15[189]}
   );
   gpc1_1 gpc1756 (
      {stage0_15[465]},
      {stage1_15[190]}
   );
   gpc1_1 gpc1757 (
      {stage0_15[466]},
      {stage1_15[191]}
   );
   gpc1_1 gpc1758 (
      {stage0_15[467]},
      {stage1_15[192]}
   );
   gpc1_1 gpc1759 (
      {stage0_15[468]},
      {stage1_15[193]}
   );
   gpc1_1 gpc1760 (
      {stage0_15[469]},
      {stage1_15[194]}
   );
   gpc1_1 gpc1761 (
      {stage0_15[470]},
      {stage1_15[195]}
   );
   gpc1_1 gpc1762 (
      {stage0_15[471]},
      {stage1_15[196]}
   );
   gpc1_1 gpc1763 (
      {stage0_15[472]},
      {stage1_15[197]}
   );
   gpc1_1 gpc1764 (
      {stage0_15[473]},
      {stage1_15[198]}
   );
   gpc1_1 gpc1765 (
      {stage0_15[474]},
      {stage1_15[199]}
   );
   gpc1_1 gpc1766 (
      {stage0_15[475]},
      {stage1_15[200]}
   );
   gpc1_1 gpc1767 (
      {stage0_15[476]},
      {stage1_15[201]}
   );
   gpc1_1 gpc1768 (
      {stage0_15[477]},
      {stage1_15[202]}
   );
   gpc1_1 gpc1769 (
      {stage0_15[478]},
      {stage1_15[203]}
   );
   gpc1_1 gpc1770 (
      {stage0_15[479]},
      {stage1_15[204]}
   );
   gpc1_1 gpc1771 (
      {stage0_15[480]},
      {stage1_15[205]}
   );
   gpc1_1 gpc1772 (
      {stage0_15[481]},
      {stage1_15[206]}
   );
   gpc1_1 gpc1773 (
      {stage0_15[482]},
      {stage1_15[207]}
   );
   gpc1_1 gpc1774 (
      {stage0_15[483]},
      {stage1_15[208]}
   );
   gpc1_1 gpc1775 (
      {stage0_15[484]},
      {stage1_15[209]}
   );
   gpc1_1 gpc1776 (
      {stage0_15[485]},
      {stage1_15[210]}
   );
   gpc1_1 gpc1777 (
      {stage0_15[486]},
      {stage1_15[211]}
   );
   gpc1_1 gpc1778 (
      {stage0_15[487]},
      {stage1_15[212]}
   );
   gpc1_1 gpc1779 (
      {stage0_15[488]},
      {stage1_15[213]}
   );
   gpc1_1 gpc1780 (
      {stage0_15[489]},
      {stage1_15[214]}
   );
   gpc1_1 gpc1781 (
      {stage0_15[490]},
      {stage1_15[215]}
   );
   gpc1_1 gpc1782 (
      {stage0_15[491]},
      {stage1_15[216]}
   );
   gpc1_1 gpc1783 (
      {stage0_15[492]},
      {stage1_15[217]}
   );
   gpc1_1 gpc1784 (
      {stage0_15[493]},
      {stage1_15[218]}
   );
   gpc1_1 gpc1785 (
      {stage0_15[494]},
      {stage1_15[219]}
   );
   gpc1_1 gpc1786 (
      {stage0_15[495]},
      {stage1_15[220]}
   );
   gpc1_1 gpc1787 (
      {stage0_15[496]},
      {stage1_15[221]}
   );
   gpc1_1 gpc1788 (
      {stage0_15[497]},
      {stage1_15[222]}
   );
   gpc1_1 gpc1789 (
      {stage0_15[498]},
      {stage1_15[223]}
   );
   gpc1_1 gpc1790 (
      {stage0_15[499]},
      {stage1_15[224]}
   );
   gpc1_1 gpc1791 (
      {stage0_15[500]},
      {stage1_15[225]}
   );
   gpc1_1 gpc1792 (
      {stage0_15[501]},
      {stage1_15[226]}
   );
   gpc1_1 gpc1793 (
      {stage0_15[502]},
      {stage1_15[227]}
   );
   gpc1_1 gpc1794 (
      {stage0_15[503]},
      {stage1_15[228]}
   );
   gpc1_1 gpc1795 (
      {stage0_15[504]},
      {stage1_15[229]}
   );
   gpc1_1 gpc1796 (
      {stage0_15[505]},
      {stage1_15[230]}
   );
   gpc1_1 gpc1797 (
      {stage0_15[506]},
      {stage1_15[231]}
   );
   gpc1_1 gpc1798 (
      {stage0_15[507]},
      {stage1_15[232]}
   );
   gpc1_1 gpc1799 (
      {stage0_15[508]},
      {stage1_15[233]}
   );
   gpc1_1 gpc1800 (
      {stage0_15[509]},
      {stage1_15[234]}
   );
   gpc1_1 gpc1801 (
      {stage0_15[510]},
      {stage1_15[235]}
   );
   gpc1_1 gpc1802 (
      {stage0_15[511]},
      {stage1_15[236]}
   );
   gpc1_1 gpc1803 (
      {stage0_17[510]},
      {stage1_17[222]}
   );
   gpc1_1 gpc1804 (
      {stage0_17[511]},
      {stage1_17[223]}
   );
   gpc1_1 gpc1805 (
      {stage0_18[511]},
      {stage1_18[202]}
   );
   gpc1_1 gpc1806 (
      {stage0_19[431]},
      {stage1_19[182]}
   );
   gpc1_1 gpc1807 (
      {stage0_19[432]},
      {stage1_19[183]}
   );
   gpc1_1 gpc1808 (
      {stage0_19[433]},
      {stage1_19[184]}
   );
   gpc1_1 gpc1809 (
      {stage0_19[434]},
      {stage1_19[185]}
   );
   gpc1_1 gpc1810 (
      {stage0_19[435]},
      {stage1_19[186]}
   );
   gpc1_1 gpc1811 (
      {stage0_19[436]},
      {stage1_19[187]}
   );
   gpc1_1 gpc1812 (
      {stage0_19[437]},
      {stage1_19[188]}
   );
   gpc1_1 gpc1813 (
      {stage0_19[438]},
      {stage1_19[189]}
   );
   gpc1_1 gpc1814 (
      {stage0_19[439]},
      {stage1_19[190]}
   );
   gpc1_1 gpc1815 (
      {stage0_19[440]},
      {stage1_19[191]}
   );
   gpc1_1 gpc1816 (
      {stage0_19[441]},
      {stage1_19[192]}
   );
   gpc1_1 gpc1817 (
      {stage0_19[442]},
      {stage1_19[193]}
   );
   gpc1_1 gpc1818 (
      {stage0_19[443]},
      {stage1_19[194]}
   );
   gpc1_1 gpc1819 (
      {stage0_19[444]},
      {stage1_19[195]}
   );
   gpc1_1 gpc1820 (
      {stage0_19[445]},
      {stage1_19[196]}
   );
   gpc1_1 gpc1821 (
      {stage0_19[446]},
      {stage1_19[197]}
   );
   gpc1_1 gpc1822 (
      {stage0_19[447]},
      {stage1_19[198]}
   );
   gpc1_1 gpc1823 (
      {stage0_19[448]},
      {stage1_19[199]}
   );
   gpc1_1 gpc1824 (
      {stage0_19[449]},
      {stage1_19[200]}
   );
   gpc1_1 gpc1825 (
      {stage0_19[450]},
      {stage1_19[201]}
   );
   gpc1_1 gpc1826 (
      {stage0_19[451]},
      {stage1_19[202]}
   );
   gpc1_1 gpc1827 (
      {stage0_19[452]},
      {stage1_19[203]}
   );
   gpc1_1 gpc1828 (
      {stage0_19[453]},
      {stage1_19[204]}
   );
   gpc1_1 gpc1829 (
      {stage0_19[454]},
      {stage1_19[205]}
   );
   gpc1_1 gpc1830 (
      {stage0_19[455]},
      {stage1_19[206]}
   );
   gpc1_1 gpc1831 (
      {stage0_19[456]},
      {stage1_19[207]}
   );
   gpc1_1 gpc1832 (
      {stage0_19[457]},
      {stage1_19[208]}
   );
   gpc1_1 gpc1833 (
      {stage0_19[458]},
      {stage1_19[209]}
   );
   gpc1_1 gpc1834 (
      {stage0_19[459]},
      {stage1_19[210]}
   );
   gpc1_1 gpc1835 (
      {stage0_19[460]},
      {stage1_19[211]}
   );
   gpc1_1 gpc1836 (
      {stage0_19[461]},
      {stage1_19[212]}
   );
   gpc1_1 gpc1837 (
      {stage0_19[462]},
      {stage1_19[213]}
   );
   gpc1_1 gpc1838 (
      {stage0_19[463]},
      {stage1_19[214]}
   );
   gpc1_1 gpc1839 (
      {stage0_19[464]},
      {stage1_19[215]}
   );
   gpc1_1 gpc1840 (
      {stage0_19[465]},
      {stage1_19[216]}
   );
   gpc1_1 gpc1841 (
      {stage0_19[466]},
      {stage1_19[217]}
   );
   gpc1_1 gpc1842 (
      {stage0_19[467]},
      {stage1_19[218]}
   );
   gpc1_1 gpc1843 (
      {stage0_19[468]},
      {stage1_19[219]}
   );
   gpc1_1 gpc1844 (
      {stage0_19[469]},
      {stage1_19[220]}
   );
   gpc1_1 gpc1845 (
      {stage0_19[470]},
      {stage1_19[221]}
   );
   gpc1_1 gpc1846 (
      {stage0_19[471]},
      {stage1_19[222]}
   );
   gpc1_1 gpc1847 (
      {stage0_19[472]},
      {stage1_19[223]}
   );
   gpc1_1 gpc1848 (
      {stage0_19[473]},
      {stage1_19[224]}
   );
   gpc1_1 gpc1849 (
      {stage0_19[474]},
      {stage1_19[225]}
   );
   gpc1_1 gpc1850 (
      {stage0_19[475]},
      {stage1_19[226]}
   );
   gpc1_1 gpc1851 (
      {stage0_19[476]},
      {stage1_19[227]}
   );
   gpc1_1 gpc1852 (
      {stage0_19[477]},
      {stage1_19[228]}
   );
   gpc1_1 gpc1853 (
      {stage0_19[478]},
      {stage1_19[229]}
   );
   gpc1_1 gpc1854 (
      {stage0_19[479]},
      {stage1_19[230]}
   );
   gpc1_1 gpc1855 (
      {stage0_19[480]},
      {stage1_19[231]}
   );
   gpc1_1 gpc1856 (
      {stage0_19[481]},
      {stage1_19[232]}
   );
   gpc1_1 gpc1857 (
      {stage0_19[482]},
      {stage1_19[233]}
   );
   gpc1_1 gpc1858 (
      {stage0_19[483]},
      {stage1_19[234]}
   );
   gpc1_1 gpc1859 (
      {stage0_19[484]},
      {stage1_19[235]}
   );
   gpc1_1 gpc1860 (
      {stage0_19[485]},
      {stage1_19[236]}
   );
   gpc1_1 gpc1861 (
      {stage0_19[486]},
      {stage1_19[237]}
   );
   gpc1_1 gpc1862 (
      {stage0_19[487]},
      {stage1_19[238]}
   );
   gpc1_1 gpc1863 (
      {stage0_19[488]},
      {stage1_19[239]}
   );
   gpc1_1 gpc1864 (
      {stage0_19[489]},
      {stage1_19[240]}
   );
   gpc1_1 gpc1865 (
      {stage0_19[490]},
      {stage1_19[241]}
   );
   gpc1_1 gpc1866 (
      {stage0_19[491]},
      {stage1_19[242]}
   );
   gpc1_1 gpc1867 (
      {stage0_19[492]},
      {stage1_19[243]}
   );
   gpc1_1 gpc1868 (
      {stage0_19[493]},
      {stage1_19[244]}
   );
   gpc1_1 gpc1869 (
      {stage0_19[494]},
      {stage1_19[245]}
   );
   gpc1_1 gpc1870 (
      {stage0_19[495]},
      {stage1_19[246]}
   );
   gpc1_1 gpc1871 (
      {stage0_19[496]},
      {stage1_19[247]}
   );
   gpc1_1 gpc1872 (
      {stage0_19[497]},
      {stage1_19[248]}
   );
   gpc1_1 gpc1873 (
      {stage0_19[498]},
      {stage1_19[249]}
   );
   gpc1_1 gpc1874 (
      {stage0_19[499]},
      {stage1_19[250]}
   );
   gpc1_1 gpc1875 (
      {stage0_19[500]},
      {stage1_19[251]}
   );
   gpc1_1 gpc1876 (
      {stage0_19[501]},
      {stage1_19[252]}
   );
   gpc1_1 gpc1877 (
      {stage0_19[502]},
      {stage1_19[253]}
   );
   gpc1_1 gpc1878 (
      {stage0_19[503]},
      {stage1_19[254]}
   );
   gpc1_1 gpc1879 (
      {stage0_19[504]},
      {stage1_19[255]}
   );
   gpc1_1 gpc1880 (
      {stage0_19[505]},
      {stage1_19[256]}
   );
   gpc1_1 gpc1881 (
      {stage0_19[506]},
      {stage1_19[257]}
   );
   gpc1_1 gpc1882 (
      {stage0_19[507]},
      {stage1_19[258]}
   );
   gpc1_1 gpc1883 (
      {stage0_19[508]},
      {stage1_19[259]}
   );
   gpc1_1 gpc1884 (
      {stage0_19[509]},
      {stage1_19[260]}
   );
   gpc1_1 gpc1885 (
      {stage0_19[510]},
      {stage1_19[261]}
   );
   gpc1_1 gpc1886 (
      {stage0_19[511]},
      {stage1_19[262]}
   );
   gpc1_1 gpc1887 (
      {stage0_20[504]},
      {stage1_20[206]}
   );
   gpc1_1 gpc1888 (
      {stage0_20[505]},
      {stage1_20[207]}
   );
   gpc1_1 gpc1889 (
      {stage0_20[506]},
      {stage1_20[208]}
   );
   gpc1_1 gpc1890 (
      {stage0_20[507]},
      {stage1_20[209]}
   );
   gpc1_1 gpc1891 (
      {stage0_20[508]},
      {stage1_20[210]}
   );
   gpc1_1 gpc1892 (
      {stage0_20[509]},
      {stage1_20[211]}
   );
   gpc1_1 gpc1893 (
      {stage0_20[510]},
      {stage1_20[212]}
   );
   gpc1_1 gpc1894 (
      {stage0_20[511]},
      {stage1_20[213]}
   );
   gpc1_1 gpc1895 (
      {stage0_21[471]},
      {stage1_21[229]}
   );
   gpc1_1 gpc1896 (
      {stage0_21[472]},
      {stage1_21[230]}
   );
   gpc1_1 gpc1897 (
      {stage0_21[473]},
      {stage1_21[231]}
   );
   gpc1_1 gpc1898 (
      {stage0_21[474]},
      {stage1_21[232]}
   );
   gpc1_1 gpc1899 (
      {stage0_21[475]},
      {stage1_21[233]}
   );
   gpc1_1 gpc1900 (
      {stage0_21[476]},
      {stage1_21[234]}
   );
   gpc1_1 gpc1901 (
      {stage0_21[477]},
      {stage1_21[235]}
   );
   gpc1_1 gpc1902 (
      {stage0_21[478]},
      {stage1_21[236]}
   );
   gpc1_1 gpc1903 (
      {stage0_21[479]},
      {stage1_21[237]}
   );
   gpc1_1 gpc1904 (
      {stage0_21[480]},
      {stage1_21[238]}
   );
   gpc1_1 gpc1905 (
      {stage0_21[481]},
      {stage1_21[239]}
   );
   gpc1_1 gpc1906 (
      {stage0_21[482]},
      {stage1_21[240]}
   );
   gpc1_1 gpc1907 (
      {stage0_21[483]},
      {stage1_21[241]}
   );
   gpc1_1 gpc1908 (
      {stage0_21[484]},
      {stage1_21[242]}
   );
   gpc1_1 gpc1909 (
      {stage0_21[485]},
      {stage1_21[243]}
   );
   gpc1_1 gpc1910 (
      {stage0_21[486]},
      {stage1_21[244]}
   );
   gpc1_1 gpc1911 (
      {stage0_21[487]},
      {stage1_21[245]}
   );
   gpc1_1 gpc1912 (
      {stage0_21[488]},
      {stage1_21[246]}
   );
   gpc1_1 gpc1913 (
      {stage0_21[489]},
      {stage1_21[247]}
   );
   gpc1_1 gpc1914 (
      {stage0_21[490]},
      {stage1_21[248]}
   );
   gpc1_1 gpc1915 (
      {stage0_21[491]},
      {stage1_21[249]}
   );
   gpc1_1 gpc1916 (
      {stage0_21[492]},
      {stage1_21[250]}
   );
   gpc1_1 gpc1917 (
      {stage0_21[493]},
      {stage1_21[251]}
   );
   gpc1_1 gpc1918 (
      {stage0_21[494]},
      {stage1_21[252]}
   );
   gpc1_1 gpc1919 (
      {stage0_21[495]},
      {stage1_21[253]}
   );
   gpc1_1 gpc1920 (
      {stage0_21[496]},
      {stage1_21[254]}
   );
   gpc1_1 gpc1921 (
      {stage0_21[497]},
      {stage1_21[255]}
   );
   gpc1_1 gpc1922 (
      {stage0_21[498]},
      {stage1_21[256]}
   );
   gpc1_1 gpc1923 (
      {stage0_21[499]},
      {stage1_21[257]}
   );
   gpc1_1 gpc1924 (
      {stage0_21[500]},
      {stage1_21[258]}
   );
   gpc1_1 gpc1925 (
      {stage0_21[501]},
      {stage1_21[259]}
   );
   gpc1_1 gpc1926 (
      {stage0_21[502]},
      {stage1_21[260]}
   );
   gpc1_1 gpc1927 (
      {stage0_21[503]},
      {stage1_21[261]}
   );
   gpc1_1 gpc1928 (
      {stage0_21[504]},
      {stage1_21[262]}
   );
   gpc1_1 gpc1929 (
      {stage0_21[505]},
      {stage1_21[263]}
   );
   gpc1_1 gpc1930 (
      {stage0_21[506]},
      {stage1_21[264]}
   );
   gpc1_1 gpc1931 (
      {stage0_21[507]},
      {stage1_21[265]}
   );
   gpc1_1 gpc1932 (
      {stage0_21[508]},
      {stage1_21[266]}
   );
   gpc1_1 gpc1933 (
      {stage0_21[509]},
      {stage1_21[267]}
   );
   gpc1_1 gpc1934 (
      {stage0_21[510]},
      {stage1_21[268]}
   );
   gpc1_1 gpc1935 (
      {stage0_21[511]},
      {stage1_21[269]}
   );
   gpc1_1 gpc1936 (
      {stage0_22[423]},
      {stage1_22[185]}
   );
   gpc1_1 gpc1937 (
      {stage0_22[424]},
      {stage1_22[186]}
   );
   gpc1_1 gpc1938 (
      {stage0_22[425]},
      {stage1_22[187]}
   );
   gpc1_1 gpc1939 (
      {stage0_22[426]},
      {stage1_22[188]}
   );
   gpc1_1 gpc1940 (
      {stage0_22[427]},
      {stage1_22[189]}
   );
   gpc1_1 gpc1941 (
      {stage0_22[428]},
      {stage1_22[190]}
   );
   gpc1_1 gpc1942 (
      {stage0_22[429]},
      {stage1_22[191]}
   );
   gpc1_1 gpc1943 (
      {stage0_22[430]},
      {stage1_22[192]}
   );
   gpc1_1 gpc1944 (
      {stage0_22[431]},
      {stage1_22[193]}
   );
   gpc1_1 gpc1945 (
      {stage0_22[432]},
      {stage1_22[194]}
   );
   gpc1_1 gpc1946 (
      {stage0_22[433]},
      {stage1_22[195]}
   );
   gpc1_1 gpc1947 (
      {stage0_22[434]},
      {stage1_22[196]}
   );
   gpc1_1 gpc1948 (
      {stage0_22[435]},
      {stage1_22[197]}
   );
   gpc1_1 gpc1949 (
      {stage0_22[436]},
      {stage1_22[198]}
   );
   gpc1_1 gpc1950 (
      {stage0_22[437]},
      {stage1_22[199]}
   );
   gpc1_1 gpc1951 (
      {stage0_22[438]},
      {stage1_22[200]}
   );
   gpc1_1 gpc1952 (
      {stage0_22[439]},
      {stage1_22[201]}
   );
   gpc1_1 gpc1953 (
      {stage0_22[440]},
      {stage1_22[202]}
   );
   gpc1_1 gpc1954 (
      {stage0_22[441]},
      {stage1_22[203]}
   );
   gpc1_1 gpc1955 (
      {stage0_22[442]},
      {stage1_22[204]}
   );
   gpc1_1 gpc1956 (
      {stage0_22[443]},
      {stage1_22[205]}
   );
   gpc1_1 gpc1957 (
      {stage0_22[444]},
      {stage1_22[206]}
   );
   gpc1_1 gpc1958 (
      {stage0_22[445]},
      {stage1_22[207]}
   );
   gpc1_1 gpc1959 (
      {stage0_22[446]},
      {stage1_22[208]}
   );
   gpc1_1 gpc1960 (
      {stage0_22[447]},
      {stage1_22[209]}
   );
   gpc1_1 gpc1961 (
      {stage0_22[448]},
      {stage1_22[210]}
   );
   gpc1_1 gpc1962 (
      {stage0_22[449]},
      {stage1_22[211]}
   );
   gpc1_1 gpc1963 (
      {stage0_22[450]},
      {stage1_22[212]}
   );
   gpc1_1 gpc1964 (
      {stage0_22[451]},
      {stage1_22[213]}
   );
   gpc1_1 gpc1965 (
      {stage0_22[452]},
      {stage1_22[214]}
   );
   gpc1_1 gpc1966 (
      {stage0_22[453]},
      {stage1_22[215]}
   );
   gpc1_1 gpc1967 (
      {stage0_22[454]},
      {stage1_22[216]}
   );
   gpc1_1 gpc1968 (
      {stage0_22[455]},
      {stage1_22[217]}
   );
   gpc1_1 gpc1969 (
      {stage0_22[456]},
      {stage1_22[218]}
   );
   gpc1_1 gpc1970 (
      {stage0_22[457]},
      {stage1_22[219]}
   );
   gpc1_1 gpc1971 (
      {stage0_22[458]},
      {stage1_22[220]}
   );
   gpc1_1 gpc1972 (
      {stage0_22[459]},
      {stage1_22[221]}
   );
   gpc1_1 gpc1973 (
      {stage0_22[460]},
      {stage1_22[222]}
   );
   gpc1_1 gpc1974 (
      {stage0_22[461]},
      {stage1_22[223]}
   );
   gpc1_1 gpc1975 (
      {stage0_22[462]},
      {stage1_22[224]}
   );
   gpc1_1 gpc1976 (
      {stage0_22[463]},
      {stage1_22[225]}
   );
   gpc1_1 gpc1977 (
      {stage0_22[464]},
      {stage1_22[226]}
   );
   gpc1_1 gpc1978 (
      {stage0_22[465]},
      {stage1_22[227]}
   );
   gpc1_1 gpc1979 (
      {stage0_22[466]},
      {stage1_22[228]}
   );
   gpc1_1 gpc1980 (
      {stage0_22[467]},
      {stage1_22[229]}
   );
   gpc1_1 gpc1981 (
      {stage0_22[468]},
      {stage1_22[230]}
   );
   gpc1_1 gpc1982 (
      {stage0_22[469]},
      {stage1_22[231]}
   );
   gpc1_1 gpc1983 (
      {stage0_22[470]},
      {stage1_22[232]}
   );
   gpc1_1 gpc1984 (
      {stage0_22[471]},
      {stage1_22[233]}
   );
   gpc1_1 gpc1985 (
      {stage0_22[472]},
      {stage1_22[234]}
   );
   gpc1_1 gpc1986 (
      {stage0_22[473]},
      {stage1_22[235]}
   );
   gpc1_1 gpc1987 (
      {stage0_22[474]},
      {stage1_22[236]}
   );
   gpc1_1 gpc1988 (
      {stage0_22[475]},
      {stage1_22[237]}
   );
   gpc1_1 gpc1989 (
      {stage0_22[476]},
      {stage1_22[238]}
   );
   gpc1_1 gpc1990 (
      {stage0_22[477]},
      {stage1_22[239]}
   );
   gpc1_1 gpc1991 (
      {stage0_22[478]},
      {stage1_22[240]}
   );
   gpc1_1 gpc1992 (
      {stage0_22[479]},
      {stage1_22[241]}
   );
   gpc1_1 gpc1993 (
      {stage0_22[480]},
      {stage1_22[242]}
   );
   gpc1_1 gpc1994 (
      {stage0_22[481]},
      {stage1_22[243]}
   );
   gpc1_1 gpc1995 (
      {stage0_22[482]},
      {stage1_22[244]}
   );
   gpc1_1 gpc1996 (
      {stage0_22[483]},
      {stage1_22[245]}
   );
   gpc1_1 gpc1997 (
      {stage0_22[484]},
      {stage1_22[246]}
   );
   gpc1_1 gpc1998 (
      {stage0_22[485]},
      {stage1_22[247]}
   );
   gpc1_1 gpc1999 (
      {stage0_22[486]},
      {stage1_22[248]}
   );
   gpc1_1 gpc2000 (
      {stage0_22[487]},
      {stage1_22[249]}
   );
   gpc1_1 gpc2001 (
      {stage0_22[488]},
      {stage1_22[250]}
   );
   gpc1_1 gpc2002 (
      {stage0_22[489]},
      {stage1_22[251]}
   );
   gpc1_1 gpc2003 (
      {stage0_22[490]},
      {stage1_22[252]}
   );
   gpc1_1 gpc2004 (
      {stage0_22[491]},
      {stage1_22[253]}
   );
   gpc1_1 gpc2005 (
      {stage0_22[492]},
      {stage1_22[254]}
   );
   gpc1_1 gpc2006 (
      {stage0_22[493]},
      {stage1_22[255]}
   );
   gpc1_1 gpc2007 (
      {stage0_22[494]},
      {stage1_22[256]}
   );
   gpc1_1 gpc2008 (
      {stage0_22[495]},
      {stage1_22[257]}
   );
   gpc1_1 gpc2009 (
      {stage0_22[496]},
      {stage1_22[258]}
   );
   gpc1_1 gpc2010 (
      {stage0_22[497]},
      {stage1_22[259]}
   );
   gpc1_1 gpc2011 (
      {stage0_22[498]},
      {stage1_22[260]}
   );
   gpc1_1 gpc2012 (
      {stage0_22[499]},
      {stage1_22[261]}
   );
   gpc1_1 gpc2013 (
      {stage0_22[500]},
      {stage1_22[262]}
   );
   gpc1_1 gpc2014 (
      {stage0_22[501]},
      {stage1_22[263]}
   );
   gpc1_1 gpc2015 (
      {stage0_22[502]},
      {stage1_22[264]}
   );
   gpc1_1 gpc2016 (
      {stage0_22[503]},
      {stage1_22[265]}
   );
   gpc1_1 gpc2017 (
      {stage0_22[504]},
      {stage1_22[266]}
   );
   gpc1_1 gpc2018 (
      {stage0_22[505]},
      {stage1_22[267]}
   );
   gpc1_1 gpc2019 (
      {stage0_22[506]},
      {stage1_22[268]}
   );
   gpc1_1 gpc2020 (
      {stage0_22[507]},
      {stage1_22[269]}
   );
   gpc1_1 gpc2021 (
      {stage0_22[508]},
      {stage1_22[270]}
   );
   gpc1_1 gpc2022 (
      {stage0_22[509]},
      {stage1_22[271]}
   );
   gpc1_1 gpc2023 (
      {stage0_22[510]},
      {stage1_22[272]}
   );
   gpc1_1 gpc2024 (
      {stage0_22[511]},
      {stage1_22[273]}
   );
   gpc1_1 gpc2025 (
      {stage0_23[500]},
      {stage1_23[154]}
   );
   gpc1_1 gpc2026 (
      {stage0_23[501]},
      {stage1_23[155]}
   );
   gpc1_1 gpc2027 (
      {stage0_23[502]},
      {stage1_23[156]}
   );
   gpc1_1 gpc2028 (
      {stage0_23[503]},
      {stage1_23[157]}
   );
   gpc1_1 gpc2029 (
      {stage0_23[504]},
      {stage1_23[158]}
   );
   gpc1_1 gpc2030 (
      {stage0_23[505]},
      {stage1_23[159]}
   );
   gpc1_1 gpc2031 (
      {stage0_23[506]},
      {stage1_23[160]}
   );
   gpc1_1 gpc2032 (
      {stage0_23[507]},
      {stage1_23[161]}
   );
   gpc1_1 gpc2033 (
      {stage0_23[508]},
      {stage1_23[162]}
   );
   gpc1_1 gpc2034 (
      {stage0_23[509]},
      {stage1_23[163]}
   );
   gpc1_1 gpc2035 (
      {stage0_23[510]},
      {stage1_23[164]}
   );
   gpc1_1 gpc2036 (
      {stage0_23[511]},
      {stage1_23[165]}
   );
   gpc1_1 gpc2037 (
      {stage0_25[482]},
      {stage1_25[244]}
   );
   gpc1_1 gpc2038 (
      {stage0_25[483]},
      {stage1_25[245]}
   );
   gpc1_1 gpc2039 (
      {stage0_25[484]},
      {stage1_25[246]}
   );
   gpc1_1 gpc2040 (
      {stage0_25[485]},
      {stage1_25[247]}
   );
   gpc1_1 gpc2041 (
      {stage0_25[486]},
      {stage1_25[248]}
   );
   gpc1_1 gpc2042 (
      {stage0_25[487]},
      {stage1_25[249]}
   );
   gpc1_1 gpc2043 (
      {stage0_25[488]},
      {stage1_25[250]}
   );
   gpc1_1 gpc2044 (
      {stage0_25[489]},
      {stage1_25[251]}
   );
   gpc1_1 gpc2045 (
      {stage0_25[490]},
      {stage1_25[252]}
   );
   gpc1_1 gpc2046 (
      {stage0_25[491]},
      {stage1_25[253]}
   );
   gpc1_1 gpc2047 (
      {stage0_25[492]},
      {stage1_25[254]}
   );
   gpc1_1 gpc2048 (
      {stage0_25[493]},
      {stage1_25[255]}
   );
   gpc1_1 gpc2049 (
      {stage0_25[494]},
      {stage1_25[256]}
   );
   gpc1_1 gpc2050 (
      {stage0_25[495]},
      {stage1_25[257]}
   );
   gpc1_1 gpc2051 (
      {stage0_25[496]},
      {stage1_25[258]}
   );
   gpc1_1 gpc2052 (
      {stage0_25[497]},
      {stage1_25[259]}
   );
   gpc1_1 gpc2053 (
      {stage0_25[498]},
      {stage1_25[260]}
   );
   gpc1_1 gpc2054 (
      {stage0_25[499]},
      {stage1_25[261]}
   );
   gpc1_1 gpc2055 (
      {stage0_25[500]},
      {stage1_25[262]}
   );
   gpc1_1 gpc2056 (
      {stage0_25[501]},
      {stage1_25[263]}
   );
   gpc1_1 gpc2057 (
      {stage0_25[502]},
      {stage1_25[264]}
   );
   gpc1_1 gpc2058 (
      {stage0_25[503]},
      {stage1_25[265]}
   );
   gpc1_1 gpc2059 (
      {stage0_25[504]},
      {stage1_25[266]}
   );
   gpc1_1 gpc2060 (
      {stage0_25[505]},
      {stage1_25[267]}
   );
   gpc1_1 gpc2061 (
      {stage0_25[506]},
      {stage1_25[268]}
   );
   gpc1_1 gpc2062 (
      {stage0_25[507]},
      {stage1_25[269]}
   );
   gpc1_1 gpc2063 (
      {stage0_25[508]},
      {stage1_25[270]}
   );
   gpc1_1 gpc2064 (
      {stage0_25[509]},
      {stage1_25[271]}
   );
   gpc1_1 gpc2065 (
      {stage0_25[510]},
      {stage1_25[272]}
   );
   gpc1_1 gpc2066 (
      {stage0_25[511]},
      {stage1_25[273]}
   );
   gpc1_1 gpc2067 (
      {stage0_26[498]},
      {stage1_26[177]}
   );
   gpc1_1 gpc2068 (
      {stage0_26[499]},
      {stage1_26[178]}
   );
   gpc1_1 gpc2069 (
      {stage0_26[500]},
      {stage1_26[179]}
   );
   gpc1_1 gpc2070 (
      {stage0_26[501]},
      {stage1_26[180]}
   );
   gpc1_1 gpc2071 (
      {stage0_26[502]},
      {stage1_26[181]}
   );
   gpc1_1 gpc2072 (
      {stage0_26[503]},
      {stage1_26[182]}
   );
   gpc1_1 gpc2073 (
      {stage0_26[504]},
      {stage1_26[183]}
   );
   gpc1_1 gpc2074 (
      {stage0_26[505]},
      {stage1_26[184]}
   );
   gpc1_1 gpc2075 (
      {stage0_26[506]},
      {stage1_26[185]}
   );
   gpc1_1 gpc2076 (
      {stage0_26[507]},
      {stage1_26[186]}
   );
   gpc1_1 gpc2077 (
      {stage0_26[508]},
      {stage1_26[187]}
   );
   gpc1_1 gpc2078 (
      {stage0_26[509]},
      {stage1_26[188]}
   );
   gpc1_1 gpc2079 (
      {stage0_26[510]},
      {stage1_26[189]}
   );
   gpc1_1 gpc2080 (
      {stage0_26[511]},
      {stage1_26[190]}
   );
   gpc1_1 gpc2081 (
      {stage0_27[479]},
      {stage1_27[167]}
   );
   gpc1_1 gpc2082 (
      {stage0_27[480]},
      {stage1_27[168]}
   );
   gpc1_1 gpc2083 (
      {stage0_27[481]},
      {stage1_27[169]}
   );
   gpc1_1 gpc2084 (
      {stage0_27[482]},
      {stage1_27[170]}
   );
   gpc1_1 gpc2085 (
      {stage0_27[483]},
      {stage1_27[171]}
   );
   gpc1_1 gpc2086 (
      {stage0_27[484]},
      {stage1_27[172]}
   );
   gpc1_1 gpc2087 (
      {stage0_27[485]},
      {stage1_27[173]}
   );
   gpc1_1 gpc2088 (
      {stage0_27[486]},
      {stage1_27[174]}
   );
   gpc1_1 gpc2089 (
      {stage0_27[487]},
      {stage1_27[175]}
   );
   gpc1_1 gpc2090 (
      {stage0_27[488]},
      {stage1_27[176]}
   );
   gpc1_1 gpc2091 (
      {stage0_27[489]},
      {stage1_27[177]}
   );
   gpc1_1 gpc2092 (
      {stage0_27[490]},
      {stage1_27[178]}
   );
   gpc1_1 gpc2093 (
      {stage0_27[491]},
      {stage1_27[179]}
   );
   gpc1_1 gpc2094 (
      {stage0_27[492]},
      {stage1_27[180]}
   );
   gpc1_1 gpc2095 (
      {stage0_27[493]},
      {stage1_27[181]}
   );
   gpc1_1 gpc2096 (
      {stage0_27[494]},
      {stage1_27[182]}
   );
   gpc1_1 gpc2097 (
      {stage0_27[495]},
      {stage1_27[183]}
   );
   gpc1_1 gpc2098 (
      {stage0_27[496]},
      {stage1_27[184]}
   );
   gpc1_1 gpc2099 (
      {stage0_27[497]},
      {stage1_27[185]}
   );
   gpc1_1 gpc2100 (
      {stage0_27[498]},
      {stage1_27[186]}
   );
   gpc1_1 gpc2101 (
      {stage0_27[499]},
      {stage1_27[187]}
   );
   gpc1_1 gpc2102 (
      {stage0_27[500]},
      {stage1_27[188]}
   );
   gpc1_1 gpc2103 (
      {stage0_27[501]},
      {stage1_27[189]}
   );
   gpc1_1 gpc2104 (
      {stage0_27[502]},
      {stage1_27[190]}
   );
   gpc1_1 gpc2105 (
      {stage0_27[503]},
      {stage1_27[191]}
   );
   gpc1_1 gpc2106 (
      {stage0_27[504]},
      {stage1_27[192]}
   );
   gpc1_1 gpc2107 (
      {stage0_27[505]},
      {stage1_27[193]}
   );
   gpc1_1 gpc2108 (
      {stage0_27[506]},
      {stage1_27[194]}
   );
   gpc1_1 gpc2109 (
      {stage0_27[507]},
      {stage1_27[195]}
   );
   gpc1_1 gpc2110 (
      {stage0_27[508]},
      {stage1_27[196]}
   );
   gpc1_1 gpc2111 (
      {stage0_27[509]},
      {stage1_27[197]}
   );
   gpc1_1 gpc2112 (
      {stage0_27[510]},
      {stage1_27[198]}
   );
   gpc1_1 gpc2113 (
      {stage0_27[511]},
      {stage1_27[199]}
   );
   gpc1_1 gpc2114 (
      {stage0_28[506]},
      {stage1_28[242]}
   );
   gpc1_1 gpc2115 (
      {stage0_28[507]},
      {stage1_28[243]}
   );
   gpc1_1 gpc2116 (
      {stage0_28[508]},
      {stage1_28[244]}
   );
   gpc1_1 gpc2117 (
      {stage0_28[509]},
      {stage1_28[245]}
   );
   gpc1_1 gpc2118 (
      {stage0_28[510]},
      {stage1_28[246]}
   );
   gpc1_1 gpc2119 (
      {stage0_28[511]},
      {stage1_28[247]}
   );
   gpc1_1 gpc2120 (
      {stage0_29[509]},
      {stage1_29[240]}
   );
   gpc1_1 gpc2121 (
      {stage0_29[510]},
      {stage1_29[241]}
   );
   gpc1_1 gpc2122 (
      {stage0_29[511]},
      {stage1_29[242]}
   );
   gpc1_1 gpc2123 (
      {stage0_30[474]},
      {stage1_30[169]}
   );
   gpc1_1 gpc2124 (
      {stage0_30[475]},
      {stage1_30[170]}
   );
   gpc1_1 gpc2125 (
      {stage0_30[476]},
      {stage1_30[171]}
   );
   gpc1_1 gpc2126 (
      {stage0_30[477]},
      {stage1_30[172]}
   );
   gpc1_1 gpc2127 (
      {stage0_30[478]},
      {stage1_30[173]}
   );
   gpc1_1 gpc2128 (
      {stage0_30[479]},
      {stage1_30[174]}
   );
   gpc1_1 gpc2129 (
      {stage0_30[480]},
      {stage1_30[175]}
   );
   gpc1_1 gpc2130 (
      {stage0_30[481]},
      {stage1_30[176]}
   );
   gpc1_1 gpc2131 (
      {stage0_30[482]},
      {stage1_30[177]}
   );
   gpc1_1 gpc2132 (
      {stage0_30[483]},
      {stage1_30[178]}
   );
   gpc1_1 gpc2133 (
      {stage0_30[484]},
      {stage1_30[179]}
   );
   gpc1_1 gpc2134 (
      {stage0_30[485]},
      {stage1_30[180]}
   );
   gpc1_1 gpc2135 (
      {stage0_30[486]},
      {stage1_30[181]}
   );
   gpc1_1 gpc2136 (
      {stage0_30[487]},
      {stage1_30[182]}
   );
   gpc1_1 gpc2137 (
      {stage0_30[488]},
      {stage1_30[183]}
   );
   gpc1_1 gpc2138 (
      {stage0_30[489]},
      {stage1_30[184]}
   );
   gpc1_1 gpc2139 (
      {stage0_30[490]},
      {stage1_30[185]}
   );
   gpc1_1 gpc2140 (
      {stage0_30[491]},
      {stage1_30[186]}
   );
   gpc1_1 gpc2141 (
      {stage0_30[492]},
      {stage1_30[187]}
   );
   gpc1_1 gpc2142 (
      {stage0_30[493]},
      {stage1_30[188]}
   );
   gpc1_1 gpc2143 (
      {stage0_30[494]},
      {stage1_30[189]}
   );
   gpc1_1 gpc2144 (
      {stage0_30[495]},
      {stage1_30[190]}
   );
   gpc1_1 gpc2145 (
      {stage0_30[496]},
      {stage1_30[191]}
   );
   gpc1_1 gpc2146 (
      {stage0_30[497]},
      {stage1_30[192]}
   );
   gpc1_1 gpc2147 (
      {stage0_30[498]},
      {stage1_30[193]}
   );
   gpc1_1 gpc2148 (
      {stage0_30[499]},
      {stage1_30[194]}
   );
   gpc1_1 gpc2149 (
      {stage0_30[500]},
      {stage1_30[195]}
   );
   gpc1_1 gpc2150 (
      {stage0_30[501]},
      {stage1_30[196]}
   );
   gpc1_1 gpc2151 (
      {stage0_30[502]},
      {stage1_30[197]}
   );
   gpc1_1 gpc2152 (
      {stage0_30[503]},
      {stage1_30[198]}
   );
   gpc1_1 gpc2153 (
      {stage0_30[504]},
      {stage1_30[199]}
   );
   gpc1_1 gpc2154 (
      {stage0_30[505]},
      {stage1_30[200]}
   );
   gpc1_1 gpc2155 (
      {stage0_30[506]},
      {stage1_30[201]}
   );
   gpc1_1 gpc2156 (
      {stage0_30[507]},
      {stage1_30[202]}
   );
   gpc1_1 gpc2157 (
      {stage0_30[508]},
      {stage1_30[203]}
   );
   gpc1_1 gpc2158 (
      {stage0_30[509]},
      {stage1_30[204]}
   );
   gpc1_1 gpc2159 (
      {stage0_30[510]},
      {stage1_30[205]}
   );
   gpc1_1 gpc2160 (
      {stage0_30[511]},
      {stage1_30[206]}
   );
   gpc1_1 gpc2161 (
      {stage0_31[426]},
      {stage1_31[157]}
   );
   gpc1_1 gpc2162 (
      {stage0_31[427]},
      {stage1_31[158]}
   );
   gpc1_1 gpc2163 (
      {stage0_31[428]},
      {stage1_31[159]}
   );
   gpc1_1 gpc2164 (
      {stage0_31[429]},
      {stage1_31[160]}
   );
   gpc1_1 gpc2165 (
      {stage0_31[430]},
      {stage1_31[161]}
   );
   gpc1_1 gpc2166 (
      {stage0_31[431]},
      {stage1_31[162]}
   );
   gpc1_1 gpc2167 (
      {stage0_31[432]},
      {stage1_31[163]}
   );
   gpc1_1 gpc2168 (
      {stage0_31[433]},
      {stage1_31[164]}
   );
   gpc1_1 gpc2169 (
      {stage0_31[434]},
      {stage1_31[165]}
   );
   gpc1_1 gpc2170 (
      {stage0_31[435]},
      {stage1_31[166]}
   );
   gpc1_1 gpc2171 (
      {stage0_31[436]},
      {stage1_31[167]}
   );
   gpc1_1 gpc2172 (
      {stage0_31[437]},
      {stage1_31[168]}
   );
   gpc1_1 gpc2173 (
      {stage0_31[438]},
      {stage1_31[169]}
   );
   gpc1_1 gpc2174 (
      {stage0_31[439]},
      {stage1_31[170]}
   );
   gpc1_1 gpc2175 (
      {stage0_31[440]},
      {stage1_31[171]}
   );
   gpc1_1 gpc2176 (
      {stage0_31[441]},
      {stage1_31[172]}
   );
   gpc1_1 gpc2177 (
      {stage0_31[442]},
      {stage1_31[173]}
   );
   gpc1_1 gpc2178 (
      {stage0_31[443]},
      {stage1_31[174]}
   );
   gpc1_1 gpc2179 (
      {stage0_31[444]},
      {stage1_31[175]}
   );
   gpc1_1 gpc2180 (
      {stage0_31[445]},
      {stage1_31[176]}
   );
   gpc1_1 gpc2181 (
      {stage0_31[446]},
      {stage1_31[177]}
   );
   gpc1_1 gpc2182 (
      {stage0_31[447]},
      {stage1_31[178]}
   );
   gpc1_1 gpc2183 (
      {stage0_31[448]},
      {stage1_31[179]}
   );
   gpc1_1 gpc2184 (
      {stage0_31[449]},
      {stage1_31[180]}
   );
   gpc1_1 gpc2185 (
      {stage0_31[450]},
      {stage1_31[181]}
   );
   gpc1_1 gpc2186 (
      {stage0_31[451]},
      {stage1_31[182]}
   );
   gpc1_1 gpc2187 (
      {stage0_31[452]},
      {stage1_31[183]}
   );
   gpc1_1 gpc2188 (
      {stage0_31[453]},
      {stage1_31[184]}
   );
   gpc1_1 gpc2189 (
      {stage0_31[454]},
      {stage1_31[185]}
   );
   gpc1_1 gpc2190 (
      {stage0_31[455]},
      {stage1_31[186]}
   );
   gpc1_1 gpc2191 (
      {stage0_31[456]},
      {stage1_31[187]}
   );
   gpc1_1 gpc2192 (
      {stage0_31[457]},
      {stage1_31[188]}
   );
   gpc1_1 gpc2193 (
      {stage0_31[458]},
      {stage1_31[189]}
   );
   gpc1_1 gpc2194 (
      {stage0_31[459]},
      {stage1_31[190]}
   );
   gpc1_1 gpc2195 (
      {stage0_31[460]},
      {stage1_31[191]}
   );
   gpc1_1 gpc2196 (
      {stage0_31[461]},
      {stage1_31[192]}
   );
   gpc1_1 gpc2197 (
      {stage0_31[462]},
      {stage1_31[193]}
   );
   gpc1_1 gpc2198 (
      {stage0_31[463]},
      {stage1_31[194]}
   );
   gpc1_1 gpc2199 (
      {stage0_31[464]},
      {stage1_31[195]}
   );
   gpc1_1 gpc2200 (
      {stage0_31[465]},
      {stage1_31[196]}
   );
   gpc1_1 gpc2201 (
      {stage0_31[466]},
      {stage1_31[197]}
   );
   gpc1_1 gpc2202 (
      {stage0_31[467]},
      {stage1_31[198]}
   );
   gpc1_1 gpc2203 (
      {stage0_31[468]},
      {stage1_31[199]}
   );
   gpc1_1 gpc2204 (
      {stage0_31[469]},
      {stage1_31[200]}
   );
   gpc1_1 gpc2205 (
      {stage0_31[470]},
      {stage1_31[201]}
   );
   gpc1_1 gpc2206 (
      {stage0_31[471]},
      {stage1_31[202]}
   );
   gpc1_1 gpc2207 (
      {stage0_31[472]},
      {stage1_31[203]}
   );
   gpc1_1 gpc2208 (
      {stage0_31[473]},
      {stage1_31[204]}
   );
   gpc1_1 gpc2209 (
      {stage0_31[474]},
      {stage1_31[205]}
   );
   gpc1_1 gpc2210 (
      {stage0_31[475]},
      {stage1_31[206]}
   );
   gpc1_1 gpc2211 (
      {stage0_31[476]},
      {stage1_31[207]}
   );
   gpc1_1 gpc2212 (
      {stage0_31[477]},
      {stage1_31[208]}
   );
   gpc1_1 gpc2213 (
      {stage0_31[478]},
      {stage1_31[209]}
   );
   gpc1_1 gpc2214 (
      {stage0_31[479]},
      {stage1_31[210]}
   );
   gpc1_1 gpc2215 (
      {stage0_31[480]},
      {stage1_31[211]}
   );
   gpc1_1 gpc2216 (
      {stage0_31[481]},
      {stage1_31[212]}
   );
   gpc1_1 gpc2217 (
      {stage0_31[482]},
      {stage1_31[213]}
   );
   gpc1_1 gpc2218 (
      {stage0_31[483]},
      {stage1_31[214]}
   );
   gpc1_1 gpc2219 (
      {stage0_31[484]},
      {stage1_31[215]}
   );
   gpc1_1 gpc2220 (
      {stage0_31[485]},
      {stage1_31[216]}
   );
   gpc1_1 gpc2221 (
      {stage0_31[486]},
      {stage1_31[217]}
   );
   gpc1_1 gpc2222 (
      {stage0_31[487]},
      {stage1_31[218]}
   );
   gpc1_1 gpc2223 (
      {stage0_31[488]},
      {stage1_31[219]}
   );
   gpc1_1 gpc2224 (
      {stage0_31[489]},
      {stage1_31[220]}
   );
   gpc1_1 gpc2225 (
      {stage0_31[490]},
      {stage1_31[221]}
   );
   gpc1_1 gpc2226 (
      {stage0_31[491]},
      {stage1_31[222]}
   );
   gpc1_1 gpc2227 (
      {stage0_31[492]},
      {stage1_31[223]}
   );
   gpc1_1 gpc2228 (
      {stage0_31[493]},
      {stage1_31[224]}
   );
   gpc1_1 gpc2229 (
      {stage0_31[494]},
      {stage1_31[225]}
   );
   gpc1_1 gpc2230 (
      {stage0_31[495]},
      {stage1_31[226]}
   );
   gpc1_1 gpc2231 (
      {stage0_31[496]},
      {stage1_31[227]}
   );
   gpc1_1 gpc2232 (
      {stage0_31[497]},
      {stage1_31[228]}
   );
   gpc1_1 gpc2233 (
      {stage0_31[498]},
      {stage1_31[229]}
   );
   gpc1_1 gpc2234 (
      {stage0_31[499]},
      {stage1_31[230]}
   );
   gpc1_1 gpc2235 (
      {stage0_31[500]},
      {stage1_31[231]}
   );
   gpc1_1 gpc2236 (
      {stage0_31[501]},
      {stage1_31[232]}
   );
   gpc1_1 gpc2237 (
      {stage0_31[502]},
      {stage1_31[233]}
   );
   gpc1_1 gpc2238 (
      {stage0_31[503]},
      {stage1_31[234]}
   );
   gpc1_1 gpc2239 (
      {stage0_31[504]},
      {stage1_31[235]}
   );
   gpc1_1 gpc2240 (
      {stage0_31[505]},
      {stage1_31[236]}
   );
   gpc1_1 gpc2241 (
      {stage0_31[506]},
      {stage1_31[237]}
   );
   gpc1_1 gpc2242 (
      {stage0_31[507]},
      {stage1_31[238]}
   );
   gpc1_1 gpc2243 (
      {stage0_31[508]},
      {stage1_31[239]}
   );
   gpc1_1 gpc2244 (
      {stage0_31[509]},
      {stage1_31[240]}
   );
   gpc1_1 gpc2245 (
      {stage0_31[510]},
      {stage1_31[241]}
   );
   gpc1_1 gpc2246 (
      {stage0_31[511]},
      {stage1_31[242]}
   );
   gpc2135_5 gpc2247 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc2248 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc2249 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc2250 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc2251 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24]},
      {stage1_1[12]},
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc2252 (
      {stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc2253 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34]},
      {stage1_1[14]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc615_5 gpc2254 (
      {stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39]},
      {stage1_1[15]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc615_5 gpc2255 (
      {stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_1[16]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc615_5 gpc2256 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_1[17]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc615_5 gpc2257 (
      {stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54]},
      {stage1_1[18]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc615_5 gpc2258 (
      {stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_1[19]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2259 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage2_5[0],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc2260 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage2_5[1],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc2261 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25]},
      {stage2_5[2],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc2262 (
      {stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42], stage1_1[43]},
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage2_5[3],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc2263 (
      {stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48], stage1_1[49]},
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage2_5[4],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc2264 (
      {stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54], stage1_1[55]},
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage2_5[5],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc2265 (
      {stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59], stage1_1[60], stage1_1[61]},
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage2_5[6],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc2266 (
      {stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65], stage1_1[66], stage1_1[67]},
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage2_5[7],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc606_5 gpc2267 (
      {stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71], stage1_1[72], stage1_1[73]},
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage2_5[8],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc606_5 gpc2268 (
      {stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78], stage1_1[79]},
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67]},
      {stage2_5[9],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc2269 (
      {stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83], stage1_1[84], stage1_1[85]},
      {stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73]},
      {stage2_5[10],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc2270 (
      {stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89], stage1_1[90], stage1_1[91]},
      {stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79]},
      {stage2_5[11],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc2271 (
      {stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95], stage1_1[96], stage1_1[97]},
      {stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage2_5[12],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc2272 (
      {stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102], stage1_1[103]},
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage2_5[13],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc2273 (
      {stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108], stage1_1[109]},
      {stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97]},
      {stage2_5[14],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc2274 (
      {stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114], stage1_1[115]},
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102], stage1_3[103]},
      {stage2_5[15],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc2275 (
      {stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120], stage1_1[121]},
      {stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109]},
      {stage2_5[16],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc2276 (
      {stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126], stage1_1[127]},
      {stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage2_5[17],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc2277 (
      {stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132], stage1_1[133]},
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120], stage1_3[121]},
      {stage2_5[18],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc2278 (
      {stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138], stage1_1[139]},
      {stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127]},
      {stage2_5[19],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc2279 (
      {stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144], stage1_1[145]},
      {stage1_3[128], stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132], stage1_3[133]},
      {stage2_5[20],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc2280 (
      {stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150], stage1_1[151]},
      {stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139]},
      {stage2_5[21],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc2281 (
      {stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156], stage1_1[157]},
      {stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage2_5[22],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc2282 (
      {stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162], stage1_1[163]},
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150], stage1_3[151]},
      {stage2_5[23],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc2283 (
      {stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168], stage1_1[169]},
      {stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157]},
      {stage2_5[24],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc2284 (
      {stage1_1[170], stage1_1[171], stage1_1[172], stage1_1[173], stage1_1[174], stage1_1[175]},
      {stage1_3[158], stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage2_5[25],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc2285 (
      {stage1_1[176], stage1_1[177], stage1_1[178], stage1_1[179], stage1_1[180], stage1_1[181]},
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169]},
      {stage2_5[26],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc615_5 gpc2286 (
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56]},
      {stage1_3[170]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[27],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc2287 (
      {stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61]},
      {stage1_3[171]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[28],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc2288 (
      {stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66]},
      {stage1_3[172]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[29],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc2289 (
      {stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_3[173]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[30],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc2290 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76]},
      {stage1_3[174]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[31],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc2291 (
      {stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage1_3[175]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[32],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc2292 (
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86]},
      {stage1_3[176]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[33],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc2293 (
      {stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91]},
      {stage1_3[177]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[34],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc2294 (
      {stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96]},
      {stage1_3[178]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[35],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc2295 (
      {stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101]},
      {stage1_3[179]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[36],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc2296 (
      {stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106]},
      {stage1_3[180]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[37],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc2297 (
      {stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage1_3[181]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[38],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc2298 (
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116]},
      {stage1_3[182]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[39],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc2299 (
      {stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121]},
      {stage1_3[183]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[40],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc2300 (
      {stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126]},
      {stage1_3[184]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[41],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc2301 (
      {stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131]},
      {stage1_3[185]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[42],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc615_5 gpc2302 (
      {stage1_2[132], stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136]},
      {stage1_3[186]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[43],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc615_5 gpc2303 (
      {stage1_2[137], stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141]},
      {stage1_3[187]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[44],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc615_5 gpc2304 (
      {stage1_2[142], stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146]},
      {stage1_3[188]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[45],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc615_5 gpc2305 (
      {stage1_2[147], stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151]},
      {stage1_3[189]},
      {stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119]},
      {stage2_6[19],stage2_5[46],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc615_5 gpc2306 (
      {stage1_3[190], stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194]},
      {stage1_4[120]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[20],stage2_5[47],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc2307 (
      {stage1_3[195], stage1_3[196], stage1_3[197], stage1_3[198], stage1_3[199]},
      {stage1_4[121]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[21],stage2_5[48],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc2308 (
      {stage1_3[200], stage1_3[201], stage1_3[202], stage1_3[203], stage1_3[204]},
      {stage1_4[122]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[22],stage2_5[49],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc2309 (
      {stage1_3[205], stage1_3[206], stage1_3[207], stage1_3[208], stage1_3[209]},
      {stage1_4[123]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[23],stage2_5[50],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc2310 (
      {stage1_3[210], stage1_3[211], stage1_3[212], stage1_3[213], stage1_3[214]},
      {stage1_4[124]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[24],stage2_5[51],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc2311 (
      {stage1_3[215], stage1_3[216], stage1_3[217], stage1_3[218], stage1_3[219]},
      {stage1_4[125]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[25],stage2_5[52],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc2312 (
      {stage1_3[220], stage1_3[221], stage1_3[222], stage1_3[223], stage1_3[224]},
      {stage1_4[126]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[26],stage2_5[53],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc2313 (
      {stage1_3[225], stage1_3[226], stage1_3[227], stage1_3[228], stage1_3[229]},
      {stage1_4[127]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[27],stage2_5[54],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc2314 (
      {stage1_3[230], stage1_3[231], stage1_3[232], stage1_3[233], stage1_3[234]},
      {stage1_4[128]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[28],stage2_5[55],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc2315 (
      {stage1_3[235], stage1_3[236], stage1_3[237], stage1_3[238], stage1_3[239]},
      {stage1_4[129]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[29],stage2_5[56],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc2316 (
      {stage1_3[240], stage1_3[241], stage1_3[242], stage1_3[243], stage1_3[244]},
      {stage1_4[130]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[30],stage2_5[57],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc2317 (
      {stage1_3[245], stage1_3[246], stage1_3[247], stage1_3[248], stage1_3[249]},
      {stage1_4[131]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[31],stage2_5[58],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc2318 (
      {stage1_3[250], stage1_3[251], stage1_3[252], stage1_3[253], stage1_3[254]},
      {stage1_4[132]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[32],stage2_5[59],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc2319 (
      {stage1_3[255], stage1_3[256], stage1_3[257], stage1_3[258], stage1_3[259]},
      {stage1_4[133]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[33],stage2_5[60],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc2320 (
      {stage1_3[260], stage1_3[261], stage1_3[262], stage1_3[263], stage1_3[264]},
      {stage1_4[134]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[34],stage2_5[61],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc2321 (
      {stage1_3[265], stage1_3[266], stage1_3[267], stage1_3[268], stage1_3[269]},
      {stage1_4[135]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[35],stage2_5[62],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc2322 (
      {stage1_3[270], stage1_3[271], stage1_3[272], stage1_3[273], stage1_3[274]},
      {stage1_4[136]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[36],stage2_5[63],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc2323 (
      {stage1_3[275], stage1_3[276], 1'b0, 1'b0, 1'b0},
      {stage1_4[137]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[37],stage2_5[64],stage2_4[76],stage2_3[76]}
   );
   gpc1163_5 gpc2324 (
      {stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[18],stage2_6[38],stage2_5[65],stage2_4[77]}
   );
   gpc606_5 gpc2325 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[19],stage2_6[39],stage2_5[66],stage2_4[78]}
   );
   gpc606_5 gpc2326 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[20],stage2_6[40],stage2_5[67],stage2_4[79]}
   );
   gpc606_5 gpc2327 (
      {stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[21],stage2_6[41],stage2_5[68],stage2_4[80]}
   );
   gpc606_5 gpc2328 (
      {stage1_4[159], stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[22],stage2_6[42],stage2_5[69],stage2_4[81]}
   );
   gpc606_5 gpc2329 (
      {stage1_4[165], stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[23],stage2_6[43],stage2_5[70],stage2_4[82]}
   );
   gpc606_5 gpc2330 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[24],stage2_6[44],stage2_5[71],stage2_4[83]}
   );
   gpc606_5 gpc2331 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[25],stage2_6[45],stage2_5[72],stage2_4[84]}
   );
   gpc606_5 gpc2332 (
      {stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[26],stage2_6[46],stage2_5[73],stage2_4[85]}
   );
   gpc606_5 gpc2333 (
      {stage1_4[189], stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[27],stage2_6[47],stage2_5[74],stage2_4[86]}
   );
   gpc606_5 gpc2334 (
      {stage1_4[195], stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[28],stage2_6[48],stage2_5[75],stage2_4[87]}
   );
   gpc606_5 gpc2335 (
      {stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[29],stage2_6[49],stage2_5[76],stage2_4[88]}
   );
   gpc615_5 gpc2336 (
      {stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211]},
      {stage1_5[114]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[30],stage2_6[50],stage2_5[77],stage2_4[89]}
   );
   gpc615_5 gpc2337 (
      {stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_5[115]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[31],stage2_6[51],stage2_5[78],stage2_4[90]}
   );
   gpc606_5 gpc2338 (
      {stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119], stage1_5[120], stage1_5[121]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[14],stage2_7[32],stage2_6[52],stage2_5[79]}
   );
   gpc606_5 gpc2339 (
      {stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125], stage1_5[126], stage1_5[127]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[15],stage2_7[33],stage2_6[53],stage2_5[80]}
   );
   gpc606_5 gpc2340 (
      {stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131], stage1_5[132], stage1_5[133]},
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage2_9[2],stage2_8[16],stage2_7[34],stage2_6[54],stage2_5[81]}
   );
   gpc606_5 gpc2341 (
      {stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137], stage1_5[138], stage1_5[139]},
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage2_9[3],stage2_8[17],stage2_7[35],stage2_6[55],stage2_5[82]}
   );
   gpc606_5 gpc2342 (
      {stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143], stage1_5[144], stage1_5[145]},
      {stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30]},
      {stage2_9[4],stage2_8[18],stage2_7[36],stage2_6[56],stage2_5[83]}
   );
   gpc606_5 gpc2343 (
      {stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149], stage1_5[150], stage1_5[151]},
      {stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage2_9[5],stage2_8[19],stage2_7[37],stage2_6[57],stage2_5[84]}
   );
   gpc606_5 gpc2344 (
      {stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157]},
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage2_9[6],stage2_8[20],stage2_7[38],stage2_6[58],stage2_5[85]}
   );
   gpc606_5 gpc2345 (
      {stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163]},
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage2_9[7],stage2_8[21],stage2_7[39],stage2_6[59],stage2_5[86]}
   );
   gpc606_5 gpc2346 (
      {stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169]},
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage2_9[8],stage2_8[22],stage2_7[40],stage2_6[60],stage2_5[87]}
   );
   gpc606_5 gpc2347 (
      {stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175]},
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60]},
      {stage2_9[9],stage2_8[23],stage2_7[41],stage2_6[61],stage2_5[88]}
   );
   gpc606_5 gpc2348 (
      {stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181]},
      {stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage2_9[10],stage2_8[24],stage2_7[42],stage2_6[62],stage2_5[89]}
   );
   gpc606_5 gpc2349 (
      {stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187]},
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71], stage1_7[72]},
      {stage2_9[11],stage2_8[25],stage2_7[43],stage2_6[63],stage2_5[90]}
   );
   gpc606_5 gpc2350 (
      {stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191], stage1_5[192], stage1_5[193]},
      {stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77], stage1_7[78]},
      {stage2_9[12],stage2_8[26],stage2_7[44],stage2_6[64],stage2_5[91]}
   );
   gpc606_5 gpc2351 (
      {stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197], stage1_5[198], stage1_5[199]},
      {stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83], stage1_7[84]},
      {stage2_9[13],stage2_8[27],stage2_7[45],stage2_6[65],stage2_5[92]}
   );
   gpc606_5 gpc2352 (
      {stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203], stage1_5[204], stage1_5[205]},
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90]},
      {stage2_9[14],stage2_8[28],stage2_7[46],stage2_6[66],stage2_5[93]}
   );
   gpc606_5 gpc2353 (
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[15],stage2_8[29],stage2_7[47],stage2_6[67]}
   );
   gpc606_5 gpc2354 (
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[16],stage2_8[30],stage2_7[48],stage2_6[68]}
   );
   gpc606_5 gpc2355 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[17],stage2_8[31],stage2_7[49],stage2_6[69]}
   );
   gpc606_5 gpc2356 (
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[18],stage2_8[32],stage2_7[50],stage2_6[70]}
   );
   gpc606_5 gpc2357 (
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[19],stage2_8[33],stage2_7[51],stage2_6[71]}
   );
   gpc606_5 gpc2358 (
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[20],stage2_8[34],stage2_7[52],stage2_6[72]}
   );
   gpc606_5 gpc2359 (
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[21],stage2_8[35],stage2_7[53],stage2_6[73]}
   );
   gpc606_5 gpc2360 (
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[22],stage2_8[36],stage2_7[54],stage2_6[74]}
   );
   gpc606_5 gpc2361 (
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131], stage1_6[132]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[23],stage2_8[37],stage2_7[55],stage2_6[75]}
   );
   gpc606_5 gpc2362 (
      {stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137], stage1_6[138]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[24],stage2_8[38],stage2_7[56],stage2_6[76]}
   );
   gpc606_5 gpc2363 (
      {stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143], stage1_6[144]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[25],stage2_8[39],stage2_7[57],stage2_6[77]}
   );
   gpc606_5 gpc2364 (
      {stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[26],stage2_8[40],stage2_7[58],stage2_6[78]}
   );
   gpc606_5 gpc2365 (
      {stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[27],stage2_8[41],stage2_7[59],stage2_6[79]}
   );
   gpc606_5 gpc2366 (
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161], stage1_6[162]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[28],stage2_8[42],stage2_7[60],stage2_6[80]}
   );
   gpc606_5 gpc2367 (
      {stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167], stage1_6[168]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[29],stage2_8[43],stage2_7[61],stage2_6[81]}
   );
   gpc606_5 gpc2368 (
      {stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173], stage1_6[174]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[30],stage2_8[44],stage2_7[62],stage2_6[82]}
   );
   gpc606_5 gpc2369 (
      {stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178], stage1_6[179], stage1_6[180]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[31],stage2_8[45],stage2_7[63],stage2_6[83]}
   );
   gpc606_5 gpc2370 (
      {stage1_6[181], stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185], stage1_6[186]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[32],stage2_8[46],stage2_7[64],stage2_6[84]}
   );
   gpc606_5 gpc2371 (
      {stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191], stage1_6[192]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[33],stage2_8[47],stage2_7[65],stage2_6[85]}
   );
   gpc615_5 gpc2372 (
      {stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196], stage1_6[197]},
      {stage1_7[91]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[34],stage2_8[48],stage2_7[66],stage2_6[86]}
   );
   gpc615_5 gpc2373 (
      {stage1_6[198], stage1_6[199], stage1_6[200], stage1_6[201], stage1_6[202]},
      {stage1_7[92]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[35],stage2_8[49],stage2_7[67],stage2_6[87]}
   );
   gpc615_5 gpc2374 (
      {stage1_6[203], stage1_6[204], stage1_6[205], stage1_6[206], stage1_6[207]},
      {stage1_7[93]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[36],stage2_8[50],stage2_7[68],stage2_6[88]}
   );
   gpc615_5 gpc2375 (
      {stage1_6[208], stage1_6[209], stage1_6[210], stage1_6[211], stage1_6[212]},
      {stage1_7[94]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[37],stage2_8[51],stage2_7[69],stage2_6[89]}
   );
   gpc615_5 gpc2376 (
      {stage1_6[213], stage1_6[214], stage1_6[215], stage1_6[216], stage1_6[217]},
      {stage1_7[95]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[38],stage2_8[52],stage2_7[70],stage2_6[90]}
   );
   gpc615_5 gpc2377 (
      {stage1_6[218], stage1_6[219], stage1_6[220], stage1_6[221], stage1_6[222]},
      {stage1_7[96]},
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage2_10[24],stage2_9[39],stage2_8[53],stage2_7[71],stage2_6[91]}
   );
   gpc615_5 gpc2378 (
      {stage1_6[223], stage1_6[224], stage1_6[225], stage1_6[226], stage1_6[227]},
      {stage1_7[97]},
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage2_10[25],stage2_9[40],stage2_8[54],stage2_7[72],stage2_6[92]}
   );
   gpc615_5 gpc2379 (
      {stage1_6[228], stage1_6[229], stage1_6[230], stage1_6[231], stage1_6[232]},
      {stage1_7[98]},
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage2_10[26],stage2_9[41],stage2_8[55],stage2_7[73],stage2_6[93]}
   );
   gpc615_5 gpc2380 (
      {stage1_6[233], stage1_6[234], stage1_6[235], stage1_6[236], stage1_6[237]},
      {stage1_7[99]},
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage2_10[27],stage2_9[42],stage2_8[56],stage2_7[74],stage2_6[94]}
   );
   gpc615_5 gpc2381 (
      {stage1_6[238], stage1_6[239], stage1_6[240], stage1_6[241], stage1_6[242]},
      {stage1_7[100]},
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172], stage1_8[173]},
      {stage2_10[28],stage2_9[43],stage2_8[57],stage2_7[75],stage2_6[95]}
   );
   gpc615_5 gpc2382 (
      {stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105]},
      {stage1_8[174]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[29],stage2_9[44],stage2_8[58],stage2_7[76]}
   );
   gpc615_5 gpc2383 (
      {stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109], stage1_7[110]},
      {stage1_8[175]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[30],stage2_9[45],stage2_8[59],stage2_7[77]}
   );
   gpc615_5 gpc2384 (
      {stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114], stage1_7[115]},
      {stage1_8[176]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[31],stage2_9[46],stage2_8[60],stage2_7[78]}
   );
   gpc615_5 gpc2385 (
      {stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120]},
      {stage1_8[177]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[32],stage2_9[47],stage2_8[61],stage2_7[79]}
   );
   gpc615_5 gpc2386 (
      {stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125]},
      {stage1_8[178]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[33],stage2_9[48],stage2_8[62],stage2_7[80]}
   );
   gpc615_5 gpc2387 (
      {stage1_7[126], stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130]},
      {stage1_8[179]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[34],stage2_9[49],stage2_8[63],stage2_7[81]}
   );
   gpc615_5 gpc2388 (
      {stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135]},
      {stage1_8[180]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[35],stage2_9[50],stage2_8[64],stage2_7[82]}
   );
   gpc615_5 gpc2389 (
      {stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140]},
      {stage1_8[181]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[36],stage2_9[51],stage2_8[65],stage2_7[83]}
   );
   gpc615_5 gpc2390 (
      {stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145]},
      {stage1_8[182]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[37],stage2_9[52],stage2_8[66],stage2_7[84]}
   );
   gpc615_5 gpc2391 (
      {stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_8[183]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[38],stage2_9[53],stage2_8[67],stage2_7[85]}
   );
   gpc615_5 gpc2392 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155]},
      {stage1_8[184]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[39],stage2_9[54],stage2_8[68],stage2_7[86]}
   );
   gpc615_5 gpc2393 (
      {stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160]},
      {stage1_8[185]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[40],stage2_9[55],stage2_8[69],stage2_7[87]}
   );
   gpc615_5 gpc2394 (
      {stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165]},
      {stage1_8[186]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[41],stage2_9[56],stage2_8[70],stage2_7[88]}
   );
   gpc606_5 gpc2395 (
      {stage1_8[187], stage1_8[188], stage1_8[189], stage1_8[190], stage1_8[191], stage1_8[192]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[13],stage2_10[42],stage2_9[57],stage2_8[71]}
   );
   gpc606_5 gpc2396 (
      {stage1_8[193], stage1_8[194], stage1_8[195], stage1_8[196], stage1_8[197], stage1_8[198]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[14],stage2_10[43],stage2_9[58],stage2_8[72]}
   );
   gpc606_5 gpc2397 (
      {stage1_8[199], stage1_8[200], stage1_8[201], stage1_8[202], stage1_8[203], stage1_8[204]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[15],stage2_10[44],stage2_9[59],stage2_8[73]}
   );
   gpc606_5 gpc2398 (
      {stage1_8[205], stage1_8[206], stage1_8[207], stage1_8[208], stage1_8[209], stage1_8[210]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[16],stage2_10[45],stage2_9[60],stage2_8[74]}
   );
   gpc606_5 gpc2399 (
      {stage1_8[211], stage1_8[212], stage1_8[213], stage1_8[214], stage1_8[215], stage1_8[216]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[17],stage2_10[46],stage2_9[61],stage2_8[75]}
   );
   gpc606_5 gpc2400 (
      {stage1_8[217], stage1_8[218], stage1_8[219], stage1_8[220], stage1_8[221], stage1_8[222]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[18],stage2_10[47],stage2_9[62],stage2_8[76]}
   );
   gpc606_5 gpc2401 (
      {stage1_8[223], stage1_8[224], stage1_8[225], stage1_8[226], stage1_8[227], stage1_8[228]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[19],stage2_10[48],stage2_9[63],stage2_8[77]}
   );
   gpc606_5 gpc2402 (
      {stage1_8[229], stage1_8[230], stage1_8[231], stage1_8[232], stage1_8[233], stage1_8[234]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[20],stage2_10[49],stage2_9[64],stage2_8[78]}
   );
   gpc606_5 gpc2403 (
      {stage1_8[235], stage1_8[236], stage1_8[237], stage1_8[238], stage1_8[239], stage1_8[240]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[21],stage2_10[50],stage2_9[65],stage2_8[79]}
   );
   gpc606_5 gpc2404 (
      {stage1_8[241], stage1_8[242], stage1_8[243], stage1_8[244], stage1_8[245], stage1_8[246]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[22],stage2_10[51],stage2_9[66],stage2_8[80]}
   );
   gpc606_5 gpc2405 (
      {stage1_8[247], stage1_8[248], stage1_8[249], stage1_8[250], stage1_8[251], stage1_8[252]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[23],stage2_10[52],stage2_9[67],stage2_8[81]}
   );
   gpc606_5 gpc2406 (
      {stage1_8[253], stage1_8[254], stage1_8[255], stage1_8[256], stage1_8[257], stage1_8[258]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[24],stage2_10[53],stage2_9[68],stage2_8[82]}
   );
   gpc606_5 gpc2407 (
      {stage1_8[259], stage1_8[260], stage1_8[261], stage1_8[262], stage1_8[263], stage1_8[264]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[25],stage2_10[54],stage2_9[69],stage2_8[83]}
   );
   gpc606_5 gpc2408 (
      {stage1_8[265], stage1_8[266], stage1_8[267], stage1_8[268], stage1_8[269], stage1_8[270]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[26],stage2_10[55],stage2_9[70],stage2_8[84]}
   );
   gpc606_5 gpc2409 (
      {stage1_8[271], stage1_8[272], stage1_8[273], stage1_8[274], stage1_8[275], stage1_8[276]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[27],stage2_10[56],stage2_9[71],stage2_8[85]}
   );
   gpc606_5 gpc2410 (
      {stage1_8[277], stage1_8[278], stage1_8[279], stage1_8[280], stage1_8[281], stage1_8[282]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[28],stage2_10[57],stage2_9[72],stage2_8[86]}
   );
   gpc606_5 gpc2411 (
      {stage1_8[283], stage1_8[284], stage1_8[285], stage1_8[286], stage1_8[287], stage1_8[288]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[29],stage2_10[58],stage2_9[73],stage2_8[87]}
   );
   gpc606_5 gpc2412 (
      {stage1_8[289], stage1_8[290], stage1_8[291], stage1_8[292], stage1_8[293], stage1_8[294]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[30],stage2_10[59],stage2_9[74],stage2_8[88]}
   );
   gpc606_5 gpc2413 (
      {stage1_8[295], stage1_8[296], stage1_8[297], stage1_8[298], stage1_8[299], stage1_8[300]},
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage2_12[18],stage2_11[31],stage2_10[60],stage2_9[75],stage2_8[89]}
   );
   gpc606_5 gpc2414 (
      {stage1_8[301], stage1_8[302], stage1_8[303], stage1_8[304], stage1_8[305], stage1_8[306]},
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage2_12[19],stage2_11[32],stage2_10[61],stage2_9[76],stage2_8[90]}
   );
   gpc606_5 gpc2415 (
      {stage1_8[307], stage1_8[308], stage1_8[309], stage1_8[310], stage1_8[311], stage1_8[312]},
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage2_12[20],stage2_11[33],stage2_10[62],stage2_9[77],stage2_8[91]}
   );
   gpc606_5 gpc2416 (
      {stage1_8[313], stage1_8[314], stage1_8[315], stage1_8[316], stage1_8[317], stage1_8[318]},
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage2_12[21],stage2_11[34],stage2_10[63],stage2_9[78],stage2_8[92]}
   );
   gpc606_5 gpc2417 (
      {stage1_8[319], stage1_8[320], stage1_8[321], stage1_8[322], stage1_8[323], stage1_8[324]},
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage2_12[22],stage2_11[35],stage2_10[64],stage2_9[79],stage2_8[93]}
   );
   gpc606_5 gpc2418 (
      {stage1_8[325], stage1_8[326], stage1_8[327], stage1_8[328], stage1_8[329], stage1_8[330]},
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage2_12[23],stage2_11[36],stage2_10[65],stage2_9[80],stage2_8[94]}
   );
   gpc606_5 gpc2419 (
      {stage1_8[331], stage1_8[332], stage1_8[333], stage1_8[334], stage1_8[335], stage1_8[336]},
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage2_12[24],stage2_11[37],stage2_10[66],stage2_9[81],stage2_8[95]}
   );
   gpc606_5 gpc2420 (
      {stage1_8[337], stage1_8[338], stage1_8[339], stage1_8[340], stage1_8[341], stage1_8[342]},
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage2_12[25],stage2_11[38],stage2_10[67],stage2_9[82],stage2_8[96]}
   );
   gpc606_5 gpc2421 (
      {stage1_8[343], stage1_8[344], stage1_8[345], stage1_8[346], stage1_8[347], stage1_8[348]},
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage2_12[26],stage2_11[39],stage2_10[68],stage2_9[83],stage2_8[97]}
   );
   gpc606_5 gpc2422 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[27],stage2_11[40],stage2_10[69],stage2_9[84]}
   );
   gpc606_5 gpc2423 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[28],stage2_11[41],stage2_10[70],stage2_9[85]}
   );
   gpc606_5 gpc2424 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[29],stage2_11[42],stage2_10[71],stage2_9[86]}
   );
   gpc606_5 gpc2425 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[30],stage2_11[43],stage2_10[72],stage2_9[87]}
   );
   gpc606_5 gpc2426 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[31],stage2_11[44],stage2_10[73],stage2_9[88]}
   );
   gpc606_5 gpc2427 (
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[32],stage2_11[45],stage2_10[74],stage2_9[89]}
   );
   gpc606_5 gpc2428 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[33],stage2_11[46],stage2_10[75],stage2_9[90]}
   );
   gpc606_5 gpc2429 (
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[34],stage2_11[47],stage2_10[76],stage2_9[91]}
   );
   gpc606_5 gpc2430 (
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[35],stage2_11[48],stage2_10[77],stage2_9[92]}
   );
   gpc606_5 gpc2431 (
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[36],stage2_11[49],stage2_10[78],stage2_9[93]}
   );
   gpc606_5 gpc2432 (
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[37],stage2_11[50],stage2_10[79],stage2_9[94]}
   );
   gpc606_5 gpc2433 (
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[38],stage2_11[51],stage2_10[80],stage2_9[95]}
   );
   gpc606_5 gpc2434 (
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[39],stage2_11[52],stage2_10[81],stage2_9[96]}
   );
   gpc606_5 gpc2435 (
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[40],stage2_11[53],stage2_10[82],stage2_9[97]}
   );
   gpc606_5 gpc2436 (
      {stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[41],stage2_11[54],stage2_10[83],stage2_9[98]}
   );
   gpc606_5 gpc2437 (
      {stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[42],stage2_11[55],stage2_10[84],stage2_9[99]}
   );
   gpc606_5 gpc2438 (
      {stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[43],stage2_11[56],stage2_10[85],stage2_9[100]}
   );
   gpc606_5 gpc2439 (
      {stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[44],stage2_11[57],stage2_10[86],stage2_9[101]}
   );
   gpc606_5 gpc2440 (
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191]},
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage2_13[18],stage2_12[45],stage2_11[58],stage2_10[87],stage2_9[102]}
   );
   gpc606_5 gpc2441 (
      {stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197]},
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage2_13[19],stage2_12[46],stage2_11[59],stage2_10[88],stage2_9[103]}
   );
   gpc606_5 gpc2442 (
      {stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203]},
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125]},
      {stage2_13[20],stage2_12[47],stage2_11[60],stage2_10[89],stage2_9[104]}
   );
   gpc606_5 gpc2443 (
      {stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209]},
      {stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131]},
      {stage2_13[21],stage2_12[48],stage2_11[61],stage2_10[90],stage2_9[105]}
   );
   gpc615_5 gpc2444 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166]},
      {stage1_11[132]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[22],stage2_12[49],stage2_11[62],stage2_10[91]}
   );
   gpc615_5 gpc2445 (
      {stage1_10[167], stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171]},
      {stage1_11[133]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[23],stage2_12[50],stage2_11[63],stage2_10[92]}
   );
   gpc615_5 gpc2446 (
      {stage1_10[172], stage1_10[173], stage1_10[174], stage1_10[175], stage1_10[176]},
      {stage1_11[134]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[24],stage2_12[51],stage2_11[64],stage2_10[93]}
   );
   gpc615_5 gpc2447 (
      {stage1_10[177], stage1_10[178], stage1_10[179], stage1_10[180], stage1_10[181]},
      {stage1_11[135]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[25],stage2_12[52],stage2_11[65],stage2_10[94]}
   );
   gpc615_5 gpc2448 (
      {stage1_11[136], stage1_11[137], stage1_11[138], stage1_11[139], stage1_11[140]},
      {stage1_12[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[4],stage2_13[26],stage2_12[53],stage2_11[66]}
   );
   gpc615_5 gpc2449 (
      {stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144], stage1_11[145]},
      {stage1_12[25]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[5],stage2_13[27],stage2_12[54],stage2_11[67]}
   );
   gpc615_5 gpc2450 (
      {stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149], stage1_11[150]},
      {stage1_12[26]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[6],stage2_13[28],stage2_12[55],stage2_11[68]}
   );
   gpc615_5 gpc2451 (
      {stage1_11[151], stage1_11[152], stage1_11[153], stage1_11[154], stage1_11[155]},
      {stage1_12[27]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[7],stage2_13[29],stage2_12[56],stage2_11[69]}
   );
   gpc615_5 gpc2452 (
      {stage1_11[156], stage1_11[157], stage1_11[158], stage1_11[159], stage1_11[160]},
      {stage1_12[28]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[8],stage2_13[30],stage2_12[57],stage2_11[70]}
   );
   gpc606_5 gpc2453 (
      {stage1_12[29], stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[5],stage2_14[9],stage2_13[31],stage2_12[58]}
   );
   gpc615_5 gpc2454 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39]},
      {stage1_13[30]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[6],stage2_14[10],stage2_13[32],stage2_12[59]}
   );
   gpc615_5 gpc2455 (
      {stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43], stage1_12[44]},
      {stage1_13[31]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[7],stage2_14[11],stage2_13[33],stage2_12[60]}
   );
   gpc615_5 gpc2456 (
      {stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage1_13[32]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[8],stage2_14[12],stage2_13[34],stage2_12[61]}
   );
   gpc615_5 gpc2457 (
      {stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53], stage1_12[54]},
      {stage1_13[33]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[9],stage2_14[13],stage2_13[35],stage2_12[62]}
   );
   gpc615_5 gpc2458 (
      {stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_13[34]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[10],stage2_14[14],stage2_13[36],stage2_12[63]}
   );
   gpc615_5 gpc2459 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64]},
      {stage1_13[35]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[11],stage2_14[15],stage2_13[37],stage2_12[64]}
   );
   gpc615_5 gpc2460 (
      {stage1_12[65], stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69]},
      {stage1_13[36]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[12],stage2_14[16],stage2_13[38],stage2_12[65]}
   );
   gpc615_5 gpc2461 (
      {stage1_12[70], stage1_12[71], stage1_12[72], stage1_12[73], stage1_12[74]},
      {stage1_13[37]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[13],stage2_14[17],stage2_13[39],stage2_12[66]}
   );
   gpc615_5 gpc2462 (
      {stage1_12[75], stage1_12[76], stage1_12[77], stage1_12[78], stage1_12[79]},
      {stage1_13[38]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[14],stage2_14[18],stage2_13[40],stage2_12[67]}
   );
   gpc615_5 gpc2463 (
      {stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83], stage1_12[84]},
      {stage1_13[39]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[15],stage2_14[19],stage2_13[41],stage2_12[68]}
   );
   gpc615_5 gpc2464 (
      {stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage1_13[40]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[16],stage2_14[20],stage2_13[42],stage2_12[69]}
   );
   gpc615_5 gpc2465 (
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94]},
      {stage1_13[41]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[17],stage2_14[21],stage2_13[43],stage2_12[70]}
   );
   gpc615_5 gpc2466 (
      {stage1_12[95], stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99]},
      {stage1_13[42]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[18],stage2_14[22],stage2_13[44],stage2_12[71]}
   );
   gpc615_5 gpc2467 (
      {stage1_12[100], stage1_12[101], stage1_12[102], stage1_12[103], stage1_12[104]},
      {stage1_13[43]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[19],stage2_14[23],stage2_13[45],stage2_12[72]}
   );
   gpc615_5 gpc2468 (
      {stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108], stage1_12[109]},
      {stage1_13[44]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[20],stage2_14[24],stage2_13[46],stage2_12[73]}
   );
   gpc615_5 gpc2469 (
      {stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_13[45]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[21],stage2_14[25],stage2_13[47],stage2_12[74]}
   );
   gpc615_5 gpc2470 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_13[46]},
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage2_16[17],stage2_15[22],stage2_14[26],stage2_13[48],stage2_12[75]}
   );
   gpc615_5 gpc2471 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124]},
      {stage1_13[47]},
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage2_16[18],stage2_15[23],stage2_14[27],stage2_13[49],stage2_12[76]}
   );
   gpc615_5 gpc2472 (
      {stage1_12[125], stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129]},
      {stage1_13[48]},
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage2_16[19],stage2_15[24],stage2_14[28],stage2_13[50],stage2_12[77]}
   );
   gpc615_5 gpc2473 (
      {stage1_12[130], stage1_12[131], stage1_12[132], stage1_12[133], stage1_12[134]},
      {stage1_13[49]},
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage2_16[20],stage2_15[25],stage2_14[29],stage2_13[51],stage2_12[78]}
   );
   gpc615_5 gpc2474 (
      {stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138], stage1_12[139]},
      {stage1_13[50]},
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage2_16[21],stage2_15[26],stage2_14[30],stage2_13[52],stage2_12[79]}
   );
   gpc615_5 gpc2475 (
      {stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_13[51]},
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage2_16[22],stage2_15[27],stage2_14[31],stage2_13[53],stage2_12[80]}
   );
   gpc615_5 gpc2476 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149]},
      {stage1_13[52]},
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage2_16[23],stage2_15[28],stage2_14[32],stage2_13[54],stage2_12[81]}
   );
   gpc615_5 gpc2477 (
      {stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154]},
      {stage1_13[53]},
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149]},
      {stage2_16[24],stage2_15[29],stage2_14[33],stage2_13[55],stage2_12[82]}
   );
   gpc615_5 gpc2478 (
      {stage1_12[155], stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159]},
      {stage1_13[54]},
      {stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155]},
      {stage2_16[25],stage2_15[30],stage2_14[34],stage2_13[56],stage2_12[83]}
   );
   gpc615_5 gpc2479 (
      {stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_13[55]},
      {stage1_14[156], stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage2_16[26],stage2_15[31],stage2_14[35],stage2_13[57],stage2_12[84]}
   );
   gpc615_5 gpc2480 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169]},
      {stage1_13[56]},
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167]},
      {stage2_16[27],stage2_15[32],stage2_14[36],stage2_13[58],stage2_12[85]}
   );
   gpc615_5 gpc2481 (
      {stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174]},
      {stage1_13[57]},
      {stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage2_16[28],stage2_15[33],stage2_14[37],stage2_13[59],stage2_12[86]}
   );
   gpc615_5 gpc2482 (
      {stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179]},
      {stage1_13[58]},
      {stage1_14[174], stage1_14[175], stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179]},
      {stage2_16[29],stage2_15[34],stage2_14[38],stage2_13[60],stage2_12[87]}
   );
   gpc615_5 gpc2483 (
      {stage1_12[180], stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184]},
      {stage1_13[59]},
      {stage1_14[180], stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage2_16[30],stage2_15[35],stage2_14[39],stage2_13[61],stage2_12[88]}
   );
   gpc615_5 gpc2484 (
      {stage1_12[185], stage1_12[186], stage1_12[187], stage1_12[188], stage1_12[189]},
      {stage1_13[60]},
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage2_16[31],stage2_15[36],stage2_14[40],stage2_13[62],stage2_12[89]}
   );
   gpc615_5 gpc2485 (
      {stage1_12[190], stage1_12[191], stage1_12[192], stage1_12[193], stage1_12[194]},
      {stage1_13[61]},
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197]},
      {stage2_16[32],stage2_15[37],stage2_14[41],stage2_13[63],stage2_12[90]}
   );
   gpc615_5 gpc2486 (
      {stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198], stage1_12[199]},
      {stage1_13[62]},
      {stage1_14[198], stage1_14[199], stage1_14[200], stage1_14[201], stage1_14[202], stage1_14[203]},
      {stage2_16[33],stage2_15[38],stage2_14[42],stage2_13[64],stage2_12[91]}
   );
   gpc615_5 gpc2487 (
      {stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203], stage1_12[204]},
      {stage1_13[63]},
      {stage1_14[204], stage1_14[205], stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209]},
      {stage2_16[34],stage2_15[39],stage2_14[43],stage2_13[65],stage2_12[92]}
   );
   gpc615_5 gpc2488 (
      {stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209]},
      {stage1_13[64]},
      {stage1_14[210], stage1_14[211], stage1_14[212], stage1_14[213], stage1_14[214], stage1_14[215]},
      {stage2_16[35],stage2_15[40],stage2_14[44],stage2_13[66],stage2_12[93]}
   );
   gpc615_5 gpc2489 (
      {stage1_12[210], stage1_12[211], stage1_12[212], stage1_12[213], stage1_12[214]},
      {stage1_13[65]},
      {stage1_14[216], stage1_14[217], stage1_14[218], stage1_14[219], stage1_14[220], stage1_14[221]},
      {stage2_16[36],stage2_15[41],stage2_14[45],stage2_13[67],stage2_12[94]}
   );
   gpc606_5 gpc2490 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[37],stage2_15[42],stage2_14[46],stage2_13[68]}
   );
   gpc606_5 gpc2491 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[38],stage2_15[43],stage2_14[47],stage2_13[69]}
   );
   gpc606_5 gpc2492 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[39],stage2_15[44],stage2_14[48],stage2_13[70]}
   );
   gpc606_5 gpc2493 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[40],stage2_15[45],stage2_14[49],stage2_13[71]}
   );
   gpc606_5 gpc2494 (
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[41],stage2_15[46],stage2_14[50],stage2_13[72]}
   );
   gpc606_5 gpc2495 (
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[42],stage2_15[47],stage2_14[51],stage2_13[73]}
   );
   gpc606_5 gpc2496 (
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[43],stage2_15[48],stage2_14[52],stage2_13[74]}
   );
   gpc606_5 gpc2497 (
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[44],stage2_15[49],stage2_14[53],stage2_13[75]}
   );
   gpc606_5 gpc2498 (
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[45],stage2_15[50],stage2_14[54],stage2_13[76]}
   );
   gpc606_5 gpc2499 (
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[46],stage2_15[51],stage2_14[55],stage2_13[77]}
   );
   gpc606_5 gpc2500 (
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[47],stage2_15[52],stage2_14[56],stage2_13[78]}
   );
   gpc606_5 gpc2501 (
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[48],stage2_15[53],stage2_14[57],stage2_13[79]}
   );
   gpc606_5 gpc2502 (
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[49],stage2_15[54],stage2_14[58],stage2_13[80]}
   );
   gpc606_5 gpc2503 (
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[50],stage2_15[55],stage2_14[59],stage2_13[81]}
   );
   gpc606_5 gpc2504 (
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[51],stage2_15[56],stage2_14[60],stage2_13[82]}
   );
   gpc606_5 gpc2505 (
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[52],stage2_15[57],stage2_14[61],stage2_13[83]}
   );
   gpc606_5 gpc2506 (
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[53],stage2_15[58],stage2_14[62],stage2_13[84]}
   );
   gpc606_5 gpc2507 (
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[54],stage2_15[59],stage2_14[63],stage2_13[85]}
   );
   gpc606_5 gpc2508 (
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[55],stage2_15[60],stage2_14[64],stage2_13[86]}
   );
   gpc606_5 gpc2509 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage2_17[19],stage2_16[56],stage2_15[61],stage2_14[65],stage2_13[87]}
   );
   gpc606_5 gpc2510 (
      {stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage2_17[20],stage2_16[57],stage2_15[62],stage2_14[66],stage2_13[88]}
   );
   gpc606_5 gpc2511 (
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196], stage1_13[197]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage2_17[21],stage2_16[58],stage2_15[63],stage2_14[67],stage2_13[89]}
   );
   gpc615_5 gpc2512 (
      {stage1_14[222], stage1_14[223], stage1_14[224], stage1_14[225], stage1_14[226]},
      {stage1_15[132]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[22],stage2_16[59],stage2_15[64],stage2_14[68]}
   );
   gpc615_5 gpc2513 (
      {stage1_14[227], stage1_14[228], stage1_14[229], stage1_14[230], stage1_14[231]},
      {stage1_15[133]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[23],stage2_16[60],stage2_15[65],stage2_14[69]}
   );
   gpc606_5 gpc2514 (
      {stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137], stage1_15[138], stage1_15[139]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[24],stage2_16[61],stage2_15[66]}
   );
   gpc606_5 gpc2515 (
      {stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143], stage1_15[144], stage1_15[145]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[25],stage2_16[62],stage2_15[67]}
   );
   gpc606_5 gpc2516 (
      {stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149], stage1_15[150], stage1_15[151]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[26],stage2_16[63],stage2_15[68]}
   );
   gpc615_5 gpc2517 (
      {stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155], stage1_15[156]},
      {stage1_16[12]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[27],stage2_16[64],stage2_15[69]}
   );
   gpc615_5 gpc2518 (
      {stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage1_16[13]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[28],stage2_16[65],stage2_15[70]}
   );
   gpc615_5 gpc2519 (
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166]},
      {stage1_16[14]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[7],stage2_17[29],stage2_16[66],stage2_15[71]}
   );
   gpc615_5 gpc2520 (
      {stage1_15[167], stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171]},
      {stage1_16[15]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[8],stage2_17[30],stage2_16[67],stage2_15[72]}
   );
   gpc615_5 gpc2521 (
      {stage1_15[172], stage1_15[173], stage1_15[174], stage1_15[175], stage1_15[176]},
      {stage1_16[16]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[9],stage2_17[31],stage2_16[68],stage2_15[73]}
   );
   gpc615_5 gpc2522 (
      {stage1_15[177], stage1_15[178], stage1_15[179], stage1_15[180], stage1_15[181]},
      {stage1_16[17]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[10],stage2_17[32],stage2_16[69],stage2_15[74]}
   );
   gpc615_5 gpc2523 (
      {stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185], stage1_15[186]},
      {stage1_16[18]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[11],stage2_17[33],stage2_16[70],stage2_15[75]}
   );
   gpc615_5 gpc2524 (
      {stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage1_16[19]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[12],stage2_17[34],stage2_16[71],stage2_15[76]}
   );
   gpc615_5 gpc2525 (
      {stage1_15[192], stage1_15[193], stage1_15[194], stage1_15[195], stage1_15[196]},
      {stage1_16[20]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[13],stage2_17[35],stage2_16[72],stage2_15[77]}
   );
   gpc615_5 gpc2526 (
      {stage1_15[197], stage1_15[198], stage1_15[199], stage1_15[200], stage1_15[201]},
      {stage1_16[21]},
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage2_19[12],stage2_18[14],stage2_17[36],stage2_16[73],stage2_15[78]}
   );
   gpc615_5 gpc2527 (
      {stage1_15[202], stage1_15[203], stage1_15[204], stage1_15[205], stage1_15[206]},
      {stage1_16[22]},
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage2_19[13],stage2_18[15],stage2_17[37],stage2_16[74],stage2_15[79]}
   );
   gpc615_5 gpc2528 (
      {stage1_15[207], stage1_15[208], stage1_15[209], stage1_15[210], stage1_15[211]},
      {stage1_16[23]},
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage2_19[14],stage2_18[16],stage2_17[38],stage2_16[75],stage2_15[80]}
   );
   gpc615_5 gpc2529 (
      {stage1_15[212], stage1_15[213], stage1_15[214], stage1_15[215], stage1_15[216]},
      {stage1_16[24]},
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage2_19[15],stage2_18[17],stage2_17[39],stage2_16[76],stage2_15[81]}
   );
   gpc615_5 gpc2530 (
      {stage1_15[217], stage1_15[218], stage1_15[219], stage1_15[220], stage1_15[221]},
      {stage1_16[25]},
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage2_19[16],stage2_18[18],stage2_17[40],stage2_16[77],stage2_15[82]}
   );
   gpc606_5 gpc2531 (
      {stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29], stage1_16[30], stage1_16[31]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[17],stage2_18[19],stage2_17[41],stage2_16[78]}
   );
   gpc606_5 gpc2532 (
      {stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35], stage1_16[36], stage1_16[37]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[18],stage2_18[20],stage2_17[42],stage2_16[79]}
   );
   gpc606_5 gpc2533 (
      {stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[19],stage2_18[21],stage2_17[43],stage2_16[80]}
   );
   gpc606_5 gpc2534 (
      {stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[20],stage2_18[22],stage2_17[44],stage2_16[81]}
   );
   gpc606_5 gpc2535 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[21],stage2_18[23],stage2_17[45],stage2_16[82]}
   );
   gpc606_5 gpc2536 (
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[22],stage2_18[24],stage2_17[46],stage2_16[83]}
   );
   gpc606_5 gpc2537 (
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[23],stage2_18[25],stage2_17[47],stage2_16[84]}
   );
   gpc606_5 gpc2538 (
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[24],stage2_18[26],stage2_17[48],stage2_16[85]}
   );
   gpc606_5 gpc2539 (
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[25],stage2_18[27],stage2_17[49],stage2_16[86]}
   );
   gpc606_5 gpc2540 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[26],stage2_18[28],stage2_17[50],stage2_16[87]}
   );
   gpc606_5 gpc2541 (
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[27],stage2_18[29],stage2_17[51],stage2_16[88]}
   );
   gpc606_5 gpc2542 (
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[28],stage2_18[30],stage2_17[52],stage2_16[89]}
   );
   gpc606_5 gpc2543 (
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[29],stage2_18[31],stage2_17[53],stage2_16[90]}
   );
   gpc606_5 gpc2544 (
      {stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107], stage1_16[108], stage1_16[109]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[30],stage2_18[32],stage2_17[54],stage2_16[91]}
   );
   gpc606_5 gpc2545 (
      {stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113], stage1_16[114], stage1_16[115]},
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage2_20[14],stage2_19[31],stage2_18[33],stage2_17[55],stage2_16[92]}
   );
   gpc606_5 gpc2546 (
      {stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119], stage1_16[120], stage1_16[121]},
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage2_20[15],stage2_19[32],stage2_18[34],stage2_17[56],stage2_16[93]}
   );
   gpc606_5 gpc2547 (
      {stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125], stage1_16[126], stage1_16[127]},
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage2_20[16],stage2_19[33],stage2_18[35],stage2_17[57],stage2_16[94]}
   );
   gpc606_5 gpc2548 (
      {stage1_16[128], stage1_16[129], stage1_16[130], stage1_16[131], stage1_16[132], stage1_16[133]},
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage2_20[17],stage2_19[34],stage2_18[36],stage2_17[58],stage2_16[95]}
   );
   gpc606_5 gpc2549 (
      {stage1_16[134], stage1_16[135], stage1_16[136], stage1_16[137], stage1_16[138], stage1_16[139]},
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage2_20[18],stage2_19[35],stage2_18[37],stage2_17[59],stage2_16[96]}
   );
   gpc606_5 gpc2550 (
      {stage1_16[140], stage1_16[141], stage1_16[142], stage1_16[143], stage1_16[144], stage1_16[145]},
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage2_20[19],stage2_19[36],stage2_18[38],stage2_17[60],stage2_16[97]}
   );
   gpc606_5 gpc2551 (
      {stage1_16[146], stage1_16[147], stage1_16[148], stage1_16[149], stage1_16[150], stage1_16[151]},
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage2_20[20],stage2_19[37],stage2_18[39],stage2_17[61],stage2_16[98]}
   );
   gpc606_5 gpc2552 (
      {stage1_16[152], stage1_16[153], stage1_16[154], stage1_16[155], stage1_16[156], stage1_16[157]},
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage2_20[21],stage2_19[38],stage2_18[40],stage2_17[62],stage2_16[99]}
   );
   gpc606_5 gpc2553 (
      {stage1_16[158], stage1_16[159], stage1_16[160], stage1_16[161], stage1_16[162], stage1_16[163]},
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage2_20[22],stage2_19[39],stage2_18[41],stage2_17[63],stage2_16[100]}
   );
   gpc606_5 gpc2554 (
      {stage1_16[164], stage1_16[165], stage1_16[166], stage1_16[167], stage1_16[168], stage1_16[169]},
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage2_20[23],stage2_19[40],stage2_18[42],stage2_17[64],stage2_16[101]}
   );
   gpc606_5 gpc2555 (
      {stage1_16[170], stage1_16[171], stage1_16[172], stage1_16[173], stage1_16[174], stage1_16[175]},
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage2_20[24],stage2_19[41],stage2_18[43],stage2_17[65],stage2_16[102]}
   );
   gpc615_5 gpc2556 (
      {stage1_16[176], stage1_16[177], stage1_16[178], stage1_16[179], stage1_16[180]},
      {stage1_17[102]},
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage2_20[25],stage2_19[42],stage2_18[44],stage2_17[66],stage2_16[103]}
   );
   gpc615_5 gpc2557 (
      {stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184], stage1_16[185]},
      {stage1_17[103]},
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage2_20[26],stage2_19[43],stage2_18[45],stage2_17[67],stage2_16[104]}
   );
   gpc615_5 gpc2558 (
      {stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190]},
      {stage1_17[104]},
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage2_20[27],stage2_19[44],stage2_18[46],stage2_17[68],stage2_16[105]}
   );
   gpc615_5 gpc2559 (
      {stage1_16[191], stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195]},
      {stage1_17[105]},
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage2_20[28],stage2_19[45],stage2_18[47],stage2_17[69],stage2_16[106]}
   );
   gpc606_5 gpc2560 (
      {stage1_17[106], stage1_17[107], stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[29],stage2_19[46],stage2_18[48],stage2_17[70]}
   );
   gpc606_5 gpc2561 (
      {stage1_17[112], stage1_17[113], stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[30],stage2_19[47],stage2_18[49],stage2_17[71]}
   );
   gpc606_5 gpc2562 (
      {stage1_17[118], stage1_17[119], stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[31],stage2_19[48],stage2_18[50],stage2_17[72]}
   );
   gpc606_5 gpc2563 (
      {stage1_17[124], stage1_17[125], stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[32],stage2_19[49],stage2_18[51],stage2_17[73]}
   );
   gpc606_5 gpc2564 (
      {stage1_17[130], stage1_17[131], stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[33],stage2_19[50],stage2_18[52],stage2_17[74]}
   );
   gpc606_5 gpc2565 (
      {stage1_17[136], stage1_17[137], stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[34],stage2_19[51],stage2_18[53],stage2_17[75]}
   );
   gpc606_5 gpc2566 (
      {stage1_17[142], stage1_17[143], stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[35],stage2_19[52],stage2_18[54],stage2_17[76]}
   );
   gpc606_5 gpc2567 (
      {stage1_17[148], stage1_17[149], stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[36],stage2_19[53],stage2_18[55],stage2_17[77]}
   );
   gpc606_5 gpc2568 (
      {stage1_17[154], stage1_17[155], stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[37],stage2_19[54],stage2_18[56],stage2_17[78]}
   );
   gpc606_5 gpc2569 (
      {stage1_17[160], stage1_17[161], stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[38],stage2_19[55],stage2_18[57],stage2_17[79]}
   );
   gpc606_5 gpc2570 (
      {stage1_17[166], stage1_17[167], stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[39],stage2_19[56],stage2_18[58],stage2_17[80]}
   );
   gpc606_5 gpc2571 (
      {stage1_17[172], stage1_17[173], stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[40],stage2_19[57],stage2_18[59],stage2_17[81]}
   );
   gpc615_5 gpc2572 (
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178]},
      {stage1_19[72]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[12],stage2_20[41],stage2_19[58],stage2_18[60]}
   );
   gpc615_5 gpc2573 (
      {stage1_18[179], stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183]},
      {stage1_19[73]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[13],stage2_20[42],stage2_19[59],stage2_18[61]}
   );
   gpc615_5 gpc2574 (
      {stage1_18[184], stage1_18[185], stage1_18[186], stage1_18[187], stage1_18[188]},
      {stage1_19[74]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[14],stage2_20[43],stage2_19[60],stage2_18[62]}
   );
   gpc615_5 gpc2575 (
      {stage1_18[189], stage1_18[190], stage1_18[191], stage1_18[192], stage1_18[193]},
      {stage1_19[75]},
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage2_22[3],stage2_21[15],stage2_20[44],stage2_19[61],stage2_18[63]}
   );
   gpc606_5 gpc2576 (
      {stage1_19[76], stage1_19[77], stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[4],stage2_21[16],stage2_20[45],stage2_19[62]}
   );
   gpc606_5 gpc2577 (
      {stage1_19[82], stage1_19[83], stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[5],stage2_21[17],stage2_20[46],stage2_19[63]}
   );
   gpc606_5 gpc2578 (
      {stage1_19[88], stage1_19[89], stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[6],stage2_21[18],stage2_20[47],stage2_19[64]}
   );
   gpc606_5 gpc2579 (
      {stage1_19[94], stage1_19[95], stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[7],stage2_21[19],stage2_20[48],stage2_19[65]}
   );
   gpc606_5 gpc2580 (
      {stage1_19[100], stage1_19[101], stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[8],stage2_21[20],stage2_20[49],stage2_19[66]}
   );
   gpc606_5 gpc2581 (
      {stage1_19[106], stage1_19[107], stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[9],stage2_21[21],stage2_20[50],stage2_19[67]}
   );
   gpc606_5 gpc2582 (
      {stage1_19[112], stage1_19[113], stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[10],stage2_21[22],stage2_20[51],stage2_19[68]}
   );
   gpc606_5 gpc2583 (
      {stage1_19[118], stage1_19[119], stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[11],stage2_21[23],stage2_20[52],stage2_19[69]}
   );
   gpc606_5 gpc2584 (
      {stage1_19[124], stage1_19[125], stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[12],stage2_21[24],stage2_20[53],stage2_19[70]}
   );
   gpc606_5 gpc2585 (
      {stage1_19[130], stage1_19[131], stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[13],stage2_21[25],stage2_20[54],stage2_19[71]}
   );
   gpc606_5 gpc2586 (
      {stage1_19[136], stage1_19[137], stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[14],stage2_21[26],stage2_20[55],stage2_19[72]}
   );
   gpc606_5 gpc2587 (
      {stage1_19[142], stage1_19[143], stage1_19[144], stage1_19[145], stage1_19[146], stage1_19[147]},
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage2_23[11],stage2_22[15],stage2_21[27],stage2_20[56],stage2_19[73]}
   );
   gpc606_5 gpc2588 (
      {stage1_19[148], stage1_19[149], stage1_19[150], stage1_19[151], stage1_19[152], stage1_19[153]},
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage2_23[12],stage2_22[16],stage2_21[28],stage2_20[57],stage2_19[74]}
   );
   gpc606_5 gpc2589 (
      {stage1_19[154], stage1_19[155], stage1_19[156], stage1_19[157], stage1_19[158], stage1_19[159]},
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage2_23[13],stage2_22[17],stage2_21[29],stage2_20[58],stage2_19[75]}
   );
   gpc606_5 gpc2590 (
      {stage1_19[160], stage1_19[161], stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165]},
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage2_23[14],stage2_22[18],stage2_21[30],stage2_20[59],stage2_19[76]}
   );
   gpc615_5 gpc2591 (
      {stage1_19[166], stage1_19[167], stage1_19[168], stage1_19[169], stage1_19[170]},
      {stage1_20[24]},
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage2_23[15],stage2_22[19],stage2_21[31],stage2_20[60],stage2_19[77]}
   );
   gpc615_5 gpc2592 (
      {stage1_19[171], stage1_19[172], stage1_19[173], stage1_19[174], stage1_19[175]},
      {stage1_20[25]},
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage2_23[16],stage2_22[20],stage2_21[32],stage2_20[61],stage2_19[78]}
   );
   gpc615_5 gpc2593 (
      {stage1_19[176], stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180]},
      {stage1_20[26]},
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage2_23[17],stage2_22[21],stage2_21[33],stage2_20[62],stage2_19[79]}
   );
   gpc615_5 gpc2594 (
      {stage1_19[181], stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185]},
      {stage1_20[27]},
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage2_23[18],stage2_22[22],stage2_21[34],stage2_20[63],stage2_19[80]}
   );
   gpc615_5 gpc2595 (
      {stage1_19[186], stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190]},
      {stage1_20[28]},
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage2_23[19],stage2_22[23],stage2_21[35],stage2_20[64],stage2_19[81]}
   );
   gpc615_5 gpc2596 (
      {stage1_19[191], stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195]},
      {stage1_20[29]},
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage2_23[20],stage2_22[24],stage2_21[36],stage2_20[65],stage2_19[82]}
   );
   gpc615_5 gpc2597 (
      {stage1_19[196], stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200]},
      {stage1_20[30]},
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage2_23[21],stage2_22[25],stage2_21[37],stage2_20[66],stage2_19[83]}
   );
   gpc615_5 gpc2598 (
      {stage1_19[201], stage1_19[202], stage1_19[203], stage1_19[204], stage1_19[205]},
      {stage1_20[31]},
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage2_23[22],stage2_22[26],stage2_21[38],stage2_20[67],stage2_19[84]}
   );
   gpc615_5 gpc2599 (
      {stage1_19[206], stage1_19[207], stage1_19[208], stage1_19[209], stage1_19[210]},
      {stage1_20[32]},
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage2_23[23],stage2_22[27],stage2_21[39],stage2_20[68],stage2_19[85]}
   );
   gpc615_5 gpc2600 (
      {stage1_19[211], stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215]},
      {stage1_20[33]},
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage2_23[24],stage2_22[28],stage2_21[40],stage2_20[69],stage2_19[86]}
   );
   gpc615_5 gpc2601 (
      {stage1_19[216], stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220]},
      {stage1_20[34]},
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage2_23[25],stage2_22[29],stage2_21[41],stage2_20[70],stage2_19[87]}
   );
   gpc615_5 gpc2602 (
      {stage1_19[221], stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225]},
      {stage1_20[35]},
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage2_23[26],stage2_22[30],stage2_21[42],stage2_20[71],stage2_19[88]}
   );
   gpc615_5 gpc2603 (
      {stage1_19[226], stage1_19[227], stage1_19[228], stage1_19[229], stage1_19[230]},
      {stage1_20[36]},
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage2_23[27],stage2_22[31],stage2_21[43],stage2_20[72],stage2_19[89]}
   );
   gpc615_5 gpc2604 (
      {stage1_19[231], stage1_19[232], stage1_19[233], stage1_19[234], stage1_19[235]},
      {stage1_20[37]},
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage2_23[28],stage2_22[32],stage2_21[44],stage2_20[73],stage2_19[90]}
   );
   gpc615_5 gpc2605 (
      {stage1_19[236], stage1_19[237], stage1_19[238], stage1_19[239], stage1_19[240]},
      {stage1_20[38]},
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage2_23[29],stage2_22[33],stage2_21[45],stage2_20[74],stage2_19[91]}
   );
   gpc615_5 gpc2606 (
      {stage1_19[241], stage1_19[242], stage1_19[243], stage1_19[244], stage1_19[245]},
      {stage1_20[39]},
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage2_23[30],stage2_22[34],stage2_21[46],stage2_20[75],stage2_19[92]}
   );
   gpc615_5 gpc2607 (
      {stage1_19[246], stage1_19[247], stage1_19[248], stage1_19[249], stage1_19[250]},
      {stage1_20[40]},
      {stage1_21[186], stage1_21[187], stage1_21[188], stage1_21[189], stage1_21[190], stage1_21[191]},
      {stage2_23[31],stage2_22[35],stage2_21[47],stage2_20[76],stage2_19[93]}
   );
   gpc615_5 gpc2608 (
      {stage1_19[251], stage1_19[252], stage1_19[253], stage1_19[254], stage1_19[255]},
      {stage1_20[41]},
      {stage1_21[192], stage1_21[193], stage1_21[194], stage1_21[195], stage1_21[196], stage1_21[197]},
      {stage2_23[32],stage2_22[36],stage2_21[48],stage2_20[77],stage2_19[94]}
   );
   gpc615_5 gpc2609 (
      {stage1_19[256], stage1_19[257], stage1_19[258], stage1_19[259], stage1_19[260]},
      {stage1_20[42]},
      {stage1_21[198], stage1_21[199], stage1_21[200], stage1_21[201], stage1_21[202], stage1_21[203]},
      {stage2_23[33],stage2_22[37],stage2_21[49],stage2_20[78],stage2_19[95]}
   );
   gpc606_5 gpc2610 (
      {stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46], stage1_20[47], stage1_20[48]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[34],stage2_22[38],stage2_21[50],stage2_20[79]}
   );
   gpc606_5 gpc2611 (
      {stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52], stage1_20[53], stage1_20[54]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[35],stage2_22[39],stage2_21[51],stage2_20[80]}
   );
   gpc606_5 gpc2612 (
      {stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58], stage1_20[59], stage1_20[60]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[36],stage2_22[40],stage2_21[52],stage2_20[81]}
   );
   gpc606_5 gpc2613 (
      {stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64], stage1_20[65], stage1_20[66]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[37],stage2_22[41],stage2_21[53],stage2_20[82]}
   );
   gpc606_5 gpc2614 (
      {stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70], stage1_20[71], stage1_20[72]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[38],stage2_22[42],stage2_21[54],stage2_20[83]}
   );
   gpc606_5 gpc2615 (
      {stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76], stage1_20[77], stage1_20[78]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[39],stage2_22[43],stage2_21[55],stage2_20[84]}
   );
   gpc606_5 gpc2616 (
      {stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82], stage1_20[83], stage1_20[84]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[40],stage2_22[44],stage2_21[56],stage2_20[85]}
   );
   gpc606_5 gpc2617 (
      {stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88], stage1_20[89], stage1_20[90]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[41],stage2_22[45],stage2_21[57],stage2_20[86]}
   );
   gpc606_5 gpc2618 (
      {stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94], stage1_20[95], stage1_20[96]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[42],stage2_22[46],stage2_21[58],stage2_20[87]}
   );
   gpc606_5 gpc2619 (
      {stage1_20[97], stage1_20[98], stage1_20[99], stage1_20[100], stage1_20[101], stage1_20[102]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[43],stage2_22[47],stage2_21[59],stage2_20[88]}
   );
   gpc606_5 gpc2620 (
      {stage1_20[103], stage1_20[104], stage1_20[105], stage1_20[106], stage1_20[107], stage1_20[108]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[44],stage2_22[48],stage2_21[60],stage2_20[89]}
   );
   gpc606_5 gpc2621 (
      {stage1_20[109], stage1_20[110], stage1_20[111], stage1_20[112], stage1_20[113], stage1_20[114]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[45],stage2_22[49],stage2_21[61],stage2_20[90]}
   );
   gpc606_5 gpc2622 (
      {stage1_20[115], stage1_20[116], stage1_20[117], stage1_20[118], stage1_20[119], stage1_20[120]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[46],stage2_22[50],stage2_21[62],stage2_20[91]}
   );
   gpc606_5 gpc2623 (
      {stage1_20[121], stage1_20[122], stage1_20[123], stage1_20[124], stage1_20[125], stage1_20[126]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[47],stage2_22[51],stage2_21[63],stage2_20[92]}
   );
   gpc606_5 gpc2624 (
      {stage1_20[127], stage1_20[128], stage1_20[129], stage1_20[130], stage1_20[131], stage1_20[132]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[48],stage2_22[52],stage2_21[64],stage2_20[93]}
   );
   gpc606_5 gpc2625 (
      {stage1_20[133], stage1_20[134], stage1_20[135], stage1_20[136], stage1_20[137], stage1_20[138]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[49],stage2_22[53],stage2_21[65],stage2_20[94]}
   );
   gpc606_5 gpc2626 (
      {stage1_20[139], stage1_20[140], stage1_20[141], stage1_20[142], stage1_20[143], stage1_20[144]},
      {stage1_22[96], stage1_22[97], stage1_22[98], stage1_22[99], stage1_22[100], stage1_22[101]},
      {stage2_24[16],stage2_23[50],stage2_22[54],stage2_21[66],stage2_20[95]}
   );
   gpc606_5 gpc2627 (
      {stage1_20[145], stage1_20[146], stage1_20[147], stage1_20[148], stage1_20[149], stage1_20[150]},
      {stage1_22[102], stage1_22[103], stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107]},
      {stage2_24[17],stage2_23[51],stage2_22[55],stage2_21[67],stage2_20[96]}
   );
   gpc606_5 gpc2628 (
      {stage1_20[151], stage1_20[152], stage1_20[153], stage1_20[154], stage1_20[155], stage1_20[156]},
      {stage1_22[108], stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage2_24[18],stage2_23[52],stage2_22[56],stage2_21[68],stage2_20[97]}
   );
   gpc606_5 gpc2629 (
      {stage1_20[157], stage1_20[158], stage1_20[159], stage1_20[160], stage1_20[161], stage1_20[162]},
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage2_24[19],stage2_23[53],stage2_22[57],stage2_21[69],stage2_20[98]}
   );
   gpc606_5 gpc2630 (
      {stage1_20[163], stage1_20[164], stage1_20[165], stage1_20[166], stage1_20[167], stage1_20[168]},
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124], stage1_22[125]},
      {stage2_24[20],stage2_23[54],stage2_22[58],stage2_21[70],stage2_20[99]}
   );
   gpc606_5 gpc2631 (
      {stage1_20[169], stage1_20[170], stage1_20[171], stage1_20[172], stage1_20[173], stage1_20[174]},
      {stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129], stage1_22[130], stage1_22[131]},
      {stage2_24[21],stage2_23[55],stage2_22[59],stage2_21[71],stage2_20[100]}
   );
   gpc606_5 gpc2632 (
      {stage1_20[175], stage1_20[176], stage1_20[177], stage1_20[178], stage1_20[179], stage1_20[180]},
      {stage1_22[132], stage1_22[133], stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137]},
      {stage2_24[22],stage2_23[56],stage2_22[60],stage2_21[72],stage2_20[101]}
   );
   gpc606_5 gpc2633 (
      {stage1_20[181], stage1_20[182], stage1_20[183], stage1_20[184], stage1_20[185], stage1_20[186]},
      {stage1_22[138], stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142], stage1_22[143]},
      {stage2_24[23],stage2_23[57],stage2_22[61],stage2_21[73],stage2_20[102]}
   );
   gpc606_5 gpc2634 (
      {stage1_20[187], stage1_20[188], stage1_20[189], stage1_20[190], stage1_20[191], stage1_20[192]},
      {stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147], stage1_22[148], stage1_22[149]},
      {stage2_24[24],stage2_23[58],stage2_22[62],stage2_21[74],stage2_20[103]}
   );
   gpc606_5 gpc2635 (
      {stage1_20[193], stage1_20[194], stage1_20[195], stage1_20[196], stage1_20[197], stage1_20[198]},
      {stage1_22[150], stage1_22[151], stage1_22[152], stage1_22[153], stage1_22[154], stage1_22[155]},
      {stage2_24[25],stage2_23[59],stage2_22[63],stage2_21[75],stage2_20[104]}
   );
   gpc606_5 gpc2636 (
      {stage1_20[199], stage1_20[200], stage1_20[201], stage1_20[202], stage1_20[203], stage1_20[204]},
      {stage1_22[156], stage1_22[157], stage1_22[158], stage1_22[159], stage1_22[160], stage1_22[161]},
      {stage2_24[26],stage2_23[60],stage2_22[64],stage2_21[76],stage2_20[105]}
   );
   gpc606_5 gpc2637 (
      {stage1_20[205], stage1_20[206], stage1_20[207], stage1_20[208], stage1_20[209], stage1_20[210]},
      {stage1_22[162], stage1_22[163], stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167]},
      {stage2_24[27],stage2_23[61],stage2_22[65],stage2_21[77],stage2_20[106]}
   );
   gpc606_5 gpc2638 (
      {stage1_21[204], stage1_21[205], stage1_21[206], stage1_21[207], stage1_21[208], stage1_21[209]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[28],stage2_23[62],stage2_22[66],stage2_21[78]}
   );
   gpc606_5 gpc2639 (
      {stage1_21[210], stage1_21[211], stage1_21[212], stage1_21[213], stage1_21[214], stage1_21[215]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[29],stage2_23[63],stage2_22[67],stage2_21[79]}
   );
   gpc606_5 gpc2640 (
      {stage1_21[216], stage1_21[217], stage1_21[218], stage1_21[219], stage1_21[220], stage1_21[221]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[30],stage2_23[64],stage2_22[68],stage2_21[80]}
   );
   gpc615_5 gpc2641 (
      {stage1_21[222], stage1_21[223], stage1_21[224], stage1_21[225], stage1_21[226]},
      {stage1_22[168]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[31],stage2_23[65],stage2_22[69],stage2_21[81]}
   );
   gpc606_5 gpc2642 (
      {stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172], stage1_22[173], stage1_22[174]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[32],stage2_23[66],stage2_22[70]}
   );
   gpc606_5 gpc2643 (
      {stage1_22[175], stage1_22[176], stage1_22[177], stage1_22[178], stage1_22[179], stage1_22[180]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[33],stage2_23[67],stage2_22[71]}
   );
   gpc606_5 gpc2644 (
      {stage1_22[181], stage1_22[182], stage1_22[183], stage1_22[184], stage1_22[185], stage1_22[186]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[34],stage2_23[68],stage2_22[72]}
   );
   gpc606_5 gpc2645 (
      {stage1_22[187], stage1_22[188], stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[35],stage2_23[69],stage2_22[73]}
   );
   gpc615_5 gpc2646 (
      {stage1_22[193], stage1_22[194], stage1_22[195], stage1_22[196], stage1_22[197]},
      {stage1_23[24]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[36],stage2_23[70],stage2_22[74]}
   );
   gpc615_5 gpc2647 (
      {stage1_22[198], stage1_22[199], stage1_22[200], stage1_22[201], stage1_22[202]},
      {stage1_23[25]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[9],stage2_24[37],stage2_23[71],stage2_22[75]}
   );
   gpc615_5 gpc2648 (
      {stage1_22[203], stage1_22[204], stage1_22[205], stage1_22[206], stage1_22[207]},
      {stage1_23[26]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[10],stage2_24[38],stage2_23[72],stage2_22[76]}
   );
   gpc615_5 gpc2649 (
      {stage1_22[208], stage1_22[209], stage1_22[210], stage1_22[211], stage1_22[212]},
      {stage1_23[27]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[11],stage2_24[39],stage2_23[73],stage2_22[77]}
   );
   gpc615_5 gpc2650 (
      {stage1_22[213], stage1_22[214], stage1_22[215], stage1_22[216], stage1_22[217]},
      {stage1_23[28]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[12],stage2_24[40],stage2_23[74],stage2_22[78]}
   );
   gpc615_5 gpc2651 (
      {stage1_22[218], stage1_22[219], stage1_22[220], stage1_22[221], stage1_22[222]},
      {stage1_23[29]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[13],stage2_24[41],stage2_23[75],stage2_22[79]}
   );
   gpc615_5 gpc2652 (
      {stage1_22[223], stage1_22[224], stage1_22[225], stage1_22[226], stage1_22[227]},
      {stage1_23[30]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[14],stage2_24[42],stage2_23[76],stage2_22[80]}
   );
   gpc615_5 gpc2653 (
      {stage1_22[228], stage1_22[229], stage1_22[230], stage1_22[231], stage1_22[232]},
      {stage1_23[31]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[15],stage2_24[43],stage2_23[77],stage2_22[81]}
   );
   gpc615_5 gpc2654 (
      {stage1_22[233], stage1_22[234], stage1_22[235], stage1_22[236], stage1_22[237]},
      {stage1_23[32]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[16],stage2_24[44],stage2_23[78],stage2_22[82]}
   );
   gpc615_5 gpc2655 (
      {stage1_22[238], stage1_22[239], stage1_22[240], stage1_22[241], stage1_22[242]},
      {stage1_23[33]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[17],stage2_24[45],stage2_23[79],stage2_22[83]}
   );
   gpc615_5 gpc2656 (
      {stage1_22[243], stage1_22[244], stage1_22[245], stage1_22[246], stage1_22[247]},
      {stage1_23[34]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[18],stage2_24[46],stage2_23[80],stage2_22[84]}
   );
   gpc615_5 gpc2657 (
      {stage1_22[248], stage1_22[249], stage1_22[250], stage1_22[251], stage1_22[252]},
      {stage1_23[35]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[19],stage2_24[47],stage2_23[81],stage2_22[85]}
   );
   gpc615_5 gpc2658 (
      {stage1_22[253], stage1_22[254], stage1_22[255], stage1_22[256], stage1_22[257]},
      {stage1_23[36]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[20],stage2_24[48],stage2_23[82],stage2_22[86]}
   );
   gpc615_5 gpc2659 (
      {stage1_22[258], stage1_22[259], stage1_22[260], stage1_22[261], stage1_22[262]},
      {stage1_23[37]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[21],stage2_24[49],stage2_23[83],stage2_22[87]}
   );
   gpc615_5 gpc2660 (
      {stage1_22[263], stage1_22[264], stage1_22[265], stage1_22[266], stage1_22[267]},
      {stage1_23[38]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[22],stage2_24[50],stage2_23[84],stage2_22[88]}
   );
   gpc606_5 gpc2661 (
      {stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42], stage1_23[43], stage1_23[44]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[19],stage2_25[23],stage2_24[51],stage2_23[85]}
   );
   gpc606_5 gpc2662 (
      {stage1_23[45], stage1_23[46], stage1_23[47], stage1_23[48], stage1_23[49], stage1_23[50]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[20],stage2_25[24],stage2_24[52],stage2_23[86]}
   );
   gpc606_5 gpc2663 (
      {stage1_23[51], stage1_23[52], stage1_23[53], stage1_23[54], stage1_23[55], stage1_23[56]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[21],stage2_25[25],stage2_24[53],stage2_23[87]}
   );
   gpc606_5 gpc2664 (
      {stage1_23[57], stage1_23[58], stage1_23[59], stage1_23[60], stage1_23[61], stage1_23[62]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[22],stage2_25[26],stage2_24[54],stage2_23[88]}
   );
   gpc606_5 gpc2665 (
      {stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66], stage1_23[67], stage1_23[68]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[23],stage2_25[27],stage2_24[55],stage2_23[89]}
   );
   gpc606_5 gpc2666 (
      {stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72], stage1_23[73], stage1_23[74]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[24],stage2_25[28],stage2_24[56],stage2_23[90]}
   );
   gpc606_5 gpc2667 (
      {stage1_23[75], stage1_23[76], stage1_23[77], stage1_23[78], stage1_23[79], stage1_23[80]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[25],stage2_25[29],stage2_24[57],stage2_23[91]}
   );
   gpc606_5 gpc2668 (
      {stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84], stage1_23[85], stage1_23[86]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[26],stage2_25[30],stage2_24[58],stage2_23[92]}
   );
   gpc606_5 gpc2669 (
      {stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90], stage1_23[91], stage1_23[92]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[27],stage2_25[31],stage2_24[59],stage2_23[93]}
   );
   gpc606_5 gpc2670 (
      {stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96], stage1_23[97], stage1_23[98]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[28],stage2_25[32],stage2_24[60],stage2_23[94]}
   );
   gpc606_5 gpc2671 (
      {stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102], stage1_23[103], stage1_23[104]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[29],stage2_25[33],stage2_24[61],stage2_23[95]}
   );
   gpc606_5 gpc2672 (
      {stage1_23[105], stage1_23[106], stage1_23[107], stage1_23[108], stage1_23[109], stage1_23[110]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[30],stage2_25[34],stage2_24[62],stage2_23[96]}
   );
   gpc606_5 gpc2673 (
      {stage1_23[111], stage1_23[112], stage1_23[113], stage1_23[114], stage1_23[115], stage1_23[116]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[31],stage2_25[35],stage2_24[63],stage2_23[97]}
   );
   gpc606_5 gpc2674 (
      {stage1_23[117], stage1_23[118], stage1_23[119], stage1_23[120], stage1_23[121], stage1_23[122]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[32],stage2_25[36],stage2_24[64],stage2_23[98]}
   );
   gpc606_5 gpc2675 (
      {stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126], stage1_23[127], stage1_23[128]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[33],stage2_25[37],stage2_24[65],stage2_23[99]}
   );
   gpc606_5 gpc2676 (
      {stage1_23[129], stage1_23[130], stage1_23[131], stage1_23[132], stage1_23[133], stage1_23[134]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[34],stage2_25[38],stage2_24[66],stage2_23[100]}
   );
   gpc606_5 gpc2677 (
      {stage1_23[135], stage1_23[136], stage1_23[137], stage1_23[138], stage1_23[139], stage1_23[140]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[35],stage2_25[39],stage2_24[67],stage2_23[101]}
   );
   gpc615_5 gpc2678 (
      {stage1_23[141], stage1_23[142], stage1_23[143], stage1_23[144], stage1_23[145]},
      {stage1_24[114]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[36],stage2_25[40],stage2_24[68],stage2_23[102]}
   );
   gpc606_5 gpc2679 (
      {stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119], stage1_24[120]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[18],stage2_26[37],stage2_25[41],stage2_24[69]}
   );
   gpc606_5 gpc2680 (
      {stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125], stage1_24[126]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[19],stage2_26[38],stage2_25[42],stage2_24[70]}
   );
   gpc606_5 gpc2681 (
      {stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131], stage1_24[132]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[20],stage2_26[39],stage2_25[43],stage2_24[71]}
   );
   gpc606_5 gpc2682 (
      {stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137], stage1_24[138]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[21],stage2_26[40],stage2_25[44],stage2_24[72]}
   );
   gpc606_5 gpc2683 (
      {stage1_24[139], stage1_24[140], stage1_24[141], stage1_24[142], stage1_24[143], stage1_24[144]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[22],stage2_26[41],stage2_25[45],stage2_24[73]}
   );
   gpc606_5 gpc2684 (
      {stage1_24[145], stage1_24[146], stage1_24[147], stage1_24[148], stage1_24[149], stage1_24[150]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[23],stage2_26[42],stage2_25[46],stage2_24[74]}
   );
   gpc606_5 gpc2685 (
      {stage1_24[151], stage1_24[152], stage1_24[153], stage1_24[154], stage1_24[155], stage1_24[156]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[24],stage2_26[43],stage2_25[47],stage2_24[75]}
   );
   gpc606_5 gpc2686 (
      {stage1_24[157], stage1_24[158], stage1_24[159], stage1_24[160], stage1_24[161], stage1_24[162]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[25],stage2_26[44],stage2_25[48],stage2_24[76]}
   );
   gpc606_5 gpc2687 (
      {stage1_24[163], stage1_24[164], stage1_24[165], stage1_24[166], stage1_24[167], stage1_24[168]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[26],stage2_26[45],stage2_25[49],stage2_24[77]}
   );
   gpc606_5 gpc2688 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173], stage1_24[174]},
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage2_28[9],stage2_27[27],stage2_26[46],stage2_25[50],stage2_24[78]}
   );
   gpc606_5 gpc2689 (
      {stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178], stage1_24[179], stage1_24[180]},
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64], stage1_26[65]},
      {stage2_28[10],stage2_27[28],stage2_26[47],stage2_25[51],stage2_24[79]}
   );
   gpc606_5 gpc2690 (
      {stage1_24[181], stage1_24[182], stage1_24[183], stage1_24[184], stage1_24[185], stage1_24[186]},
      {stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69], stage1_26[70], stage1_26[71]},
      {stage2_28[11],stage2_27[29],stage2_26[48],stage2_25[52],stage2_24[80]}
   );
   gpc606_5 gpc2691 (
      {stage1_24[187], stage1_24[188], stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192]},
      {stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77]},
      {stage2_28[12],stage2_27[30],stage2_26[49],stage2_25[53],stage2_24[81]}
   );
   gpc606_5 gpc2692 (
      {stage1_24[193], stage1_24[194], stage1_24[195], stage1_24[196], stage1_24[197], stage1_24[198]},
      {stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83]},
      {stage2_28[13],stage2_27[31],stage2_26[50],stage2_25[54],stage2_24[82]}
   );
   gpc606_5 gpc2693 (
      {stage1_24[199], stage1_24[200], stage1_24[201], stage1_24[202], stage1_24[203], stage1_24[204]},
      {stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage2_28[14],stage2_27[32],stage2_26[51],stage2_25[55],stage2_24[83]}
   );
   gpc606_5 gpc2694 (
      {stage1_24[205], stage1_24[206], stage1_24[207], stage1_24[208], stage1_24[209], stage1_24[210]},
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94], stage1_26[95]},
      {stage2_28[15],stage2_27[33],stage2_26[52],stage2_25[56],stage2_24[84]}
   );
   gpc606_5 gpc2695 (
      {stage1_24[211], stage1_24[212], stage1_24[213], stage1_24[214], stage1_24[215], stage1_24[216]},
      {stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99], stage1_26[100], stage1_26[101]},
      {stage2_28[16],stage2_27[34],stage2_26[53],stage2_25[57],stage2_24[85]}
   );
   gpc606_5 gpc2696 (
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[17],stage2_27[35],stage2_26[54],stage2_25[58]}
   );
   gpc606_5 gpc2697 (
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[18],stage2_27[36],stage2_26[55],stage2_25[59]}
   );
   gpc606_5 gpc2698 (
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[19],stage2_27[37],stage2_26[56],stage2_25[60]}
   );
   gpc606_5 gpc2699 (
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[20],stage2_27[38],stage2_26[57],stage2_25[61]}
   );
   gpc606_5 gpc2700 (
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[21],stage2_27[39],stage2_26[58],stage2_25[62]}
   );
   gpc606_5 gpc2701 (
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[22],stage2_27[40],stage2_26[59],stage2_25[63]}
   );
   gpc606_5 gpc2702 (
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[23],stage2_27[41],stage2_26[60],stage2_25[64]}
   );
   gpc606_5 gpc2703 (
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage1_27[42], stage1_27[43], stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47]},
      {stage2_29[7],stage2_28[24],stage2_27[42],stage2_26[61],stage2_25[65]}
   );
   gpc606_5 gpc2704 (
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53]},
      {stage2_29[8],stage2_28[25],stage2_27[43],stage2_26[62],stage2_25[66]}
   );
   gpc606_5 gpc2705 (
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage2_29[9],stage2_28[26],stage2_27[44],stage2_26[63],stage2_25[67]}
   );
   gpc606_5 gpc2706 (
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage1_27[60], stage1_27[61], stage1_27[62], stage1_27[63], stage1_27[64], stage1_27[65]},
      {stage2_29[10],stage2_28[27],stage2_27[45],stage2_26[64],stage2_25[68]}
   );
   gpc606_5 gpc2707 (
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage1_27[66], stage1_27[67], stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71]},
      {stage2_29[11],stage2_28[28],stage2_27[46],stage2_26[65],stage2_25[69]}
   );
   gpc606_5 gpc2708 (
      {stage1_25[180], stage1_25[181], stage1_25[182], stage1_25[183], stage1_25[184], stage1_25[185]},
      {stage1_27[72], stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage2_29[12],stage2_28[29],stage2_27[47],stage2_26[66],stage2_25[70]}
   );
   gpc606_5 gpc2709 (
      {stage1_25[186], stage1_25[187], stage1_25[188], stage1_25[189], stage1_25[190], stage1_25[191]},
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82], stage1_27[83]},
      {stage2_29[13],stage2_28[30],stage2_27[48],stage2_26[67],stage2_25[71]}
   );
   gpc606_5 gpc2710 (
      {stage1_25[192], stage1_25[193], stage1_25[194], stage1_25[195], stage1_25[196], stage1_25[197]},
      {stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87], stage1_27[88], stage1_27[89]},
      {stage2_29[14],stage2_28[31],stage2_27[49],stage2_26[68],stage2_25[72]}
   );
   gpc606_5 gpc2711 (
      {stage1_25[198], stage1_25[199], stage1_25[200], stage1_25[201], stage1_25[202], stage1_25[203]},
      {stage1_27[90], stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94], stage1_27[95]},
      {stage2_29[15],stage2_28[32],stage2_27[50],stage2_26[69],stage2_25[73]}
   );
   gpc606_5 gpc2712 (
      {stage1_25[204], stage1_25[205], stage1_25[206], stage1_25[207], stage1_25[208], stage1_25[209]},
      {stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99], stage1_27[100], stage1_27[101]},
      {stage2_29[16],stage2_28[33],stage2_27[51],stage2_26[70],stage2_25[74]}
   );
   gpc615_5 gpc2713 (
      {stage1_25[210], stage1_25[211], stage1_25[212], stage1_25[213], stage1_25[214]},
      {stage1_26[102]},
      {stage1_27[102], stage1_27[103], stage1_27[104], stage1_27[105], stage1_27[106], stage1_27[107]},
      {stage2_29[17],stage2_28[34],stage2_27[52],stage2_26[71],stage2_25[75]}
   );
   gpc615_5 gpc2714 (
      {stage1_25[215], stage1_25[216], stage1_25[217], stage1_25[218], stage1_25[219]},
      {stage1_26[103]},
      {stage1_27[108], stage1_27[109], stage1_27[110], stage1_27[111], stage1_27[112], stage1_27[113]},
      {stage2_29[18],stage2_28[35],stage2_27[53],stage2_26[72],stage2_25[76]}
   );
   gpc615_5 gpc2715 (
      {stage1_25[220], stage1_25[221], stage1_25[222], stage1_25[223], stage1_25[224]},
      {stage1_26[104]},
      {stage1_27[114], stage1_27[115], stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119]},
      {stage2_29[19],stage2_28[36],stage2_27[54],stage2_26[73],stage2_25[77]}
   );
   gpc615_5 gpc2716 (
      {stage1_25[225], stage1_25[226], stage1_25[227], stage1_25[228], stage1_25[229]},
      {stage1_26[105]},
      {stage1_27[120], stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124], stage1_27[125]},
      {stage2_29[20],stage2_28[37],stage2_27[55],stage2_26[74],stage2_25[78]}
   );
   gpc615_5 gpc2717 (
      {stage1_25[230], stage1_25[231], stage1_25[232], stage1_25[233], stage1_25[234]},
      {stage1_26[106]},
      {stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129], stage1_27[130], stage1_27[131]},
      {stage2_29[21],stage2_28[38],stage2_27[56],stage2_26[75],stage2_25[79]}
   );
   gpc615_5 gpc2718 (
      {stage1_25[235], stage1_25[236], stage1_25[237], stage1_25[238], stage1_25[239]},
      {stage1_26[107]},
      {stage1_27[132], stage1_27[133], stage1_27[134], stage1_27[135], stage1_27[136], stage1_27[137]},
      {stage2_29[22],stage2_28[39],stage2_27[57],stage2_26[76],stage2_25[80]}
   );
   gpc615_5 gpc2719 (
      {stage1_25[240], stage1_25[241], stage1_25[242], stage1_25[243], stage1_25[244]},
      {stage1_26[108]},
      {stage1_27[138], stage1_27[139], stage1_27[140], stage1_27[141], stage1_27[142], stage1_27[143]},
      {stage2_29[23],stage2_28[40],stage2_27[58],stage2_26[77],stage2_25[81]}
   );
   gpc615_5 gpc2720 (
      {stage1_25[245], stage1_25[246], stage1_25[247], stage1_25[248], stage1_25[249]},
      {stage1_26[109]},
      {stage1_27[144], stage1_27[145], stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149]},
      {stage2_29[24],stage2_28[41],stage2_27[59],stage2_26[78],stage2_25[82]}
   );
   gpc615_5 gpc2721 (
      {stage1_25[250], stage1_25[251], stage1_25[252], stage1_25[253], stage1_25[254]},
      {stage1_26[110]},
      {stage1_27[150], stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154], stage1_27[155]},
      {stage2_29[25],stage2_28[42],stage2_27[60],stage2_26[79],stage2_25[83]}
   );
   gpc615_5 gpc2722 (
      {stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114], stage1_26[115]},
      {stage1_27[156]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[26],stage2_28[43],stage2_27[61],stage2_26[80]}
   );
   gpc615_5 gpc2723 (
      {stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119], stage1_26[120]},
      {stage1_27[157]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[27],stage2_28[44],stage2_27[62],stage2_26[81]}
   );
   gpc615_5 gpc2724 (
      {stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124], stage1_26[125]},
      {stage1_27[158]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[28],stage2_28[45],stage2_27[63],stage2_26[82]}
   );
   gpc615_5 gpc2725 (
      {stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129], stage1_26[130]},
      {stage1_27[159]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[29],stage2_28[46],stage2_27[64],stage2_26[83]}
   );
   gpc615_5 gpc2726 (
      {stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134], stage1_26[135]},
      {stage1_27[160]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[30],stage2_28[47],stage2_27[65],stage2_26[84]}
   );
   gpc615_5 gpc2727 (
      {stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139], stage1_26[140]},
      {stage1_27[161]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[31],stage2_28[48],stage2_27[66],stage2_26[85]}
   );
   gpc615_5 gpc2728 (
      {stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144], stage1_26[145]},
      {stage1_27[162]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[32],stage2_28[49],stage2_27[67],stage2_26[86]}
   );
   gpc615_5 gpc2729 (
      {stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149], stage1_26[150]},
      {stage1_27[163]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[33],stage2_28[50],stage2_27[68],stage2_26[87]}
   );
   gpc615_5 gpc2730 (
      {stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154], stage1_26[155]},
      {stage1_27[164]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[34],stage2_28[51],stage2_27[69],stage2_26[88]}
   );
   gpc615_5 gpc2731 (
      {stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159], stage1_26[160]},
      {stage1_27[165]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[35],stage2_28[52],stage2_27[70],stage2_26[89]}
   );
   gpc615_5 gpc2732 (
      {stage1_26[161], stage1_26[162], stage1_26[163], stage1_26[164], stage1_26[165]},
      {stage1_27[166]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[36],stage2_28[53],stage2_27[71],stage2_26[90]}
   );
   gpc615_5 gpc2733 (
      {stage1_26[166], stage1_26[167], stage1_26[168], stage1_26[169], stage1_26[170]},
      {stage1_27[167]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[37],stage2_28[54],stage2_27[72],stage2_26[91]}
   );
   gpc615_5 gpc2734 (
      {stage1_26[171], stage1_26[172], stage1_26[173], stage1_26[174], stage1_26[175]},
      {stage1_27[168]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[38],stage2_28[55],stage2_27[73],stage2_26[92]}
   );
   gpc615_5 gpc2735 (
      {stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179], stage1_26[180]},
      {stage1_27[169]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[39],stage2_28[56],stage2_27[74],stage2_26[93]}
   );
   gpc615_5 gpc2736 (
      {stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184], stage1_26[185]},
      {stage1_27[170]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[40],stage2_28[57],stage2_27[75],stage2_26[94]}
   );
   gpc615_5 gpc2737 (
      {stage1_27[171], stage1_27[172], stage1_27[173], stage1_27[174], stage1_27[175]},
      {stage1_28[90]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[15],stage2_29[41],stage2_28[58],stage2_27[76]}
   );
   gpc615_5 gpc2738 (
      {stage1_27[176], stage1_27[177], stage1_27[178], stage1_27[179], stage1_27[180]},
      {stage1_28[91]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[16],stage2_29[42],stage2_28[59],stage2_27[77]}
   );
   gpc615_5 gpc2739 (
      {stage1_27[181], stage1_27[182], stage1_27[183], stage1_27[184], stage1_27[185]},
      {stage1_28[92]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[17],stage2_29[43],stage2_28[60],stage2_27[78]}
   );
   gpc615_5 gpc2740 (
      {stage1_27[186], stage1_27[187], stage1_27[188], stage1_27[189], stage1_27[190]},
      {stage1_28[93]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[18],stage2_29[44],stage2_28[61],stage2_27[79]}
   );
   gpc615_5 gpc2741 (
      {stage1_27[191], stage1_27[192], stage1_27[193], stage1_27[194], stage1_27[195]},
      {stage1_28[94]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[19],stage2_29[45],stage2_28[62],stage2_27[80]}
   );
   gpc606_5 gpc2742 (
      {stage1_28[95], stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[5],stage2_30[20],stage2_29[46],stage2_28[63]}
   );
   gpc606_5 gpc2743 (
      {stage1_28[101], stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[6],stage2_30[21],stage2_29[47],stage2_28[64]}
   );
   gpc606_5 gpc2744 (
      {stage1_28[107], stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[7],stage2_30[22],stage2_29[48],stage2_28[65]}
   );
   gpc606_5 gpc2745 (
      {stage1_28[113], stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[8],stage2_30[23],stage2_29[49],stage2_28[66]}
   );
   gpc606_5 gpc2746 (
      {stage1_28[119], stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[9],stage2_30[24],stage2_29[50],stage2_28[67]}
   );
   gpc606_5 gpc2747 (
      {stage1_28[125], stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[10],stage2_30[25],stage2_29[51],stage2_28[68]}
   );
   gpc606_5 gpc2748 (
      {stage1_28[131], stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[11],stage2_30[26],stage2_29[52],stage2_28[69]}
   );
   gpc606_5 gpc2749 (
      {stage1_28[137], stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[12],stage2_30[27],stage2_29[53],stage2_28[70]}
   );
   gpc606_5 gpc2750 (
      {stage1_28[143], stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[13],stage2_30[28],stage2_29[54],stage2_28[71]}
   );
   gpc606_5 gpc2751 (
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[9],stage2_31[14],stage2_30[29],stage2_29[55]}
   );
   gpc606_5 gpc2752 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[10],stage2_31[15],stage2_30[30],stage2_29[56]}
   );
   gpc606_5 gpc2753 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[11],stage2_31[16],stage2_30[31],stage2_29[57]}
   );
   gpc606_5 gpc2754 (
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[12],stage2_31[17],stage2_30[32],stage2_29[58]}
   );
   gpc606_5 gpc2755 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[13],stage2_31[18],stage2_30[33],stage2_29[59]}
   );
   gpc606_5 gpc2756 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[14],stage2_31[19],stage2_30[34],stage2_29[60]}
   );
   gpc606_5 gpc2757 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[15],stage2_31[20],stage2_30[35],stage2_29[61]}
   );
   gpc606_5 gpc2758 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[16],stage2_31[21],stage2_30[36],stage2_29[62]}
   );
   gpc606_5 gpc2759 (
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[17],stage2_31[22],stage2_30[37],stage2_29[63]}
   );
   gpc606_5 gpc2760 (
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[18],stage2_31[23],stage2_30[38],stage2_29[64]}
   );
   gpc606_5 gpc2761 (
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage2_33[10],stage2_32[19],stage2_31[24],stage2_30[39],stage2_29[65]}
   );
   gpc606_5 gpc2762 (
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage2_33[11],stage2_32[20],stage2_31[25],stage2_30[40],stage2_29[66]}
   );
   gpc606_5 gpc2763 (
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage2_33[12],stage2_32[21],stage2_31[26],stage2_30[41],stage2_29[67]}
   );
   gpc606_5 gpc2764 (
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage2_33[13],stage2_32[22],stage2_31[27],stage2_30[42],stage2_29[68]}
   );
   gpc606_5 gpc2765 (
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage2_33[14],stage2_32[23],stage2_31[28],stage2_30[43],stage2_29[69]}
   );
   gpc606_5 gpc2766 (
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94], stage1_31[95]},
      {stage2_33[15],stage2_32[24],stage2_31[29],stage2_30[44],stage2_29[70]}
   );
   gpc606_5 gpc2767 (
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100], stage1_31[101]},
      {stage2_33[16],stage2_32[25],stage2_31[30],stage2_30[45],stage2_29[71]}
   );
   gpc606_5 gpc2768 (
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106], stage1_31[107]},
      {stage2_33[17],stage2_32[26],stage2_31[31],stage2_30[46],stage2_29[72]}
   );
   gpc606_5 gpc2769 (
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113]},
      {stage2_33[18],stage2_32[27],stage2_31[32],stage2_30[47],stage2_29[73]}
   );
   gpc606_5 gpc2770 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage2_33[19],stage2_32[28],stage2_31[33],stage2_30[48],stage2_29[74]}
   );
   gpc606_5 gpc2771 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124], stage1_31[125]},
      {stage2_33[20],stage2_32[29],stage2_31[34],stage2_30[49],stage2_29[75]}
   );
   gpc606_5 gpc2772 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129], stage1_31[130], stage1_31[131]},
      {stage2_33[21],stage2_32[30],stage2_31[35],stage2_30[50],stage2_29[76]}
   );
   gpc606_5 gpc2773 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[132], stage1_31[133], stage1_31[134], stage1_31[135], stage1_31[136], stage1_31[137]},
      {stage2_33[22],stage2_32[31],stage2_31[36],stage2_30[51],stage2_29[77]}
   );
   gpc606_5 gpc2774 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[138], stage1_31[139], stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143]},
      {stage2_33[23],stage2_32[32],stage2_31[37],stage2_30[52],stage2_29[78]}
   );
   gpc606_5 gpc2775 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[144], stage1_31[145], stage1_31[146], stage1_31[147], stage1_31[148], stage1_31[149]},
      {stage2_33[24],stage2_32[33],stage2_31[38],stage2_30[53],stage2_29[79]}
   );
   gpc606_5 gpc2776 (
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[25],stage2_32[34],stage2_31[39],stage2_30[54]}
   );
   gpc606_5 gpc2777 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[26],stage2_32[35],stage2_31[40],stage2_30[55]}
   );
   gpc606_5 gpc2778 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[27],stage2_32[36],stage2_31[41],stage2_30[56]}
   );
   gpc606_5 gpc2779 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[28],stage2_32[37],stage2_31[42],stage2_30[57]}
   );
   gpc606_5 gpc2780 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[29],stage2_32[38],stage2_31[43],stage2_30[58]}
   );
   gpc606_5 gpc2781 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[30],stage2_32[39],stage2_31[44],stage2_30[59]}
   );
   gpc606_5 gpc2782 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[31],stage2_32[40],stage2_31[45],stage2_30[60]}
   );
   gpc606_5 gpc2783 (
      {stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99], stage1_30[100], stage1_30[101]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[32],stage2_32[41],stage2_31[46],stage2_30[61]}
   );
   gpc606_5 gpc2784 (
      {stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105], stage1_30[106], stage1_30[107]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[33],stage2_32[42],stage2_31[47],stage2_30[62]}
   );
   gpc606_5 gpc2785 (
      {stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[34],stage2_32[43],stage2_31[48],stage2_30[63]}
   );
   gpc606_5 gpc2786 (
      {stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[35],stage2_32[44],stage2_31[49],stage2_30[64]}
   );
   gpc606_5 gpc2787 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124], stage1_30[125]},
      {stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70], stage1_32[71]},
      {stage2_34[11],stage2_33[36],stage2_32[45],stage2_31[50],stage2_30[65]}
   );
   gpc606_5 gpc2788 (
      {stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129], stage1_30[130], stage1_30[131]},
      {stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76], stage1_32[77]},
      {stage2_34[12],stage2_33[37],stage2_32[46],stage2_31[51],stage2_30[66]}
   );
   gpc606_5 gpc2789 (
      {stage1_30[132], stage1_30[133], stage1_30[134], stage1_30[135], stage1_30[136], stage1_30[137]},
      {stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82], stage1_32[83]},
      {stage2_34[13],stage2_33[38],stage2_32[47],stage2_31[52],stage2_30[67]}
   );
   gpc606_5 gpc2790 (
      {stage1_30[138], stage1_30[139], stage1_30[140], stage1_30[141], stage1_30[142], stage1_30[143]},
      {stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88], stage1_32[89]},
      {stage2_34[14],stage2_33[39],stage2_32[48],stage2_31[53],stage2_30[68]}
   );
   gpc606_5 gpc2791 (
      {stage1_30[144], stage1_30[145], stage1_30[146], stage1_30[147], stage1_30[148], stage1_30[149]},
      {stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94], stage1_32[95]},
      {stage2_34[15],stage2_33[40],stage2_32[49],stage2_31[54],stage2_30[69]}
   );
   gpc606_5 gpc2792 (
      {stage1_30[150], stage1_30[151], stage1_30[152], stage1_30[153], stage1_30[154], stage1_30[155]},
      {stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100], stage1_32[101]},
      {stage2_34[16],stage2_33[41],stage2_32[50],stage2_31[55],stage2_30[70]}
   );
   gpc606_5 gpc2793 (
      {stage1_30[156], stage1_30[157], stage1_30[158], stage1_30[159], stage1_30[160], stage1_30[161]},
      {stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106], stage1_32[107]},
      {stage2_34[17],stage2_33[42],stage2_32[51],stage2_31[56],stage2_30[71]}
   );
   gpc606_5 gpc2794 (
      {stage1_30[162], stage1_30[163], stage1_30[164], stage1_30[165], stage1_30[166], stage1_30[167]},
      {stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112], stage1_32[113]},
      {stage2_34[18],stage2_33[43],stage2_32[52],stage2_31[57],stage2_30[72]}
   );
   gpc606_5 gpc2795 (
      {stage1_30[168], stage1_30[169], stage1_30[170], stage1_30[171], stage1_30[172], stage1_30[173]},
      {stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118], stage1_32[119]},
      {stage2_34[19],stage2_33[44],stage2_32[53],stage2_31[58],stage2_30[73]}
   );
   gpc606_5 gpc2796 (
      {stage1_30[174], stage1_30[175], stage1_30[176], stage1_30[177], stage1_30[178], stage1_30[179]},
      {stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124], stage1_32[125]},
      {stage2_34[20],stage2_33[45],stage2_32[54],stage2_31[59],stage2_30[74]}
   );
   gpc606_5 gpc2797 (
      {stage1_30[180], stage1_30[181], stage1_30[182], stage1_30[183], stage1_30[184], stage1_30[185]},
      {stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130], stage1_32[131]},
      {stage2_34[21],stage2_33[46],stage2_32[55],stage2_31[60],stage2_30[75]}
   );
   gpc606_5 gpc2798 (
      {stage1_30[186], stage1_30[187], stage1_30[188], stage1_30[189], stage1_30[190], stage1_30[191]},
      {stage1_32[132], stage1_32[133], stage1_32[134], stage1_32[135], stage1_32[136], stage1_32[137]},
      {stage2_34[22],stage2_33[47],stage2_32[56],stage2_31[61],stage2_30[76]}
   );
   gpc606_5 gpc2799 (
      {stage1_31[150], stage1_31[151], stage1_31[152], stage1_31[153], stage1_31[154], stage1_31[155]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[23],stage2_33[48],stage2_32[57],stage2_31[62]}
   );
   gpc606_5 gpc2800 (
      {stage1_31[156], stage1_31[157], stage1_31[158], stage1_31[159], stage1_31[160], stage1_31[161]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[24],stage2_33[49],stage2_32[58],stage2_31[63]}
   );
   gpc606_5 gpc2801 (
      {stage1_31[162], stage1_31[163], stage1_31[164], stage1_31[165], stage1_31[166], stage1_31[167]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[25],stage2_33[50],stage2_32[59],stage2_31[64]}
   );
   gpc606_5 gpc2802 (
      {stage1_31[168], stage1_31[169], stage1_31[170], stage1_31[171], stage1_31[172], stage1_31[173]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[26],stage2_33[51],stage2_32[60],stage2_31[65]}
   );
   gpc606_5 gpc2803 (
      {stage1_31[174], stage1_31[175], stage1_31[176], stage1_31[177], stage1_31[178], stage1_31[179]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[27],stage2_33[52],stage2_32[61],stage2_31[66]}
   );
   gpc615_5 gpc2804 (
      {stage1_31[180], stage1_31[181], stage1_31[182], stage1_31[183], stage1_31[184]},
      {stage1_32[138]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[28],stage2_33[53],stage2_32[62],stage2_31[67]}
   );
   gpc615_5 gpc2805 (
      {stage1_31[185], stage1_31[186], stage1_31[187], stage1_31[188], stage1_31[189]},
      {stage1_32[139]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[29],stage2_33[54],stage2_32[63],stage2_31[68]}
   );
   gpc615_5 gpc2806 (
      {stage1_31[190], stage1_31[191], stage1_31[192], stage1_31[193], stage1_31[194]},
      {stage1_32[140]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[30],stage2_33[55],stage2_32[64],stage2_31[69]}
   );
   gpc615_5 gpc2807 (
      {stage1_31[195], stage1_31[196], stage1_31[197], stage1_31[198], stage1_31[199]},
      {stage1_32[141]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[31],stage2_33[56],stage2_32[65],stage2_31[70]}
   );
   gpc615_5 gpc2808 (
      {stage1_31[200], stage1_31[201], stage1_31[202], stage1_31[203], stage1_31[204]},
      {stage1_32[142]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[32],stage2_33[57],stage2_32[66],stage2_31[71]}
   );
   gpc615_5 gpc2809 (
      {stage1_31[205], stage1_31[206], stage1_31[207], stage1_31[208], stage1_31[209]},
      {stage1_32[143]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[33],stage2_33[58],stage2_32[67],stage2_31[72]}
   );
   gpc615_5 gpc2810 (
      {stage1_31[210], stage1_31[211], stage1_31[212], stage1_31[213], stage1_31[214]},
      {stage1_32[144]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], 1'b0},
      {stage2_35[11],stage2_34[34],stage2_33[59],stage2_32[68],stage2_31[73]}
   );
   gpc1_1 gpc2811 (
      {stage1_0[60]},
      {stage2_0[12]}
   );
   gpc1_1 gpc2812 (
      {stage1_0[61]},
      {stage2_0[13]}
   );
   gpc1_1 gpc2813 (
      {stage1_0[62]},
      {stage2_0[14]}
   );
   gpc1_1 gpc2814 (
      {stage1_0[63]},
      {stage2_0[15]}
   );
   gpc1_1 gpc2815 (
      {stage1_0[64]},
      {stage2_0[16]}
   );
   gpc1_1 gpc2816 (
      {stage1_0[65]},
      {stage2_0[17]}
   );
   gpc1_1 gpc2817 (
      {stage1_0[66]},
      {stage2_0[18]}
   );
   gpc1_1 gpc2818 (
      {stage1_0[67]},
      {stage2_0[19]}
   );
   gpc1_1 gpc2819 (
      {stage1_0[68]},
      {stage2_0[20]}
   );
   gpc1_1 gpc2820 (
      {stage1_0[69]},
      {stage2_0[21]}
   );
   gpc1_1 gpc2821 (
      {stage1_0[70]},
      {stage2_0[22]}
   );
   gpc1_1 gpc2822 (
      {stage1_0[71]},
      {stage2_0[23]}
   );
   gpc1_1 gpc2823 (
      {stage1_0[72]},
      {stage2_0[24]}
   );
   gpc1_1 gpc2824 (
      {stage1_0[73]},
      {stage2_0[25]}
   );
   gpc1_1 gpc2825 (
      {stage1_0[74]},
      {stage2_0[26]}
   );
   gpc1_1 gpc2826 (
      {stage1_0[75]},
      {stage2_0[27]}
   );
   gpc1_1 gpc2827 (
      {stage1_0[76]},
      {stage2_0[28]}
   );
   gpc1_1 gpc2828 (
      {stage1_0[77]},
      {stage2_0[29]}
   );
   gpc1_1 gpc2829 (
      {stage1_0[78]},
      {stage2_0[30]}
   );
   gpc1_1 gpc2830 (
      {stage1_0[79]},
      {stage2_0[31]}
   );
   gpc1_1 gpc2831 (
      {stage1_0[80]},
      {stage2_0[32]}
   );
   gpc1_1 gpc2832 (
      {stage1_0[81]},
      {stage2_0[33]}
   );
   gpc1_1 gpc2833 (
      {stage1_0[82]},
      {stage2_0[34]}
   );
   gpc1_1 gpc2834 (
      {stage1_0[83]},
      {stage2_0[35]}
   );
   gpc1_1 gpc2835 (
      {stage1_0[84]},
      {stage2_0[36]}
   );
   gpc1_1 gpc2836 (
      {stage1_0[85]},
      {stage2_0[37]}
   );
   gpc1_1 gpc2837 (
      {stage1_0[86]},
      {stage2_0[38]}
   );
   gpc1_1 gpc2838 (
      {stage1_0[87]},
      {stage2_0[39]}
   );
   gpc1_1 gpc2839 (
      {stage1_0[88]},
      {stage2_0[40]}
   );
   gpc1_1 gpc2840 (
      {stage1_0[89]},
      {stage2_0[41]}
   );
   gpc1_1 gpc2841 (
      {stage1_0[90]},
      {stage2_0[42]}
   );
   gpc1_1 gpc2842 (
      {stage1_0[91]},
      {stage2_0[43]}
   );
   gpc1_1 gpc2843 (
      {stage1_0[92]},
      {stage2_0[44]}
   );
   gpc1_1 gpc2844 (
      {stage1_0[93]},
      {stage2_0[45]}
   );
   gpc1_1 gpc2845 (
      {stage1_0[94]},
      {stage2_0[46]}
   );
   gpc1_1 gpc2846 (
      {stage1_0[95]},
      {stage2_0[47]}
   );
   gpc1_1 gpc2847 (
      {stage1_0[96]},
      {stage2_0[48]}
   );
   gpc1_1 gpc2848 (
      {stage1_0[97]},
      {stage2_0[49]}
   );
   gpc1_1 gpc2849 (
      {stage1_0[98]},
      {stage2_0[50]}
   );
   gpc1_1 gpc2850 (
      {stage1_0[99]},
      {stage2_0[51]}
   );
   gpc1_1 gpc2851 (
      {stage1_0[100]},
      {stage2_0[52]}
   );
   gpc1_1 gpc2852 (
      {stage1_0[101]},
      {stage2_0[53]}
   );
   gpc1_1 gpc2853 (
      {stage1_0[102]},
      {stage2_0[54]}
   );
   gpc1_1 gpc2854 (
      {stage1_0[103]},
      {stage2_0[55]}
   );
   gpc1_1 gpc2855 (
      {stage1_0[104]},
      {stage2_0[56]}
   );
   gpc1_1 gpc2856 (
      {stage1_0[105]},
      {stage2_0[57]}
   );
   gpc1_1 gpc2857 (
      {stage1_0[106]},
      {stage2_0[58]}
   );
   gpc1_1 gpc2858 (
      {stage1_0[107]},
      {stage2_0[59]}
   );
   gpc1_1 gpc2859 (
      {stage1_0[108]},
      {stage2_0[60]}
   );
   gpc1_1 gpc2860 (
      {stage1_0[109]},
      {stage2_0[61]}
   );
   gpc1_1 gpc2861 (
      {stage1_0[110]},
      {stage2_0[62]}
   );
   gpc1_1 gpc2862 (
      {stage1_1[182]},
      {stage2_1[39]}
   );
   gpc1_1 gpc2863 (
      {stage1_1[183]},
      {stage2_1[40]}
   );
   gpc1_1 gpc2864 (
      {stage1_1[184]},
      {stage2_1[41]}
   );
   gpc1_1 gpc2865 (
      {stage1_1[185]},
      {stage2_1[42]}
   );
   gpc1_1 gpc2866 (
      {stage1_1[186]},
      {stage2_1[43]}
   );
   gpc1_1 gpc2867 (
      {stage1_1[187]},
      {stage2_1[44]}
   );
   gpc1_1 gpc2868 (
      {stage1_1[188]},
      {stage2_1[45]}
   );
   gpc1_1 gpc2869 (
      {stage1_1[189]},
      {stage2_1[46]}
   );
   gpc1_1 gpc2870 (
      {stage1_1[190]},
      {stage2_1[47]}
   );
   gpc1_1 gpc2871 (
      {stage1_1[191]},
      {stage2_1[48]}
   );
   gpc1_1 gpc2872 (
      {stage1_1[192]},
      {stage2_1[49]}
   );
   gpc1_1 gpc2873 (
      {stage1_1[193]},
      {stage2_1[50]}
   );
   gpc1_1 gpc2874 (
      {stage1_1[194]},
      {stage2_1[51]}
   );
   gpc1_1 gpc2875 (
      {stage1_1[195]},
      {stage2_1[52]}
   );
   gpc1_1 gpc2876 (
      {stage1_1[196]},
      {stage2_1[53]}
   );
   gpc1_1 gpc2877 (
      {stage1_1[197]},
      {stage2_1[54]}
   );
   gpc1_1 gpc2878 (
      {stage1_1[198]},
      {stage2_1[55]}
   );
   gpc1_1 gpc2879 (
      {stage1_2[152]},
      {stage2_2[59]}
   );
   gpc1_1 gpc2880 (
      {stage1_2[153]},
      {stage2_2[60]}
   );
   gpc1_1 gpc2881 (
      {stage1_2[154]},
      {stage2_2[61]}
   );
   gpc1_1 gpc2882 (
      {stage1_2[155]},
      {stage2_2[62]}
   );
   gpc1_1 gpc2883 (
      {stage1_2[156]},
      {stage2_2[63]}
   );
   gpc1_1 gpc2884 (
      {stage1_2[157]},
      {stage2_2[64]}
   );
   gpc1_1 gpc2885 (
      {stage1_2[158]},
      {stage2_2[65]}
   );
   gpc1_1 gpc2886 (
      {stage1_2[159]},
      {stage2_2[66]}
   );
   gpc1_1 gpc2887 (
      {stage1_2[160]},
      {stage2_2[67]}
   );
   gpc1_1 gpc2888 (
      {stage1_2[161]},
      {stage2_2[68]}
   );
   gpc1_1 gpc2889 (
      {stage1_2[162]},
      {stage2_2[69]}
   );
   gpc1_1 gpc2890 (
      {stage1_2[163]},
      {stage2_2[70]}
   );
   gpc1_1 gpc2891 (
      {stage1_2[164]},
      {stage2_2[71]}
   );
   gpc1_1 gpc2892 (
      {stage1_2[165]},
      {stage2_2[72]}
   );
   gpc1_1 gpc2893 (
      {stage1_2[166]},
      {stage2_2[73]}
   );
   gpc1_1 gpc2894 (
      {stage1_2[167]},
      {stage2_2[74]}
   );
   gpc1_1 gpc2895 (
      {stage1_2[168]},
      {stage2_2[75]}
   );
   gpc1_1 gpc2896 (
      {stage1_2[169]},
      {stage2_2[76]}
   );
   gpc1_1 gpc2897 (
      {stage1_2[170]},
      {stage2_2[77]}
   );
   gpc1_1 gpc2898 (
      {stage1_2[171]},
      {stage2_2[78]}
   );
   gpc1_1 gpc2899 (
      {stage1_2[172]},
      {stage2_2[79]}
   );
   gpc1_1 gpc2900 (
      {stage1_2[173]},
      {stage2_2[80]}
   );
   gpc1_1 gpc2901 (
      {stage1_2[174]},
      {stage2_2[81]}
   );
   gpc1_1 gpc2902 (
      {stage1_2[175]},
      {stage2_2[82]}
   );
   gpc1_1 gpc2903 (
      {stage1_2[176]},
      {stage2_2[83]}
   );
   gpc1_1 gpc2904 (
      {stage1_2[177]},
      {stage2_2[84]}
   );
   gpc1_1 gpc2905 (
      {stage1_2[178]},
      {stage2_2[85]}
   );
   gpc1_1 gpc2906 (
      {stage1_2[179]},
      {stage2_2[86]}
   );
   gpc1_1 gpc2907 (
      {stage1_2[180]},
      {stage2_2[87]}
   );
   gpc1_1 gpc2908 (
      {stage1_2[181]},
      {stage2_2[88]}
   );
   gpc1_1 gpc2909 (
      {stage1_2[182]},
      {stage2_2[89]}
   );
   gpc1_1 gpc2910 (
      {stage1_2[183]},
      {stage2_2[90]}
   );
   gpc1_1 gpc2911 (
      {stage1_2[184]},
      {stage2_2[91]}
   );
   gpc1_1 gpc2912 (
      {stage1_2[185]},
      {stage2_2[92]}
   );
   gpc1_1 gpc2913 (
      {stage1_2[186]},
      {stage2_2[93]}
   );
   gpc1_1 gpc2914 (
      {stage1_2[187]},
      {stage2_2[94]}
   );
   gpc1_1 gpc2915 (
      {stage1_4[217]},
      {stage2_4[91]}
   );
   gpc1_1 gpc2916 (
      {stage1_4[218]},
      {stage2_4[92]}
   );
   gpc1_1 gpc2917 (
      {stage1_4[219]},
      {stage2_4[93]}
   );
   gpc1_1 gpc2918 (
      {stage1_4[220]},
      {stage2_4[94]}
   );
   gpc1_1 gpc2919 (
      {stage1_4[221]},
      {stage2_4[95]}
   );
   gpc1_1 gpc2920 (
      {stage1_4[222]},
      {stage2_4[96]}
   );
   gpc1_1 gpc2921 (
      {stage1_4[223]},
      {stage2_4[97]}
   );
   gpc1_1 gpc2922 (
      {stage1_4[224]},
      {stage2_4[98]}
   );
   gpc1_1 gpc2923 (
      {stage1_4[225]},
      {stage2_4[99]}
   );
   gpc1_1 gpc2924 (
      {stage1_4[226]},
      {stage2_4[100]}
   );
   gpc1_1 gpc2925 (
      {stage1_4[227]},
      {stage2_4[101]}
   );
   gpc1_1 gpc2926 (
      {stage1_4[228]},
      {stage2_4[102]}
   );
   gpc1_1 gpc2927 (
      {stage1_4[229]},
      {stage2_4[103]}
   );
   gpc1_1 gpc2928 (
      {stage1_4[230]},
      {stage2_4[104]}
   );
   gpc1_1 gpc2929 (
      {stage1_4[231]},
      {stage2_4[105]}
   );
   gpc1_1 gpc2930 (
      {stage1_4[232]},
      {stage2_4[106]}
   );
   gpc1_1 gpc2931 (
      {stage1_4[233]},
      {stage2_4[107]}
   );
   gpc1_1 gpc2932 (
      {stage1_4[234]},
      {stage2_4[108]}
   );
   gpc1_1 gpc2933 (
      {stage1_4[235]},
      {stage2_4[109]}
   );
   gpc1_1 gpc2934 (
      {stage1_4[236]},
      {stage2_4[110]}
   );
   gpc1_1 gpc2935 (
      {stage1_4[237]},
      {stage2_4[111]}
   );
   gpc1_1 gpc2936 (
      {stage1_4[238]},
      {stage2_4[112]}
   );
   gpc1_1 gpc2937 (
      {stage1_4[239]},
      {stage2_4[113]}
   );
   gpc1_1 gpc2938 (
      {stage1_4[240]},
      {stage2_4[114]}
   );
   gpc1_1 gpc2939 (
      {stage1_4[241]},
      {stage2_4[115]}
   );
   gpc1_1 gpc2940 (
      {stage1_4[242]},
      {stage2_4[116]}
   );
   gpc1_1 gpc2941 (
      {stage1_4[243]},
      {stage2_4[117]}
   );
   gpc1_1 gpc2942 (
      {stage1_4[244]},
      {stage2_4[118]}
   );
   gpc1_1 gpc2943 (
      {stage1_7[166]},
      {stage2_7[89]}
   );
   gpc1_1 gpc2944 (
      {stage1_7[167]},
      {stage2_7[90]}
   );
   gpc1_1 gpc2945 (
      {stage1_7[168]},
      {stage2_7[91]}
   );
   gpc1_1 gpc2946 (
      {stage1_7[169]},
      {stage2_7[92]}
   );
   gpc1_1 gpc2947 (
      {stage1_7[170]},
      {stage2_7[93]}
   );
   gpc1_1 gpc2948 (
      {stage1_7[171]},
      {stage2_7[94]}
   );
   gpc1_1 gpc2949 (
      {stage1_7[172]},
      {stage2_7[95]}
   );
   gpc1_1 gpc2950 (
      {stage1_7[173]},
      {stage2_7[96]}
   );
   gpc1_1 gpc2951 (
      {stage1_7[174]},
      {stage2_7[97]}
   );
   gpc1_1 gpc2952 (
      {stage1_7[175]},
      {stage2_7[98]}
   );
   gpc1_1 gpc2953 (
      {stage1_7[176]},
      {stage2_7[99]}
   );
   gpc1_1 gpc2954 (
      {stage1_7[177]},
      {stage2_7[100]}
   );
   gpc1_1 gpc2955 (
      {stage1_7[178]},
      {stage2_7[101]}
   );
   gpc1_1 gpc2956 (
      {stage1_7[179]},
      {stage2_7[102]}
   );
   gpc1_1 gpc2957 (
      {stage1_7[180]},
      {stage2_7[103]}
   );
   gpc1_1 gpc2958 (
      {stage1_7[181]},
      {stage2_7[104]}
   );
   gpc1_1 gpc2959 (
      {stage1_7[182]},
      {stage2_7[105]}
   );
   gpc1_1 gpc2960 (
      {stage1_7[183]},
      {stage2_7[106]}
   );
   gpc1_1 gpc2961 (
      {stage1_7[184]},
      {stage2_7[107]}
   );
   gpc1_1 gpc2962 (
      {stage1_7[185]},
      {stage2_7[108]}
   );
   gpc1_1 gpc2963 (
      {stage1_9[210]},
      {stage2_9[106]}
   );
   gpc1_1 gpc2964 (
      {stage1_9[211]},
      {stage2_9[107]}
   );
   gpc1_1 gpc2965 (
      {stage1_11[161]},
      {stage2_11[71]}
   );
   gpc1_1 gpc2966 (
      {stage1_11[162]},
      {stage2_11[72]}
   );
   gpc1_1 gpc2967 (
      {stage1_11[163]},
      {stage2_11[73]}
   );
   gpc1_1 gpc2968 (
      {stage1_11[164]},
      {stage2_11[74]}
   );
   gpc1_1 gpc2969 (
      {stage1_11[165]},
      {stage2_11[75]}
   );
   gpc1_1 gpc2970 (
      {stage1_11[166]},
      {stage2_11[76]}
   );
   gpc1_1 gpc2971 (
      {stage1_11[167]},
      {stage2_11[77]}
   );
   gpc1_1 gpc2972 (
      {stage1_11[168]},
      {stage2_11[78]}
   );
   gpc1_1 gpc2973 (
      {stage1_11[169]},
      {stage2_11[79]}
   );
   gpc1_1 gpc2974 (
      {stage1_11[170]},
      {stage2_11[80]}
   );
   gpc1_1 gpc2975 (
      {stage1_11[171]},
      {stage2_11[81]}
   );
   gpc1_1 gpc2976 (
      {stage1_11[172]},
      {stage2_11[82]}
   );
   gpc1_1 gpc2977 (
      {stage1_11[173]},
      {stage2_11[83]}
   );
   gpc1_1 gpc2978 (
      {stage1_11[174]},
      {stage2_11[84]}
   );
   gpc1_1 gpc2979 (
      {stage1_11[175]},
      {stage2_11[85]}
   );
   gpc1_1 gpc2980 (
      {stage1_11[176]},
      {stage2_11[86]}
   );
   gpc1_1 gpc2981 (
      {stage1_11[177]},
      {stage2_11[87]}
   );
   gpc1_1 gpc2982 (
      {stage1_11[178]},
      {stage2_11[88]}
   );
   gpc1_1 gpc2983 (
      {stage1_11[179]},
      {stage2_11[89]}
   );
   gpc1_1 gpc2984 (
      {stage1_11[180]},
      {stage2_11[90]}
   );
   gpc1_1 gpc2985 (
      {stage1_11[181]},
      {stage2_11[91]}
   );
   gpc1_1 gpc2986 (
      {stage1_11[182]},
      {stage2_11[92]}
   );
   gpc1_1 gpc2987 (
      {stage1_11[183]},
      {stage2_11[93]}
   );
   gpc1_1 gpc2988 (
      {stage1_11[184]},
      {stage2_11[94]}
   );
   gpc1_1 gpc2989 (
      {stage1_11[185]},
      {stage2_11[95]}
   );
   gpc1_1 gpc2990 (
      {stage1_11[186]},
      {stage2_11[96]}
   );
   gpc1_1 gpc2991 (
      {stage1_11[187]},
      {stage2_11[97]}
   );
   gpc1_1 gpc2992 (
      {stage1_11[188]},
      {stage2_11[98]}
   );
   gpc1_1 gpc2993 (
      {stage1_11[189]},
      {stage2_11[99]}
   );
   gpc1_1 gpc2994 (
      {stage1_11[190]},
      {stage2_11[100]}
   );
   gpc1_1 gpc2995 (
      {stage1_11[191]},
      {stage2_11[101]}
   );
   gpc1_1 gpc2996 (
      {stage1_11[192]},
      {stage2_11[102]}
   );
   gpc1_1 gpc2997 (
      {stage1_11[193]},
      {stage2_11[103]}
   );
   gpc1_1 gpc2998 (
      {stage1_11[194]},
      {stage2_11[104]}
   );
   gpc1_1 gpc2999 (
      {stage1_11[195]},
      {stage2_11[105]}
   );
   gpc1_1 gpc3000 (
      {stage1_11[196]},
      {stage2_11[106]}
   );
   gpc1_1 gpc3001 (
      {stage1_11[197]},
      {stage2_11[107]}
   );
   gpc1_1 gpc3002 (
      {stage1_11[198]},
      {stage2_11[108]}
   );
   gpc1_1 gpc3003 (
      {stage1_11[199]},
      {stage2_11[109]}
   );
   gpc1_1 gpc3004 (
      {stage1_11[200]},
      {stage2_11[110]}
   );
   gpc1_1 gpc3005 (
      {stage1_11[201]},
      {stage2_11[111]}
   );
   gpc1_1 gpc3006 (
      {stage1_11[202]},
      {stage2_11[112]}
   );
   gpc1_1 gpc3007 (
      {stage1_11[203]},
      {stage2_11[113]}
   );
   gpc1_1 gpc3008 (
      {stage1_11[204]},
      {stage2_11[114]}
   );
   gpc1_1 gpc3009 (
      {stage1_11[205]},
      {stage2_11[115]}
   );
   gpc1_1 gpc3010 (
      {stage1_12[215]},
      {stage2_12[95]}
   );
   gpc1_1 gpc3011 (
      {stage1_12[216]},
      {stage2_12[96]}
   );
   gpc1_1 gpc3012 (
      {stage1_12[217]},
      {stage2_12[97]}
   );
   gpc1_1 gpc3013 (
      {stage1_12[218]},
      {stage2_12[98]}
   );
   gpc1_1 gpc3014 (
      {stage1_12[219]},
      {stage2_12[99]}
   );
   gpc1_1 gpc3015 (
      {stage1_12[220]},
      {stage2_12[100]}
   );
   gpc1_1 gpc3016 (
      {stage1_12[221]},
      {stage2_12[101]}
   );
   gpc1_1 gpc3017 (
      {stage1_13[198]},
      {stage2_13[90]}
   );
   gpc1_1 gpc3018 (
      {stage1_13[199]},
      {stage2_13[91]}
   );
   gpc1_1 gpc3019 (
      {stage1_13[200]},
      {stage2_13[92]}
   );
   gpc1_1 gpc3020 (
      {stage1_13[201]},
      {stage2_13[93]}
   );
   gpc1_1 gpc3021 (
      {stage1_13[202]},
      {stage2_13[94]}
   );
   gpc1_1 gpc3022 (
      {stage1_13[203]},
      {stage2_13[95]}
   );
   gpc1_1 gpc3023 (
      {stage1_13[204]},
      {stage2_13[96]}
   );
   gpc1_1 gpc3024 (
      {stage1_13[205]},
      {stage2_13[97]}
   );
   gpc1_1 gpc3025 (
      {stage1_13[206]},
      {stage2_13[98]}
   );
   gpc1_1 gpc3026 (
      {stage1_13[207]},
      {stage2_13[99]}
   );
   gpc1_1 gpc3027 (
      {stage1_13[208]},
      {stage2_13[100]}
   );
   gpc1_1 gpc3028 (
      {stage1_13[209]},
      {stage2_13[101]}
   );
   gpc1_1 gpc3029 (
      {stage1_13[210]},
      {stage2_13[102]}
   );
   gpc1_1 gpc3030 (
      {stage1_13[211]},
      {stage2_13[103]}
   );
   gpc1_1 gpc3031 (
      {stage1_13[212]},
      {stage2_13[104]}
   );
   gpc1_1 gpc3032 (
      {stage1_13[213]},
      {stage2_13[105]}
   );
   gpc1_1 gpc3033 (
      {stage1_13[214]},
      {stage2_13[106]}
   );
   gpc1_1 gpc3034 (
      {stage1_13[215]},
      {stage2_13[107]}
   );
   gpc1_1 gpc3035 (
      {stage1_13[216]},
      {stage2_13[108]}
   );
   gpc1_1 gpc3036 (
      {stage1_13[217]},
      {stage2_13[109]}
   );
   gpc1_1 gpc3037 (
      {stage1_13[218]},
      {stage2_13[110]}
   );
   gpc1_1 gpc3038 (
      {stage1_13[219]},
      {stage2_13[111]}
   );
   gpc1_1 gpc3039 (
      {stage1_13[220]},
      {stage2_13[112]}
   );
   gpc1_1 gpc3040 (
      {stage1_13[221]},
      {stage2_13[113]}
   );
   gpc1_1 gpc3041 (
      {stage1_13[222]},
      {stage2_13[114]}
   );
   gpc1_1 gpc3042 (
      {stage1_13[223]},
      {stage2_13[115]}
   );
   gpc1_1 gpc3043 (
      {stage1_13[224]},
      {stage2_13[116]}
   );
   gpc1_1 gpc3044 (
      {stage1_13[225]},
      {stage2_13[117]}
   );
   gpc1_1 gpc3045 (
      {stage1_13[226]},
      {stage2_13[118]}
   );
   gpc1_1 gpc3046 (
      {stage1_13[227]},
      {stage2_13[119]}
   );
   gpc1_1 gpc3047 (
      {stage1_13[228]},
      {stage2_13[120]}
   );
   gpc1_1 gpc3048 (
      {stage1_13[229]},
      {stage2_13[121]}
   );
   gpc1_1 gpc3049 (
      {stage1_13[230]},
      {stage2_13[122]}
   );
   gpc1_1 gpc3050 (
      {stage1_13[231]},
      {stage2_13[123]}
   );
   gpc1_1 gpc3051 (
      {stage1_15[222]},
      {stage2_15[83]}
   );
   gpc1_1 gpc3052 (
      {stage1_15[223]},
      {stage2_15[84]}
   );
   gpc1_1 gpc3053 (
      {stage1_15[224]},
      {stage2_15[85]}
   );
   gpc1_1 gpc3054 (
      {stage1_15[225]},
      {stage2_15[86]}
   );
   gpc1_1 gpc3055 (
      {stage1_15[226]},
      {stage2_15[87]}
   );
   gpc1_1 gpc3056 (
      {stage1_15[227]},
      {stage2_15[88]}
   );
   gpc1_1 gpc3057 (
      {stage1_15[228]},
      {stage2_15[89]}
   );
   gpc1_1 gpc3058 (
      {stage1_15[229]},
      {stage2_15[90]}
   );
   gpc1_1 gpc3059 (
      {stage1_15[230]},
      {stage2_15[91]}
   );
   gpc1_1 gpc3060 (
      {stage1_15[231]},
      {stage2_15[92]}
   );
   gpc1_1 gpc3061 (
      {stage1_15[232]},
      {stage2_15[93]}
   );
   gpc1_1 gpc3062 (
      {stage1_15[233]},
      {stage2_15[94]}
   );
   gpc1_1 gpc3063 (
      {stage1_15[234]},
      {stage2_15[95]}
   );
   gpc1_1 gpc3064 (
      {stage1_15[235]},
      {stage2_15[96]}
   );
   gpc1_1 gpc3065 (
      {stage1_15[236]},
      {stage2_15[97]}
   );
   gpc1_1 gpc3066 (
      {stage1_16[196]},
      {stage2_16[107]}
   );
   gpc1_1 gpc3067 (
      {stage1_16[197]},
      {stage2_16[108]}
   );
   gpc1_1 gpc3068 (
      {stage1_16[198]},
      {stage2_16[109]}
   );
   gpc1_1 gpc3069 (
      {stage1_16[199]},
      {stage2_16[110]}
   );
   gpc1_1 gpc3070 (
      {stage1_16[200]},
      {stage2_16[111]}
   );
   gpc1_1 gpc3071 (
      {stage1_16[201]},
      {stage2_16[112]}
   );
   gpc1_1 gpc3072 (
      {stage1_16[202]},
      {stage2_16[113]}
   );
   gpc1_1 gpc3073 (
      {stage1_16[203]},
      {stage2_16[114]}
   );
   gpc1_1 gpc3074 (
      {stage1_16[204]},
      {stage2_16[115]}
   );
   gpc1_1 gpc3075 (
      {stage1_16[205]},
      {stage2_16[116]}
   );
   gpc1_1 gpc3076 (
      {stage1_16[206]},
      {stage2_16[117]}
   );
   gpc1_1 gpc3077 (
      {stage1_16[207]},
      {stage2_16[118]}
   );
   gpc1_1 gpc3078 (
      {stage1_16[208]},
      {stage2_16[119]}
   );
   gpc1_1 gpc3079 (
      {stage1_16[209]},
      {stage2_16[120]}
   );
   gpc1_1 gpc3080 (
      {stage1_16[210]},
      {stage2_16[121]}
   );
   gpc1_1 gpc3081 (
      {stage1_16[211]},
      {stage2_16[122]}
   );
   gpc1_1 gpc3082 (
      {stage1_16[212]},
      {stage2_16[123]}
   );
   gpc1_1 gpc3083 (
      {stage1_16[213]},
      {stage2_16[124]}
   );
   gpc1_1 gpc3084 (
      {stage1_17[178]},
      {stage2_17[82]}
   );
   gpc1_1 gpc3085 (
      {stage1_17[179]},
      {stage2_17[83]}
   );
   gpc1_1 gpc3086 (
      {stage1_17[180]},
      {stage2_17[84]}
   );
   gpc1_1 gpc3087 (
      {stage1_17[181]},
      {stage2_17[85]}
   );
   gpc1_1 gpc3088 (
      {stage1_17[182]},
      {stage2_17[86]}
   );
   gpc1_1 gpc3089 (
      {stage1_17[183]},
      {stage2_17[87]}
   );
   gpc1_1 gpc3090 (
      {stage1_17[184]},
      {stage2_17[88]}
   );
   gpc1_1 gpc3091 (
      {stage1_17[185]},
      {stage2_17[89]}
   );
   gpc1_1 gpc3092 (
      {stage1_17[186]},
      {stage2_17[90]}
   );
   gpc1_1 gpc3093 (
      {stage1_17[187]},
      {stage2_17[91]}
   );
   gpc1_1 gpc3094 (
      {stage1_17[188]},
      {stage2_17[92]}
   );
   gpc1_1 gpc3095 (
      {stage1_17[189]},
      {stage2_17[93]}
   );
   gpc1_1 gpc3096 (
      {stage1_17[190]},
      {stage2_17[94]}
   );
   gpc1_1 gpc3097 (
      {stage1_17[191]},
      {stage2_17[95]}
   );
   gpc1_1 gpc3098 (
      {stage1_17[192]},
      {stage2_17[96]}
   );
   gpc1_1 gpc3099 (
      {stage1_17[193]},
      {stage2_17[97]}
   );
   gpc1_1 gpc3100 (
      {stage1_17[194]},
      {stage2_17[98]}
   );
   gpc1_1 gpc3101 (
      {stage1_17[195]},
      {stage2_17[99]}
   );
   gpc1_1 gpc3102 (
      {stage1_17[196]},
      {stage2_17[100]}
   );
   gpc1_1 gpc3103 (
      {stage1_17[197]},
      {stage2_17[101]}
   );
   gpc1_1 gpc3104 (
      {stage1_17[198]},
      {stage2_17[102]}
   );
   gpc1_1 gpc3105 (
      {stage1_17[199]},
      {stage2_17[103]}
   );
   gpc1_1 gpc3106 (
      {stage1_17[200]},
      {stage2_17[104]}
   );
   gpc1_1 gpc3107 (
      {stage1_17[201]},
      {stage2_17[105]}
   );
   gpc1_1 gpc3108 (
      {stage1_17[202]},
      {stage2_17[106]}
   );
   gpc1_1 gpc3109 (
      {stage1_17[203]},
      {stage2_17[107]}
   );
   gpc1_1 gpc3110 (
      {stage1_17[204]},
      {stage2_17[108]}
   );
   gpc1_1 gpc3111 (
      {stage1_17[205]},
      {stage2_17[109]}
   );
   gpc1_1 gpc3112 (
      {stage1_17[206]},
      {stage2_17[110]}
   );
   gpc1_1 gpc3113 (
      {stage1_17[207]},
      {stage2_17[111]}
   );
   gpc1_1 gpc3114 (
      {stage1_17[208]},
      {stage2_17[112]}
   );
   gpc1_1 gpc3115 (
      {stage1_17[209]},
      {stage2_17[113]}
   );
   gpc1_1 gpc3116 (
      {stage1_17[210]},
      {stage2_17[114]}
   );
   gpc1_1 gpc3117 (
      {stage1_17[211]},
      {stage2_17[115]}
   );
   gpc1_1 gpc3118 (
      {stage1_17[212]},
      {stage2_17[116]}
   );
   gpc1_1 gpc3119 (
      {stage1_17[213]},
      {stage2_17[117]}
   );
   gpc1_1 gpc3120 (
      {stage1_17[214]},
      {stage2_17[118]}
   );
   gpc1_1 gpc3121 (
      {stage1_17[215]},
      {stage2_17[119]}
   );
   gpc1_1 gpc3122 (
      {stage1_17[216]},
      {stage2_17[120]}
   );
   gpc1_1 gpc3123 (
      {stage1_17[217]},
      {stage2_17[121]}
   );
   gpc1_1 gpc3124 (
      {stage1_17[218]},
      {stage2_17[122]}
   );
   gpc1_1 gpc3125 (
      {stage1_17[219]},
      {stage2_17[123]}
   );
   gpc1_1 gpc3126 (
      {stage1_17[220]},
      {stage2_17[124]}
   );
   gpc1_1 gpc3127 (
      {stage1_17[221]},
      {stage2_17[125]}
   );
   gpc1_1 gpc3128 (
      {stage1_17[222]},
      {stage2_17[126]}
   );
   gpc1_1 gpc3129 (
      {stage1_17[223]},
      {stage2_17[127]}
   );
   gpc1_1 gpc3130 (
      {stage1_18[194]},
      {stage2_18[64]}
   );
   gpc1_1 gpc3131 (
      {stage1_18[195]},
      {stage2_18[65]}
   );
   gpc1_1 gpc3132 (
      {stage1_18[196]},
      {stage2_18[66]}
   );
   gpc1_1 gpc3133 (
      {stage1_18[197]},
      {stage2_18[67]}
   );
   gpc1_1 gpc3134 (
      {stage1_18[198]},
      {stage2_18[68]}
   );
   gpc1_1 gpc3135 (
      {stage1_18[199]},
      {stage2_18[69]}
   );
   gpc1_1 gpc3136 (
      {stage1_18[200]},
      {stage2_18[70]}
   );
   gpc1_1 gpc3137 (
      {stage1_18[201]},
      {stage2_18[71]}
   );
   gpc1_1 gpc3138 (
      {stage1_18[202]},
      {stage2_18[72]}
   );
   gpc1_1 gpc3139 (
      {stage1_19[261]},
      {stage2_19[96]}
   );
   gpc1_1 gpc3140 (
      {stage1_19[262]},
      {stage2_19[97]}
   );
   gpc1_1 gpc3141 (
      {stage1_20[211]},
      {stage2_20[107]}
   );
   gpc1_1 gpc3142 (
      {stage1_20[212]},
      {stage2_20[108]}
   );
   gpc1_1 gpc3143 (
      {stage1_20[213]},
      {stage2_20[109]}
   );
   gpc1_1 gpc3144 (
      {stage1_21[227]},
      {stage2_21[82]}
   );
   gpc1_1 gpc3145 (
      {stage1_21[228]},
      {stage2_21[83]}
   );
   gpc1_1 gpc3146 (
      {stage1_21[229]},
      {stage2_21[84]}
   );
   gpc1_1 gpc3147 (
      {stage1_21[230]},
      {stage2_21[85]}
   );
   gpc1_1 gpc3148 (
      {stage1_21[231]},
      {stage2_21[86]}
   );
   gpc1_1 gpc3149 (
      {stage1_21[232]},
      {stage2_21[87]}
   );
   gpc1_1 gpc3150 (
      {stage1_21[233]},
      {stage2_21[88]}
   );
   gpc1_1 gpc3151 (
      {stage1_21[234]},
      {stage2_21[89]}
   );
   gpc1_1 gpc3152 (
      {stage1_21[235]},
      {stage2_21[90]}
   );
   gpc1_1 gpc3153 (
      {stage1_21[236]},
      {stage2_21[91]}
   );
   gpc1_1 gpc3154 (
      {stage1_21[237]},
      {stage2_21[92]}
   );
   gpc1_1 gpc3155 (
      {stage1_21[238]},
      {stage2_21[93]}
   );
   gpc1_1 gpc3156 (
      {stage1_21[239]},
      {stage2_21[94]}
   );
   gpc1_1 gpc3157 (
      {stage1_21[240]},
      {stage2_21[95]}
   );
   gpc1_1 gpc3158 (
      {stage1_21[241]},
      {stage2_21[96]}
   );
   gpc1_1 gpc3159 (
      {stage1_21[242]},
      {stage2_21[97]}
   );
   gpc1_1 gpc3160 (
      {stage1_21[243]},
      {stage2_21[98]}
   );
   gpc1_1 gpc3161 (
      {stage1_21[244]},
      {stage2_21[99]}
   );
   gpc1_1 gpc3162 (
      {stage1_21[245]},
      {stage2_21[100]}
   );
   gpc1_1 gpc3163 (
      {stage1_21[246]},
      {stage2_21[101]}
   );
   gpc1_1 gpc3164 (
      {stage1_21[247]},
      {stage2_21[102]}
   );
   gpc1_1 gpc3165 (
      {stage1_21[248]},
      {stage2_21[103]}
   );
   gpc1_1 gpc3166 (
      {stage1_21[249]},
      {stage2_21[104]}
   );
   gpc1_1 gpc3167 (
      {stage1_21[250]},
      {stage2_21[105]}
   );
   gpc1_1 gpc3168 (
      {stage1_21[251]},
      {stage2_21[106]}
   );
   gpc1_1 gpc3169 (
      {stage1_21[252]},
      {stage2_21[107]}
   );
   gpc1_1 gpc3170 (
      {stage1_21[253]},
      {stage2_21[108]}
   );
   gpc1_1 gpc3171 (
      {stage1_21[254]},
      {stage2_21[109]}
   );
   gpc1_1 gpc3172 (
      {stage1_21[255]},
      {stage2_21[110]}
   );
   gpc1_1 gpc3173 (
      {stage1_21[256]},
      {stage2_21[111]}
   );
   gpc1_1 gpc3174 (
      {stage1_21[257]},
      {stage2_21[112]}
   );
   gpc1_1 gpc3175 (
      {stage1_21[258]},
      {stage2_21[113]}
   );
   gpc1_1 gpc3176 (
      {stage1_21[259]},
      {stage2_21[114]}
   );
   gpc1_1 gpc3177 (
      {stage1_21[260]},
      {stage2_21[115]}
   );
   gpc1_1 gpc3178 (
      {stage1_21[261]},
      {stage2_21[116]}
   );
   gpc1_1 gpc3179 (
      {stage1_21[262]},
      {stage2_21[117]}
   );
   gpc1_1 gpc3180 (
      {stage1_21[263]},
      {stage2_21[118]}
   );
   gpc1_1 gpc3181 (
      {stage1_21[264]},
      {stage2_21[119]}
   );
   gpc1_1 gpc3182 (
      {stage1_21[265]},
      {stage2_21[120]}
   );
   gpc1_1 gpc3183 (
      {stage1_21[266]},
      {stage2_21[121]}
   );
   gpc1_1 gpc3184 (
      {stage1_21[267]},
      {stage2_21[122]}
   );
   gpc1_1 gpc3185 (
      {stage1_21[268]},
      {stage2_21[123]}
   );
   gpc1_1 gpc3186 (
      {stage1_21[269]},
      {stage2_21[124]}
   );
   gpc1_1 gpc3187 (
      {stage1_22[268]},
      {stage2_22[89]}
   );
   gpc1_1 gpc3188 (
      {stage1_22[269]},
      {stage2_22[90]}
   );
   gpc1_1 gpc3189 (
      {stage1_22[270]},
      {stage2_22[91]}
   );
   gpc1_1 gpc3190 (
      {stage1_22[271]},
      {stage2_22[92]}
   );
   gpc1_1 gpc3191 (
      {stage1_22[272]},
      {stage2_22[93]}
   );
   gpc1_1 gpc3192 (
      {stage1_22[273]},
      {stage2_22[94]}
   );
   gpc1_1 gpc3193 (
      {stage1_23[146]},
      {stage2_23[103]}
   );
   gpc1_1 gpc3194 (
      {stage1_23[147]},
      {stage2_23[104]}
   );
   gpc1_1 gpc3195 (
      {stage1_23[148]},
      {stage2_23[105]}
   );
   gpc1_1 gpc3196 (
      {stage1_23[149]},
      {stage2_23[106]}
   );
   gpc1_1 gpc3197 (
      {stage1_23[150]},
      {stage2_23[107]}
   );
   gpc1_1 gpc3198 (
      {stage1_23[151]},
      {stage2_23[108]}
   );
   gpc1_1 gpc3199 (
      {stage1_23[152]},
      {stage2_23[109]}
   );
   gpc1_1 gpc3200 (
      {stage1_23[153]},
      {stage2_23[110]}
   );
   gpc1_1 gpc3201 (
      {stage1_23[154]},
      {stage2_23[111]}
   );
   gpc1_1 gpc3202 (
      {stage1_23[155]},
      {stage2_23[112]}
   );
   gpc1_1 gpc3203 (
      {stage1_23[156]},
      {stage2_23[113]}
   );
   gpc1_1 gpc3204 (
      {stage1_23[157]},
      {stage2_23[114]}
   );
   gpc1_1 gpc3205 (
      {stage1_23[158]},
      {stage2_23[115]}
   );
   gpc1_1 gpc3206 (
      {stage1_23[159]},
      {stage2_23[116]}
   );
   gpc1_1 gpc3207 (
      {stage1_23[160]},
      {stage2_23[117]}
   );
   gpc1_1 gpc3208 (
      {stage1_23[161]},
      {stage2_23[118]}
   );
   gpc1_1 gpc3209 (
      {stage1_23[162]},
      {stage2_23[119]}
   );
   gpc1_1 gpc3210 (
      {stage1_23[163]},
      {stage2_23[120]}
   );
   gpc1_1 gpc3211 (
      {stage1_23[164]},
      {stage2_23[121]}
   );
   gpc1_1 gpc3212 (
      {stage1_23[165]},
      {stage2_23[122]}
   );
   gpc1_1 gpc3213 (
      {stage1_24[217]},
      {stage2_24[86]}
   );
   gpc1_1 gpc3214 (
      {stage1_24[218]},
      {stage2_24[87]}
   );
   gpc1_1 gpc3215 (
      {stage1_24[219]},
      {stage2_24[88]}
   );
   gpc1_1 gpc3216 (
      {stage1_24[220]},
      {stage2_24[89]}
   );
   gpc1_1 gpc3217 (
      {stage1_25[255]},
      {stage2_25[84]}
   );
   gpc1_1 gpc3218 (
      {stage1_25[256]},
      {stage2_25[85]}
   );
   gpc1_1 gpc3219 (
      {stage1_25[257]},
      {stage2_25[86]}
   );
   gpc1_1 gpc3220 (
      {stage1_25[258]},
      {stage2_25[87]}
   );
   gpc1_1 gpc3221 (
      {stage1_25[259]},
      {stage2_25[88]}
   );
   gpc1_1 gpc3222 (
      {stage1_25[260]},
      {stage2_25[89]}
   );
   gpc1_1 gpc3223 (
      {stage1_25[261]},
      {stage2_25[90]}
   );
   gpc1_1 gpc3224 (
      {stage1_25[262]},
      {stage2_25[91]}
   );
   gpc1_1 gpc3225 (
      {stage1_25[263]},
      {stage2_25[92]}
   );
   gpc1_1 gpc3226 (
      {stage1_25[264]},
      {stage2_25[93]}
   );
   gpc1_1 gpc3227 (
      {stage1_25[265]},
      {stage2_25[94]}
   );
   gpc1_1 gpc3228 (
      {stage1_25[266]},
      {stage2_25[95]}
   );
   gpc1_1 gpc3229 (
      {stage1_25[267]},
      {stage2_25[96]}
   );
   gpc1_1 gpc3230 (
      {stage1_25[268]},
      {stage2_25[97]}
   );
   gpc1_1 gpc3231 (
      {stage1_25[269]},
      {stage2_25[98]}
   );
   gpc1_1 gpc3232 (
      {stage1_25[270]},
      {stage2_25[99]}
   );
   gpc1_1 gpc3233 (
      {stage1_25[271]},
      {stage2_25[100]}
   );
   gpc1_1 gpc3234 (
      {stage1_25[272]},
      {stage2_25[101]}
   );
   gpc1_1 gpc3235 (
      {stage1_25[273]},
      {stage2_25[102]}
   );
   gpc1_1 gpc3236 (
      {stage1_26[186]},
      {stage2_26[95]}
   );
   gpc1_1 gpc3237 (
      {stage1_26[187]},
      {stage2_26[96]}
   );
   gpc1_1 gpc3238 (
      {stage1_26[188]},
      {stage2_26[97]}
   );
   gpc1_1 gpc3239 (
      {stage1_26[189]},
      {stage2_26[98]}
   );
   gpc1_1 gpc3240 (
      {stage1_26[190]},
      {stage2_26[99]}
   );
   gpc1_1 gpc3241 (
      {stage1_27[196]},
      {stage2_27[81]}
   );
   gpc1_1 gpc3242 (
      {stage1_27[197]},
      {stage2_27[82]}
   );
   gpc1_1 gpc3243 (
      {stage1_27[198]},
      {stage2_27[83]}
   );
   gpc1_1 gpc3244 (
      {stage1_27[199]},
      {stage2_27[84]}
   );
   gpc1_1 gpc3245 (
      {stage1_28[149]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3246 (
      {stage1_28[150]},
      {stage2_28[73]}
   );
   gpc1_1 gpc3247 (
      {stage1_28[151]},
      {stage2_28[74]}
   );
   gpc1_1 gpc3248 (
      {stage1_28[152]},
      {stage2_28[75]}
   );
   gpc1_1 gpc3249 (
      {stage1_28[153]},
      {stage2_28[76]}
   );
   gpc1_1 gpc3250 (
      {stage1_28[154]},
      {stage2_28[77]}
   );
   gpc1_1 gpc3251 (
      {stage1_28[155]},
      {stage2_28[78]}
   );
   gpc1_1 gpc3252 (
      {stage1_28[156]},
      {stage2_28[79]}
   );
   gpc1_1 gpc3253 (
      {stage1_28[157]},
      {stage2_28[80]}
   );
   gpc1_1 gpc3254 (
      {stage1_28[158]},
      {stage2_28[81]}
   );
   gpc1_1 gpc3255 (
      {stage1_28[159]},
      {stage2_28[82]}
   );
   gpc1_1 gpc3256 (
      {stage1_28[160]},
      {stage2_28[83]}
   );
   gpc1_1 gpc3257 (
      {stage1_28[161]},
      {stage2_28[84]}
   );
   gpc1_1 gpc3258 (
      {stage1_28[162]},
      {stage2_28[85]}
   );
   gpc1_1 gpc3259 (
      {stage1_28[163]},
      {stage2_28[86]}
   );
   gpc1_1 gpc3260 (
      {stage1_28[164]},
      {stage2_28[87]}
   );
   gpc1_1 gpc3261 (
      {stage1_28[165]},
      {stage2_28[88]}
   );
   gpc1_1 gpc3262 (
      {stage1_28[166]},
      {stage2_28[89]}
   );
   gpc1_1 gpc3263 (
      {stage1_28[167]},
      {stage2_28[90]}
   );
   gpc1_1 gpc3264 (
      {stage1_28[168]},
      {stage2_28[91]}
   );
   gpc1_1 gpc3265 (
      {stage1_28[169]},
      {stage2_28[92]}
   );
   gpc1_1 gpc3266 (
      {stage1_28[170]},
      {stage2_28[93]}
   );
   gpc1_1 gpc3267 (
      {stage1_28[171]},
      {stage2_28[94]}
   );
   gpc1_1 gpc3268 (
      {stage1_28[172]},
      {stage2_28[95]}
   );
   gpc1_1 gpc3269 (
      {stage1_28[173]},
      {stage2_28[96]}
   );
   gpc1_1 gpc3270 (
      {stage1_28[174]},
      {stage2_28[97]}
   );
   gpc1_1 gpc3271 (
      {stage1_28[175]},
      {stage2_28[98]}
   );
   gpc1_1 gpc3272 (
      {stage1_28[176]},
      {stage2_28[99]}
   );
   gpc1_1 gpc3273 (
      {stage1_28[177]},
      {stage2_28[100]}
   );
   gpc1_1 gpc3274 (
      {stage1_28[178]},
      {stage2_28[101]}
   );
   gpc1_1 gpc3275 (
      {stage1_28[179]},
      {stage2_28[102]}
   );
   gpc1_1 gpc3276 (
      {stage1_28[180]},
      {stage2_28[103]}
   );
   gpc1_1 gpc3277 (
      {stage1_28[181]},
      {stage2_28[104]}
   );
   gpc1_1 gpc3278 (
      {stage1_28[182]},
      {stage2_28[105]}
   );
   gpc1_1 gpc3279 (
      {stage1_28[183]},
      {stage2_28[106]}
   );
   gpc1_1 gpc3280 (
      {stage1_28[184]},
      {stage2_28[107]}
   );
   gpc1_1 gpc3281 (
      {stage1_28[185]},
      {stage2_28[108]}
   );
   gpc1_1 gpc3282 (
      {stage1_28[186]},
      {stage2_28[109]}
   );
   gpc1_1 gpc3283 (
      {stage1_28[187]},
      {stage2_28[110]}
   );
   gpc1_1 gpc3284 (
      {stage1_28[188]},
      {stage2_28[111]}
   );
   gpc1_1 gpc3285 (
      {stage1_28[189]},
      {stage2_28[112]}
   );
   gpc1_1 gpc3286 (
      {stage1_28[190]},
      {stage2_28[113]}
   );
   gpc1_1 gpc3287 (
      {stage1_28[191]},
      {stage2_28[114]}
   );
   gpc1_1 gpc3288 (
      {stage1_28[192]},
      {stage2_28[115]}
   );
   gpc1_1 gpc3289 (
      {stage1_28[193]},
      {stage2_28[116]}
   );
   gpc1_1 gpc3290 (
      {stage1_28[194]},
      {stage2_28[117]}
   );
   gpc1_1 gpc3291 (
      {stage1_28[195]},
      {stage2_28[118]}
   );
   gpc1_1 gpc3292 (
      {stage1_28[196]},
      {stage2_28[119]}
   );
   gpc1_1 gpc3293 (
      {stage1_28[197]},
      {stage2_28[120]}
   );
   gpc1_1 gpc3294 (
      {stage1_28[198]},
      {stage2_28[121]}
   );
   gpc1_1 gpc3295 (
      {stage1_28[199]},
      {stage2_28[122]}
   );
   gpc1_1 gpc3296 (
      {stage1_28[200]},
      {stage2_28[123]}
   );
   gpc1_1 gpc3297 (
      {stage1_28[201]},
      {stage2_28[124]}
   );
   gpc1_1 gpc3298 (
      {stage1_28[202]},
      {stage2_28[125]}
   );
   gpc1_1 gpc3299 (
      {stage1_28[203]},
      {stage2_28[126]}
   );
   gpc1_1 gpc3300 (
      {stage1_28[204]},
      {stage2_28[127]}
   );
   gpc1_1 gpc3301 (
      {stage1_28[205]},
      {stage2_28[128]}
   );
   gpc1_1 gpc3302 (
      {stage1_28[206]},
      {stage2_28[129]}
   );
   gpc1_1 gpc3303 (
      {stage1_28[207]},
      {stage2_28[130]}
   );
   gpc1_1 gpc3304 (
      {stage1_28[208]},
      {stage2_28[131]}
   );
   gpc1_1 gpc3305 (
      {stage1_28[209]},
      {stage2_28[132]}
   );
   gpc1_1 gpc3306 (
      {stage1_28[210]},
      {stage2_28[133]}
   );
   gpc1_1 gpc3307 (
      {stage1_28[211]},
      {stage2_28[134]}
   );
   gpc1_1 gpc3308 (
      {stage1_28[212]},
      {stage2_28[135]}
   );
   gpc1_1 gpc3309 (
      {stage1_28[213]},
      {stage2_28[136]}
   );
   gpc1_1 gpc3310 (
      {stage1_28[214]},
      {stage2_28[137]}
   );
   gpc1_1 gpc3311 (
      {stage1_28[215]},
      {stage2_28[138]}
   );
   gpc1_1 gpc3312 (
      {stage1_28[216]},
      {stage2_28[139]}
   );
   gpc1_1 gpc3313 (
      {stage1_28[217]},
      {stage2_28[140]}
   );
   gpc1_1 gpc3314 (
      {stage1_28[218]},
      {stage2_28[141]}
   );
   gpc1_1 gpc3315 (
      {stage1_28[219]},
      {stage2_28[142]}
   );
   gpc1_1 gpc3316 (
      {stage1_28[220]},
      {stage2_28[143]}
   );
   gpc1_1 gpc3317 (
      {stage1_28[221]},
      {stage2_28[144]}
   );
   gpc1_1 gpc3318 (
      {stage1_28[222]},
      {stage2_28[145]}
   );
   gpc1_1 gpc3319 (
      {stage1_28[223]},
      {stage2_28[146]}
   );
   gpc1_1 gpc3320 (
      {stage1_28[224]},
      {stage2_28[147]}
   );
   gpc1_1 gpc3321 (
      {stage1_28[225]},
      {stage2_28[148]}
   );
   gpc1_1 gpc3322 (
      {stage1_28[226]},
      {stage2_28[149]}
   );
   gpc1_1 gpc3323 (
      {stage1_28[227]},
      {stage2_28[150]}
   );
   gpc1_1 gpc3324 (
      {stage1_28[228]},
      {stage2_28[151]}
   );
   gpc1_1 gpc3325 (
      {stage1_28[229]},
      {stage2_28[152]}
   );
   gpc1_1 gpc3326 (
      {stage1_28[230]},
      {stage2_28[153]}
   );
   gpc1_1 gpc3327 (
      {stage1_28[231]},
      {stage2_28[154]}
   );
   gpc1_1 gpc3328 (
      {stage1_28[232]},
      {stage2_28[155]}
   );
   gpc1_1 gpc3329 (
      {stage1_28[233]},
      {stage2_28[156]}
   );
   gpc1_1 gpc3330 (
      {stage1_28[234]},
      {stage2_28[157]}
   );
   gpc1_1 gpc3331 (
      {stage1_28[235]},
      {stage2_28[158]}
   );
   gpc1_1 gpc3332 (
      {stage1_28[236]},
      {stage2_28[159]}
   );
   gpc1_1 gpc3333 (
      {stage1_28[237]},
      {stage2_28[160]}
   );
   gpc1_1 gpc3334 (
      {stage1_28[238]},
      {stage2_28[161]}
   );
   gpc1_1 gpc3335 (
      {stage1_28[239]},
      {stage2_28[162]}
   );
   gpc1_1 gpc3336 (
      {stage1_28[240]},
      {stage2_28[163]}
   );
   gpc1_1 gpc3337 (
      {stage1_28[241]},
      {stage2_28[164]}
   );
   gpc1_1 gpc3338 (
      {stage1_28[242]},
      {stage2_28[165]}
   );
   gpc1_1 gpc3339 (
      {stage1_28[243]},
      {stage2_28[166]}
   );
   gpc1_1 gpc3340 (
      {stage1_28[244]},
      {stage2_28[167]}
   );
   gpc1_1 gpc3341 (
      {stage1_28[245]},
      {stage2_28[168]}
   );
   gpc1_1 gpc3342 (
      {stage1_28[246]},
      {stage2_28[169]}
   );
   gpc1_1 gpc3343 (
      {stage1_28[247]},
      {stage2_28[170]}
   );
   gpc1_1 gpc3344 (
      {stage1_29[180]},
      {stage2_29[80]}
   );
   gpc1_1 gpc3345 (
      {stage1_29[181]},
      {stage2_29[81]}
   );
   gpc1_1 gpc3346 (
      {stage1_29[182]},
      {stage2_29[82]}
   );
   gpc1_1 gpc3347 (
      {stage1_29[183]},
      {stage2_29[83]}
   );
   gpc1_1 gpc3348 (
      {stage1_29[184]},
      {stage2_29[84]}
   );
   gpc1_1 gpc3349 (
      {stage1_29[185]},
      {stage2_29[85]}
   );
   gpc1_1 gpc3350 (
      {stage1_29[186]},
      {stage2_29[86]}
   );
   gpc1_1 gpc3351 (
      {stage1_29[187]},
      {stage2_29[87]}
   );
   gpc1_1 gpc3352 (
      {stage1_29[188]},
      {stage2_29[88]}
   );
   gpc1_1 gpc3353 (
      {stage1_29[189]},
      {stage2_29[89]}
   );
   gpc1_1 gpc3354 (
      {stage1_29[190]},
      {stage2_29[90]}
   );
   gpc1_1 gpc3355 (
      {stage1_29[191]},
      {stage2_29[91]}
   );
   gpc1_1 gpc3356 (
      {stage1_29[192]},
      {stage2_29[92]}
   );
   gpc1_1 gpc3357 (
      {stage1_29[193]},
      {stage2_29[93]}
   );
   gpc1_1 gpc3358 (
      {stage1_29[194]},
      {stage2_29[94]}
   );
   gpc1_1 gpc3359 (
      {stage1_29[195]},
      {stage2_29[95]}
   );
   gpc1_1 gpc3360 (
      {stage1_29[196]},
      {stage2_29[96]}
   );
   gpc1_1 gpc3361 (
      {stage1_29[197]},
      {stage2_29[97]}
   );
   gpc1_1 gpc3362 (
      {stage1_29[198]},
      {stage2_29[98]}
   );
   gpc1_1 gpc3363 (
      {stage1_29[199]},
      {stage2_29[99]}
   );
   gpc1_1 gpc3364 (
      {stage1_29[200]},
      {stage2_29[100]}
   );
   gpc1_1 gpc3365 (
      {stage1_29[201]},
      {stage2_29[101]}
   );
   gpc1_1 gpc3366 (
      {stage1_29[202]},
      {stage2_29[102]}
   );
   gpc1_1 gpc3367 (
      {stage1_29[203]},
      {stage2_29[103]}
   );
   gpc1_1 gpc3368 (
      {stage1_29[204]},
      {stage2_29[104]}
   );
   gpc1_1 gpc3369 (
      {stage1_29[205]},
      {stage2_29[105]}
   );
   gpc1_1 gpc3370 (
      {stage1_29[206]},
      {stage2_29[106]}
   );
   gpc1_1 gpc3371 (
      {stage1_29[207]},
      {stage2_29[107]}
   );
   gpc1_1 gpc3372 (
      {stage1_29[208]},
      {stage2_29[108]}
   );
   gpc1_1 gpc3373 (
      {stage1_29[209]},
      {stage2_29[109]}
   );
   gpc1_1 gpc3374 (
      {stage1_29[210]},
      {stage2_29[110]}
   );
   gpc1_1 gpc3375 (
      {stage1_29[211]},
      {stage2_29[111]}
   );
   gpc1_1 gpc3376 (
      {stage1_29[212]},
      {stage2_29[112]}
   );
   gpc1_1 gpc3377 (
      {stage1_29[213]},
      {stage2_29[113]}
   );
   gpc1_1 gpc3378 (
      {stage1_29[214]},
      {stage2_29[114]}
   );
   gpc1_1 gpc3379 (
      {stage1_29[215]},
      {stage2_29[115]}
   );
   gpc1_1 gpc3380 (
      {stage1_29[216]},
      {stage2_29[116]}
   );
   gpc1_1 gpc3381 (
      {stage1_29[217]},
      {stage2_29[117]}
   );
   gpc1_1 gpc3382 (
      {stage1_29[218]},
      {stage2_29[118]}
   );
   gpc1_1 gpc3383 (
      {stage1_29[219]},
      {stage2_29[119]}
   );
   gpc1_1 gpc3384 (
      {stage1_29[220]},
      {stage2_29[120]}
   );
   gpc1_1 gpc3385 (
      {stage1_29[221]},
      {stage2_29[121]}
   );
   gpc1_1 gpc3386 (
      {stage1_29[222]},
      {stage2_29[122]}
   );
   gpc1_1 gpc3387 (
      {stage1_29[223]},
      {stage2_29[123]}
   );
   gpc1_1 gpc3388 (
      {stage1_29[224]},
      {stage2_29[124]}
   );
   gpc1_1 gpc3389 (
      {stage1_29[225]},
      {stage2_29[125]}
   );
   gpc1_1 gpc3390 (
      {stage1_29[226]},
      {stage2_29[126]}
   );
   gpc1_1 gpc3391 (
      {stage1_29[227]},
      {stage2_29[127]}
   );
   gpc1_1 gpc3392 (
      {stage1_29[228]},
      {stage2_29[128]}
   );
   gpc1_1 gpc3393 (
      {stage1_29[229]},
      {stage2_29[129]}
   );
   gpc1_1 gpc3394 (
      {stage1_29[230]},
      {stage2_29[130]}
   );
   gpc1_1 gpc3395 (
      {stage1_29[231]},
      {stage2_29[131]}
   );
   gpc1_1 gpc3396 (
      {stage1_29[232]},
      {stage2_29[132]}
   );
   gpc1_1 gpc3397 (
      {stage1_29[233]},
      {stage2_29[133]}
   );
   gpc1_1 gpc3398 (
      {stage1_29[234]},
      {stage2_29[134]}
   );
   gpc1_1 gpc3399 (
      {stage1_29[235]},
      {stage2_29[135]}
   );
   gpc1_1 gpc3400 (
      {stage1_29[236]},
      {stage2_29[136]}
   );
   gpc1_1 gpc3401 (
      {stage1_29[237]},
      {stage2_29[137]}
   );
   gpc1_1 gpc3402 (
      {stage1_29[238]},
      {stage2_29[138]}
   );
   gpc1_1 gpc3403 (
      {stage1_29[239]},
      {stage2_29[139]}
   );
   gpc1_1 gpc3404 (
      {stage1_29[240]},
      {stage2_29[140]}
   );
   gpc1_1 gpc3405 (
      {stage1_29[241]},
      {stage2_29[141]}
   );
   gpc1_1 gpc3406 (
      {stage1_29[242]},
      {stage2_29[142]}
   );
   gpc1_1 gpc3407 (
      {stage1_30[192]},
      {stage2_30[77]}
   );
   gpc1_1 gpc3408 (
      {stage1_30[193]},
      {stage2_30[78]}
   );
   gpc1_1 gpc3409 (
      {stage1_30[194]},
      {stage2_30[79]}
   );
   gpc1_1 gpc3410 (
      {stage1_30[195]},
      {stage2_30[80]}
   );
   gpc1_1 gpc3411 (
      {stage1_30[196]},
      {stage2_30[81]}
   );
   gpc1_1 gpc3412 (
      {stage1_30[197]},
      {stage2_30[82]}
   );
   gpc1_1 gpc3413 (
      {stage1_30[198]},
      {stage2_30[83]}
   );
   gpc1_1 gpc3414 (
      {stage1_30[199]},
      {stage2_30[84]}
   );
   gpc1_1 gpc3415 (
      {stage1_30[200]},
      {stage2_30[85]}
   );
   gpc1_1 gpc3416 (
      {stage1_30[201]},
      {stage2_30[86]}
   );
   gpc1_1 gpc3417 (
      {stage1_30[202]},
      {stage2_30[87]}
   );
   gpc1_1 gpc3418 (
      {stage1_30[203]},
      {stage2_30[88]}
   );
   gpc1_1 gpc3419 (
      {stage1_30[204]},
      {stage2_30[89]}
   );
   gpc1_1 gpc3420 (
      {stage1_30[205]},
      {stage2_30[90]}
   );
   gpc1_1 gpc3421 (
      {stage1_30[206]},
      {stage2_30[91]}
   );
   gpc1_1 gpc3422 (
      {stage1_31[215]},
      {stage2_31[74]}
   );
   gpc1_1 gpc3423 (
      {stage1_31[216]},
      {stage2_31[75]}
   );
   gpc1_1 gpc3424 (
      {stage1_31[217]},
      {stage2_31[76]}
   );
   gpc1_1 gpc3425 (
      {stage1_31[218]},
      {stage2_31[77]}
   );
   gpc1_1 gpc3426 (
      {stage1_31[219]},
      {stage2_31[78]}
   );
   gpc1_1 gpc3427 (
      {stage1_31[220]},
      {stage2_31[79]}
   );
   gpc1_1 gpc3428 (
      {stage1_31[221]},
      {stage2_31[80]}
   );
   gpc1_1 gpc3429 (
      {stage1_31[222]},
      {stage2_31[81]}
   );
   gpc1_1 gpc3430 (
      {stage1_31[223]},
      {stage2_31[82]}
   );
   gpc1_1 gpc3431 (
      {stage1_31[224]},
      {stage2_31[83]}
   );
   gpc1_1 gpc3432 (
      {stage1_31[225]},
      {stage2_31[84]}
   );
   gpc1_1 gpc3433 (
      {stage1_31[226]},
      {stage2_31[85]}
   );
   gpc1_1 gpc3434 (
      {stage1_31[227]},
      {stage2_31[86]}
   );
   gpc1_1 gpc3435 (
      {stage1_31[228]},
      {stage2_31[87]}
   );
   gpc1_1 gpc3436 (
      {stage1_31[229]},
      {stage2_31[88]}
   );
   gpc1_1 gpc3437 (
      {stage1_31[230]},
      {stage2_31[89]}
   );
   gpc1_1 gpc3438 (
      {stage1_31[231]},
      {stage2_31[90]}
   );
   gpc1_1 gpc3439 (
      {stage1_31[232]},
      {stage2_31[91]}
   );
   gpc1_1 gpc3440 (
      {stage1_31[233]},
      {stage2_31[92]}
   );
   gpc1_1 gpc3441 (
      {stage1_31[234]},
      {stage2_31[93]}
   );
   gpc1_1 gpc3442 (
      {stage1_31[235]},
      {stage2_31[94]}
   );
   gpc1_1 gpc3443 (
      {stage1_31[236]},
      {stage2_31[95]}
   );
   gpc1_1 gpc3444 (
      {stage1_31[237]},
      {stage2_31[96]}
   );
   gpc1_1 gpc3445 (
      {stage1_31[238]},
      {stage2_31[97]}
   );
   gpc1_1 gpc3446 (
      {stage1_31[239]},
      {stage2_31[98]}
   );
   gpc1_1 gpc3447 (
      {stage1_31[240]},
      {stage2_31[99]}
   );
   gpc1_1 gpc3448 (
      {stage1_31[241]},
      {stage2_31[100]}
   );
   gpc1_1 gpc3449 (
      {stage1_31[242]},
      {stage2_31[101]}
   );
   gpc1_1 gpc3450 (
      {stage1_32[145]},
      {stage2_32[69]}
   );
   gpc1_1 gpc3451 (
      {stage1_32[146]},
      {stage2_32[70]}
   );
   gpc1_1 gpc3452 (
      {stage1_32[147]},
      {stage2_32[71]}
   );
   gpc1_1 gpc3453 (
      {stage1_32[148]},
      {stage2_32[72]}
   );
   gpc1_1 gpc3454 (
      {stage1_32[149]},
      {stage2_32[73]}
   );
   gpc1163_5 gpc3455 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc3456 (
      {stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc3457 (
      {stage2_0[9], stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc606_5 gpc3458 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc3459 (
      {stage2_0[21], stage2_0[22], stage2_0[23], stage2_0[24], stage2_0[25], stage2_0[26]},
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc3460 (
      {stage2_0[27], stage2_0[28], stage2_0[29], stage2_0[30], stage2_0[31], stage2_0[32]},
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc3461 (
      {stage2_0[33], stage2_0[34], stage2_0[35], stage2_0[36], stage2_0[37], stage2_0[38]},
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34], stage2_2[35], stage2_2[36]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc606_5 gpc3462 (
      {stage2_0[39], stage2_0[40], stage2_0[41], stage2_0[42], stage2_0[43], stage2_0[44]},
      {stage2_2[37], stage2_2[38], stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42]},
      {stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7],stage3_0[7]}
   );
   gpc606_5 gpc3463 (
      {stage2_0[45], stage2_0[46], stage2_0[47], stage2_0[48], stage2_0[49], stage2_0[50]},
      {stage2_2[43], stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8],stage3_0[8]}
   );
   gpc606_5 gpc3464 (
      {stage2_0[51], stage2_0[52], stage2_0[53], stage2_0[54], stage2_0[55], stage2_0[56]},
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54]},
      {stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9],stage3_0[9]}
   );
   gpc606_5 gpc3465 (
      {stage2_0[57], stage2_0[58], stage2_0[59], stage2_0[60], stage2_0[61], stage2_0[62]},
      {stage2_2[55], stage2_2[56], stage2_2[57], stage2_2[58], stage2_2[59], stage2_2[60]},
      {stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10],stage3_0[10]}
   );
   gpc606_5 gpc3466 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc3467 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[12],stage3_3[12],stage3_2[12],stage3_1[12]}
   );
   gpc606_5 gpc3468 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[13],stage3_3[13],stage3_2[13],stage3_1[13]}
   );
   gpc606_5 gpc3469 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[3],stage3_4[14],stage3_3[14],stage3_2[14],stage3_1[14]}
   );
   gpc606_5 gpc3470 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[4],stage3_4[15],stage3_3[15],stage3_2[15],stage3_1[15]}
   );
   gpc606_5 gpc3471 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[5],stage3_4[16],stage3_3[16],stage3_2[16],stage3_1[16]}
   );
   gpc606_5 gpc3472 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41], stage2_3[42]},
      {stage3_5[6],stage3_4[17],stage3_3[17],stage3_2[17],stage3_1[17]}
   );
   gpc615_5 gpc3473 (
      {stage2_2[61], stage2_2[62], stage2_2[63], stage2_2[64], stage2_2[65]},
      {stage2_3[43]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[7],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc615_5 gpc3474 (
      {stage2_2[66], stage2_2[67], stage2_2[68], stage2_2[69], stage2_2[70]},
      {stage2_3[44]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[8],stage3_4[19],stage3_3[19],stage3_2[19]}
   );
   gpc615_5 gpc3475 (
      {stage2_2[71], stage2_2[72], stage2_2[73], stage2_2[74], stage2_2[75]},
      {stage2_3[45]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[9],stage3_4[20],stage3_3[20],stage3_2[20]}
   );
   gpc615_5 gpc3476 (
      {stage2_2[76], stage2_2[77], stage2_2[78], stage2_2[79], stage2_2[80]},
      {stage2_3[46]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[10],stage3_4[21],stage3_3[21],stage3_2[21]}
   );
   gpc615_5 gpc3477 (
      {stage2_3[47], stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51]},
      {stage2_4[24]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[4],stage3_5[11],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc3478 (
      {stage2_3[52], stage2_3[53], stage2_3[54], stage2_3[55], stage2_3[56]},
      {stage2_4[25]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[5],stage3_5[12],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc3479 (
      {stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61]},
      {stage2_4[26]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[6],stage3_5[13],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc3480 (
      {stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66]},
      {stage2_4[27]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[7],stage3_5[14],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc3481 (
      {stage2_3[67], stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71]},
      {stage2_4[28]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[8],stage3_5[15],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc3482 (
      {stage2_3[72], stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76]},
      {stage2_4[29]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[9],stage3_5[16],stage3_4[27],stage3_3[27]}
   );
   gpc606_5 gpc3483 (
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[6],stage3_6[10],stage3_5[17],stage3_4[28]}
   );
   gpc606_5 gpc3484 (
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[7],stage3_6[11],stage3_5[18],stage3_4[29]}
   );
   gpc606_5 gpc3485 (
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46], stage2_4[47]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[8],stage3_6[12],stage3_5[19],stage3_4[30]}
   );
   gpc606_5 gpc3486 (
      {stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51], stage2_4[52], stage2_4[53]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[9],stage3_6[13],stage3_5[20],stage3_4[31]}
   );
   gpc606_5 gpc3487 (
      {stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58], stage2_4[59]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[10],stage3_6[14],stage3_5[21],stage3_4[32]}
   );
   gpc606_5 gpc3488 (
      {stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[11],stage3_6[15],stage3_5[22],stage3_4[33]}
   );
   gpc606_5 gpc3489 (
      {stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[12],stage3_6[16],stage3_5[23],stage3_4[34]}
   );
   gpc606_5 gpc3490 (
      {stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76], stage2_4[77]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[13],stage3_6[17],stage3_5[24],stage3_4[35]}
   );
   gpc606_5 gpc3491 (
      {stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82], stage2_4[83]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[14],stage3_6[18],stage3_5[25],stage3_4[36]}
   );
   gpc606_5 gpc3492 (
      {stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88], stage2_4[89]},
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58], stage2_6[59]},
      {stage3_8[9],stage3_7[15],stage3_6[19],stage3_5[26],stage3_4[37]}
   );
   gpc606_5 gpc3493 (
      {stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94], stage2_4[95]},
      {stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63], stage2_6[64], stage2_6[65]},
      {stage3_8[10],stage3_7[16],stage3_6[20],stage3_5[27],stage3_4[38]}
   );
   gpc606_5 gpc3494 (
      {stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100], stage2_4[101]},
      {stage2_6[66], stage2_6[67], stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71]},
      {stage3_8[11],stage3_7[17],stage3_6[21],stage3_5[28],stage3_4[39]}
   );
   gpc606_5 gpc3495 (
      {stage2_4[102], stage2_4[103], stage2_4[104], stage2_4[105], stage2_4[106], stage2_4[107]},
      {stage2_6[72], stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage3_8[12],stage3_7[18],stage3_6[22],stage3_5[29],stage3_4[40]}
   );
   gpc606_5 gpc3496 (
      {stage2_4[108], stage2_4[109], stage2_4[110], stage2_4[111], stage2_4[112], stage2_4[113]},
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83]},
      {stage3_8[13],stage3_7[19],stage3_6[23],stage3_5[30],stage3_4[41]}
   );
   gpc606_5 gpc3497 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[14],stage3_7[20],stage3_6[24],stage3_5[31]}
   );
   gpc606_5 gpc3498 (
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[15],stage3_7[21],stage3_6[25],stage3_5[32]}
   );
   gpc606_5 gpc3499 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[16],stage3_7[22],stage3_6[26],stage3_5[33]}
   );
   gpc606_5 gpc3500 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[17],stage3_7[23],stage3_6[27],stage3_5[34]}
   );
   gpc606_5 gpc3501 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[18],stage3_7[24],stage3_6[28],stage3_5[35]}
   );
   gpc606_5 gpc3502 (
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[19],stage3_7[25],stage3_6[29],stage3_5[36]}
   );
   gpc615_5 gpc3503 (
      {stage2_6[84], stage2_6[85], stage2_6[86], stage2_6[87], stage2_6[88]},
      {stage2_7[36]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[6],stage3_8[20],stage3_7[26],stage3_6[30]}
   );
   gpc615_5 gpc3504 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[7],stage3_8[21],stage3_7[27]}
   );
   gpc615_5 gpc3505 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[8],stage3_8[22],stage3_7[28]}
   );
   gpc615_5 gpc3506 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[9],stage3_8[23],stage3_7[29]}
   );
   gpc615_5 gpc3507 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[10],stage3_8[24],stage3_7[30]}
   );
   gpc615_5 gpc3508 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61]},
      {stage2_8[10]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[5],stage3_9[11],stage3_8[25],stage3_7[31]}
   );
   gpc615_5 gpc3509 (
      {stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66]},
      {stage2_8[11]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[6],stage3_9[12],stage3_8[26],stage3_7[32]}
   );
   gpc615_5 gpc3510 (
      {stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage2_8[12]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[7],stage3_9[13],stage3_8[27],stage3_7[33]}
   );
   gpc615_5 gpc3511 (
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76]},
      {stage2_8[13]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[8],stage3_9[14],stage3_8[28],stage3_7[34]}
   );
   gpc615_5 gpc3512 (
      {stage2_7[77], stage2_7[78], stage2_7[79], stage2_7[80], stage2_7[81]},
      {stage2_8[14]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[9],stage3_9[15],stage3_8[29],stage3_7[35]}
   );
   gpc615_5 gpc3513 (
      {stage2_7[82], stage2_7[83], stage2_7[84], stage2_7[85], stage2_7[86]},
      {stage2_8[15]},
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage3_11[9],stage3_10[10],stage3_9[16],stage3_8[30],stage3_7[36]}
   );
   gpc615_5 gpc3514 (
      {stage2_7[87], stage2_7[88], stage2_7[89], stage2_7[90], stage2_7[91]},
      {stage2_8[16]},
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage3_11[10],stage3_10[11],stage3_9[17],stage3_8[31],stage3_7[37]}
   );
   gpc615_5 gpc3515 (
      {stage2_7[92], stage2_7[93], stage2_7[94], stage2_7[95], stage2_7[96]},
      {stage2_8[17]},
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage3_11[11],stage3_10[12],stage3_9[18],stage3_8[32],stage3_7[38]}
   );
   gpc615_5 gpc3516 (
      {stage2_7[97], stage2_7[98], stage2_7[99], stage2_7[100], stage2_7[101]},
      {stage2_8[18]},
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage3_11[12],stage3_10[13],stage3_9[19],stage3_8[33],stage3_7[39]}
   );
   gpc606_5 gpc3517 (
      {stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[13],stage3_10[14],stage3_9[20],stage3_8[34]}
   );
   gpc606_5 gpc3518 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[14],stage3_10[15],stage3_9[21],stage3_8[35]}
   );
   gpc606_5 gpc3519 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[15],stage3_10[16],stage3_9[22],stage3_8[36]}
   );
   gpc606_5 gpc3520 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[16],stage3_10[17],stage3_9[23],stage3_8[37]}
   );
   gpc615_5 gpc3521 (
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82]},
      {stage2_10[24]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[4],stage3_11[17],stage3_10[18],stage3_9[24]}
   );
   gpc606_5 gpc3522 (
      {stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[5],stage3_11[18],stage3_10[19]}
   );
   gpc606_5 gpc3523 (
      {stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[6],stage3_11[19],stage3_10[20]}
   );
   gpc606_5 gpc3524 (
      {stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[7],stage3_11[20],stage3_10[21]}
   );
   gpc606_5 gpc3525 (
      {stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[4],stage3_12[8],stage3_11[21],stage3_10[22]}
   );
   gpc606_5 gpc3526 (
      {stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[5],stage3_12[9],stage3_11[22],stage3_10[23]}
   );
   gpc606_5 gpc3527 (
      {stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[6],stage3_12[10],stage3_11[23],stage3_10[24]}
   );
   gpc606_5 gpc3528 (
      {stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[7],stage3_12[11],stage3_11[24],stage3_10[25]}
   );
   gpc615_5 gpc3529 (
      {stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage2_11[6]},
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage3_14[7],stage3_13[8],stage3_12[12],stage3_11[25],stage3_10[26]}
   );
   gpc615_5 gpc3530 (
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76]},
      {stage2_11[7]},
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage3_14[8],stage3_13[9],stage3_12[13],stage3_11[26],stage3_10[27]}
   );
   gpc615_5 gpc3531 (
      {stage2_10[77], stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81]},
      {stage2_11[8]},
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage3_14[9],stage3_13[10],stage3_12[14],stage3_11[27],stage3_10[28]}
   );
   gpc615_5 gpc3532 (
      {stage2_10[82], stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86]},
      {stage2_11[9]},
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage3_14[10],stage3_13[11],stage3_12[15],stage3_11[28],stage3_10[29]}
   );
   gpc615_5 gpc3533 (
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[66]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[11],stage3_13[12],stage3_12[16],stage3_11[29]}
   );
   gpc615_5 gpc3534 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_12[67]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[12],stage3_13[13],stage3_12[17],stage3_11[30]}
   );
   gpc615_5 gpc3535 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_12[68]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[13],stage3_13[14],stage3_12[18],stage3_11[31]}
   );
   gpc615_5 gpc3536 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_12[69]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[14],stage3_13[15],stage3_12[19],stage3_11[32]}
   );
   gpc615_5 gpc3537 (
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34]},
      {stage2_12[70]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[15],stage3_13[16],stage3_12[20],stage3_11[33]}
   );
   gpc615_5 gpc3538 (
      {stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage2_12[71]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[16],stage3_13[17],stage3_12[21],stage3_11[34]}
   );
   gpc615_5 gpc3539 (
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_12[72]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[17],stage3_13[18],stage3_12[22],stage3_11[35]}
   );
   gpc615_5 gpc3540 (
      {stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49]},
      {stage2_12[73]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[18],stage3_13[19],stage3_12[23],stage3_11[36]}
   );
   gpc615_5 gpc3541 (
      {stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54]},
      {stage2_12[74]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[19],stage3_13[20],stage3_12[24],stage3_11[37]}
   );
   gpc615_5 gpc3542 (
      {stage2_11[55], stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59]},
      {stage2_12[75]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[20],stage3_13[21],stage3_12[25],stage3_11[38]}
   );
   gpc615_5 gpc3543 (
      {stage2_11[60], stage2_11[61], stage2_11[62], stage2_11[63], stage2_11[64]},
      {stage2_12[76]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[21],stage3_13[22],stage3_12[26],stage3_11[39]}
   );
   gpc615_5 gpc3544 (
      {stage2_11[65], stage2_11[66], stage2_11[67], stage2_11[68], stage2_11[69]},
      {stage2_12[77]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[22],stage3_13[23],stage3_12[27],stage3_11[40]}
   );
   gpc615_5 gpc3545 (
      {stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73], stage2_11[74]},
      {stage2_12[78]},
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage3_15[12],stage3_14[23],stage3_13[24],stage3_12[28],stage3_11[41]}
   );
   gpc615_5 gpc3546 (
      {stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79]},
      {stage2_12[79]},
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage3_15[13],stage3_14[24],stage3_13[25],stage3_12[29],stage3_11[42]}
   );
   gpc615_5 gpc3547 (
      {stage2_11[80], stage2_11[81], stage2_11[82], stage2_11[83], stage2_11[84]},
      {stage2_12[80]},
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage3_15[14],stage3_14[25],stage3_13[26],stage3_12[30],stage3_11[43]}
   );
   gpc615_5 gpc3548 (
      {stage2_11[85], stage2_11[86], stage2_11[87], stage2_11[88], stage2_11[89]},
      {stage2_12[81]},
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94], stage2_13[95]},
      {stage3_15[15],stage3_14[26],stage3_13[27],stage3_12[31],stage3_11[44]}
   );
   gpc615_5 gpc3549 (
      {stage2_11[90], stage2_11[91], stage2_11[92], stage2_11[93], stage2_11[94]},
      {stage2_12[82]},
      {stage2_13[96], stage2_13[97], stage2_13[98], stage2_13[99], stage2_13[100], stage2_13[101]},
      {stage3_15[16],stage3_14[27],stage3_13[28],stage3_12[32],stage3_11[45]}
   );
   gpc615_5 gpc3550 (
      {stage2_11[95], stage2_11[96], stage2_11[97], stage2_11[98], stage2_11[99]},
      {stage2_12[83]},
      {stage2_13[102], stage2_13[103], stage2_13[104], stage2_13[105], stage2_13[106], stage2_13[107]},
      {stage3_15[17],stage3_14[28],stage3_13[29],stage3_12[33],stage3_11[46]}
   );
   gpc615_5 gpc3551 (
      {stage2_11[100], stage2_11[101], stage2_11[102], stage2_11[103], stage2_11[104]},
      {stage2_12[84]},
      {stage2_13[108], stage2_13[109], stage2_13[110], stage2_13[111], stage2_13[112], stage2_13[113]},
      {stage3_15[18],stage3_14[29],stage3_13[30],stage3_12[34],stage3_11[47]}
   );
   gpc615_5 gpc3552 (
      {stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108], stage2_11[109]},
      {stage2_12[85]},
      {stage2_13[114], stage2_13[115], stage2_13[116], stage2_13[117], stage2_13[118], stage2_13[119]},
      {stage3_15[19],stage3_14[30],stage3_13[31],stage3_12[35],stage3_11[48]}
   );
   gpc606_5 gpc3553 (
      {stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89], stage2_12[90], stage2_12[91]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[20],stage3_14[31],stage3_13[32],stage3_12[36]}
   );
   gpc615_5 gpc3554 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[21],stage3_14[32]}
   );
   gpc615_5 gpc3555 (
      {stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[22],stage3_14[33]}
   );
   gpc615_5 gpc3556 (
      {stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[23],stage3_14[34]}
   );
   gpc615_5 gpc3557 (
      {stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[4],stage3_15[24],stage3_14[35]}
   );
   gpc615_5 gpc3558 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30]},
      {stage2_15[4]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[4],stage3_16[5],stage3_15[25],stage3_14[36]}
   );
   gpc615_5 gpc3559 (
      {stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_15[5]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[5],stage3_16[6],stage3_15[26],stage3_14[37]}
   );
   gpc615_5 gpc3560 (
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40]},
      {stage2_15[6]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[6],stage3_16[7],stage3_15[27],stage3_14[38]}
   );
   gpc615_5 gpc3561 (
      {stage2_14[41], stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45]},
      {stage2_15[7]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[7],stage3_16[8],stage3_15[28],stage3_14[39]}
   );
   gpc615_5 gpc3562 (
      {stage2_14[46], stage2_14[47], stage2_14[48], stage2_14[49], stage2_14[50]},
      {stage2_15[8]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[8],stage3_16[9],stage3_15[29],stage3_14[40]}
   );
   gpc615_5 gpc3563 (
      {stage2_14[51], stage2_14[52], stage2_14[53], stage2_14[54], stage2_14[55]},
      {stage2_15[9]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[9],stage3_16[10],stage3_15[30],stage3_14[41]}
   );
   gpc615_5 gpc3564 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[60]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[10],stage3_17[10],stage3_16[11],stage3_15[31]}
   );
   gpc615_5 gpc3565 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[61]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[11],stage3_17[11],stage3_16[12],stage3_15[32]}
   );
   gpc615_5 gpc3566 (
      {stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23], stage2_15[24]},
      {stage2_16[62]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[12],stage3_17[12],stage3_16[13],stage3_15[33]}
   );
   gpc615_5 gpc3567 (
      {stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage2_16[63]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[13],stage3_17[13],stage3_16[14],stage3_15[34]}
   );
   gpc615_5 gpc3568 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[64]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[14],stage3_17[14],stage3_16[15],stage3_15[35]}
   );
   gpc615_5 gpc3569 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[65]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[15],stage3_17[15],stage3_16[16],stage3_15[36]}
   );
   gpc615_5 gpc3570 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[66]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[16],stage3_17[16],stage3_16[17],stage3_15[37]}
   );
   gpc615_5 gpc3571 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[67]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[17],stage3_17[17],stage3_16[18],stage3_15[38]}
   );
   gpc615_5 gpc3572 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[68]},
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage3_19[8],stage3_18[18],stage3_17[18],stage3_16[19],stage3_15[39]}
   );
   gpc615_5 gpc3573 (
      {stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59]},
      {stage2_16[69]},
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage3_19[9],stage3_18[19],stage3_17[19],stage3_16[20],stage3_15[40]}
   );
   gpc615_5 gpc3574 (
      {stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_16[70]},
      {stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65]},
      {stage3_19[10],stage3_18[20],stage3_17[20],stage3_16[21],stage3_15[41]}
   );
   gpc615_5 gpc3575 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69]},
      {stage2_16[71]},
      {stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71]},
      {stage3_19[11],stage3_18[21],stage3_17[21],stage3_16[22],stage3_15[42]}
   );
   gpc135_4 gpc3576 (
      {stage2_16[72], stage2_16[73], stage2_16[74], stage2_16[75], stage2_16[76]},
      {stage2_17[72], stage2_17[73], stage2_17[74]},
      {stage2_18[0]},
      {stage3_19[12],stage3_18[22],stage3_17[22],stage3_16[23]}
   );
   gpc606_5 gpc3577 (
      {stage2_16[77], stage2_16[78], stage2_16[79], stage2_16[80], stage2_16[81], stage2_16[82]},
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[0],stage3_19[13],stage3_18[23],stage3_17[23],stage3_16[24]}
   );
   gpc606_5 gpc3578 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[14],stage3_18[24]}
   );
   gpc606_5 gpc3579 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[15],stage3_18[25]}
   );
   gpc606_5 gpc3580 (
      {stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[3],stage3_19[16],stage3_18[26]}
   );
   gpc606_5 gpc3581 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[4],stage3_19[17],stage3_18[27]}
   );
   gpc606_5 gpc3582 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35], stage2_18[36]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[5],stage3_19[18],stage3_18[28]}
   );
   gpc606_5 gpc3583 (
      {stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40], stage2_18[41], stage2_18[42]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[6],stage3_19[19],stage3_18[29]}
   );
   gpc606_5 gpc3584 (
      {stage2_18[43], stage2_18[44], stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[7],stage3_19[20],stage3_18[30]}
   );
   gpc606_5 gpc3585 (
      {stage2_18[49], stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[7],stage3_20[8],stage3_19[21],stage3_18[31]}
   );
   gpc606_5 gpc3586 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[8],stage3_20[9],stage3_19[22],stage3_18[32]}
   );
   gpc606_5 gpc3587 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65], stage2_18[66]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[9],stage3_20[10],stage3_19[23],stage3_18[33]}
   );
   gpc606_5 gpc3588 (
      {stage2_18[67], stage2_18[68], stage2_18[69], stage2_18[70], stage2_18[71], stage2_18[72]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[10],stage3_20[11],stage3_19[24],stage3_18[34]}
   );
   gpc606_5 gpc3589 (
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[11],stage3_21[11],stage3_20[12],stage3_19[25]}
   );
   gpc606_5 gpc3590 (
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[12],stage3_21[12],stage3_20[13],stage3_19[26]}
   );
   gpc606_5 gpc3591 (
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage3_23[2],stage3_22[13],stage3_21[13],stage3_20[14],stage3_19[27]}
   );
   gpc606_5 gpc3592 (
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage3_23[3],stage3_22[14],stage3_21[14],stage3_20[15],stage3_19[28]}
   );
   gpc606_5 gpc3593 (
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage3_23[4],stage3_22[15],stage3_21[15],stage3_20[16],stage3_19[29]}
   );
   gpc606_5 gpc3594 (
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34], stage2_21[35]},
      {stage3_23[5],stage3_22[16],stage3_21[16],stage3_20[17],stage3_19[30]}
   );
   gpc606_5 gpc3595 (
      {stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39], stage2_21[40], stage2_21[41]},
      {stage3_23[6],stage3_22[17],stage3_21[17],stage3_20[18],stage3_19[31]}
   );
   gpc606_5 gpc3596 (
      {stage2_19[42], stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47]},
      {stage3_23[7],stage3_22[18],stage3_21[18],stage3_20[19],stage3_19[32]}
   );
   gpc606_5 gpc3597 (
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51], stage2_21[52], stage2_21[53]},
      {stage3_23[8],stage3_22[19],stage3_21[19],stage3_20[20],stage3_19[33]}
   );
   gpc615_5 gpc3598 (
      {stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57], stage2_19[58]},
      {stage2_20[66]},
      {stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57], stage2_21[58], stage2_21[59]},
      {stage3_23[9],stage3_22[20],stage3_21[20],stage3_20[21],stage3_19[34]}
   );
   gpc615_5 gpc3599 (
      {stage2_19[59], stage2_19[60], stage2_19[61], stage2_19[62], stage2_19[63]},
      {stage2_20[67]},
      {stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63], stage2_21[64], stage2_21[65]},
      {stage3_23[10],stage3_22[21],stage3_21[21],stage3_20[22],stage3_19[35]}
   );
   gpc606_5 gpc3600 (
      {stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71], stage2_20[72], stage2_20[73]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[11],stage3_22[22],stage3_21[22],stage3_20[23]}
   );
   gpc606_5 gpc3601 (
      {stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77], stage2_20[78], stage2_20[79]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[12],stage3_22[23],stage3_21[23],stage3_20[24]}
   );
   gpc606_5 gpc3602 (
      {stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83], stage2_20[84], stage2_20[85]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[13],stage3_22[24],stage3_21[24],stage3_20[25]}
   );
   gpc606_5 gpc3603 (
      {stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89], stage2_20[90], stage2_20[91]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[14],stage3_22[25],stage3_21[25],stage3_20[26]}
   );
   gpc606_5 gpc3604 (
      {stage2_20[92], stage2_20[93], stage2_20[94], stage2_20[95], stage2_20[96], stage2_20[97]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[15],stage3_22[26],stage3_21[26],stage3_20[27]}
   );
   gpc606_5 gpc3605 (
      {stage2_20[98], stage2_20[99], stage2_20[100], stage2_20[101], stage2_20[102], stage2_20[103]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage3_24[5],stage3_23[16],stage3_22[27],stage3_21[27],stage3_20[28]}
   );
   gpc606_5 gpc3606 (
      {stage2_20[104], stage2_20[105], stage2_20[106], stage2_20[107], stage2_20[108], stage2_20[109]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage3_24[6],stage3_23[17],stage3_22[28],stage3_21[28],stage3_20[29]}
   );
   gpc606_5 gpc3607 (
      {stage2_21[66], stage2_21[67], stage2_21[68], stage2_21[69], stage2_21[70], stage2_21[71]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[7],stage3_23[18],stage3_22[29],stage3_21[29]}
   );
   gpc606_5 gpc3608 (
      {stage2_21[72], stage2_21[73], stage2_21[74], stage2_21[75], stage2_21[76], stage2_21[77]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[8],stage3_23[19],stage3_22[30],stage3_21[30]}
   );
   gpc606_5 gpc3609 (
      {stage2_21[78], stage2_21[79], stage2_21[80], stage2_21[81], stage2_21[82], stage2_21[83]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[9],stage3_23[20],stage3_22[31],stage3_21[31]}
   );
   gpc606_5 gpc3610 (
      {stage2_21[84], stage2_21[85], stage2_21[86], stage2_21[87], stage2_21[88], stage2_21[89]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[10],stage3_23[21],stage3_22[32],stage3_21[32]}
   );
   gpc606_5 gpc3611 (
      {stage2_21[90], stage2_21[91], stage2_21[92], stage2_21[93], stage2_21[94], stage2_21[95]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[11],stage3_23[22],stage3_22[33],stage3_21[33]}
   );
   gpc615_5 gpc3612 (
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46]},
      {stage2_23[30]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[5],stage3_24[12],stage3_23[23],stage3_22[34]}
   );
   gpc615_5 gpc3613 (
      {stage2_22[47], stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51]},
      {stage2_23[31]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[6],stage3_24[13],stage3_23[24],stage3_22[35]}
   );
   gpc615_5 gpc3614 (
      {stage2_22[52], stage2_22[53], stage2_22[54], stage2_22[55], stage2_22[56]},
      {stage2_23[32]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[7],stage3_24[14],stage3_23[25],stage3_22[36]}
   );
   gpc615_5 gpc3615 (
      {stage2_22[57], stage2_22[58], stage2_22[59], stage2_22[60], stage2_22[61]},
      {stage2_23[33]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[8],stage3_24[15],stage3_23[26],stage3_22[37]}
   );
   gpc615_5 gpc3616 (
      {stage2_22[62], stage2_22[63], stage2_22[64], stage2_22[65], stage2_22[66]},
      {stage2_23[34]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[9],stage3_24[16],stage3_23[27],stage3_22[38]}
   );
   gpc615_5 gpc3617 (
      {stage2_22[67], stage2_22[68], stage2_22[69], stage2_22[70], stage2_22[71]},
      {stage2_23[35]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[10],stage3_24[17],stage3_23[28],stage3_22[39]}
   );
   gpc615_5 gpc3618 (
      {stage2_22[72], stage2_22[73], stage2_22[74], stage2_22[75], stage2_22[76]},
      {stage2_23[36]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[11],stage3_24[18],stage3_23[29],stage3_22[40]}
   );
   gpc615_5 gpc3619 (
      {stage2_22[77], stage2_22[78], stage2_22[79], stage2_22[80], stage2_22[81]},
      {stage2_23[37]},
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage3_26[7],stage3_25[12],stage3_24[19],stage3_23[30],stage3_22[41]}
   );
   gpc615_5 gpc3620 (
      {stage2_22[82], stage2_22[83], stage2_22[84], stage2_22[85], stage2_22[86]},
      {stage2_23[38]},
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage3_26[8],stage3_25[13],stage3_24[20],stage3_23[31],stage3_22[42]}
   );
   gpc606_5 gpc3621 (
      {stage2_23[39], stage2_23[40], stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[9],stage3_25[14],stage3_24[21],stage3_23[32]}
   );
   gpc606_5 gpc3622 (
      {stage2_23[45], stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[10],stage3_25[15],stage3_24[22],stage3_23[33]}
   );
   gpc606_5 gpc3623 (
      {stage2_23[51], stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55], stage2_23[56]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[11],stage3_25[16],stage3_24[23],stage3_23[34]}
   );
   gpc606_5 gpc3624 (
      {stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60], stage2_23[61], stage2_23[62]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[12],stage3_25[17],stage3_24[24],stage3_23[35]}
   );
   gpc606_5 gpc3625 (
      {stage2_23[63], stage2_23[64], stage2_23[65], stage2_23[66], stage2_23[67], stage2_23[68]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[13],stage3_25[18],stage3_24[25],stage3_23[36]}
   );
   gpc606_5 gpc3626 (
      {stage2_23[69], stage2_23[70], stage2_23[71], stage2_23[72], stage2_23[73], stage2_23[74]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[14],stage3_25[19],stage3_24[26],stage3_23[37]}
   );
   gpc606_5 gpc3627 (
      {stage2_23[75], stage2_23[76], stage2_23[77], stage2_23[78], stage2_23[79], stage2_23[80]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[15],stage3_25[20],stage3_24[27],stage3_23[38]}
   );
   gpc606_5 gpc3628 (
      {stage2_23[81], stage2_23[82], stage2_23[83], stage2_23[84], stage2_23[85], stage2_23[86]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[16],stage3_25[21],stage3_24[28],stage3_23[39]}
   );
   gpc606_5 gpc3629 (
      {stage2_23[87], stage2_23[88], stage2_23[89], stage2_23[90], stage2_23[91], stage2_23[92]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[17],stage3_25[22],stage3_24[29],stage3_23[40]}
   );
   gpc606_5 gpc3630 (
      {stage2_23[93], stage2_23[94], stage2_23[95], stage2_23[96], stage2_23[97], stage2_23[98]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[18],stage3_25[23],stage3_24[30],stage3_23[41]}
   );
   gpc606_5 gpc3631 (
      {stage2_23[99], stage2_23[100], stage2_23[101], stage2_23[102], stage2_23[103], stage2_23[104]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[19],stage3_25[24],stage3_24[31],stage3_23[42]}
   );
   gpc606_5 gpc3632 (
      {stage2_23[105], stage2_23[106], stage2_23[107], stage2_23[108], stage2_23[109], stage2_23[110]},
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage3_27[11],stage3_26[20],stage3_25[25],stage3_24[32],stage3_23[43]}
   );
   gpc606_5 gpc3633 (
      {stage2_23[111], stage2_23[112], stage2_23[113], stage2_23[114], stage2_23[115], stage2_23[116]},
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage3_27[12],stage3_26[21],stage3_25[26],stage3_24[33],stage3_23[44]}
   );
   gpc606_5 gpc3634 (
      {stage2_23[117], stage2_23[118], stage2_23[119], stage2_23[120], stage2_23[121], stage2_23[122]},
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage3_27[13],stage3_26[22],stage3_25[27],stage3_24[34],stage3_23[45]}
   );
   gpc606_5 gpc3635 (
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[14],stage3_26[23],stage3_25[28],stage3_24[35]}
   );
   gpc606_5 gpc3636 (
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[15],stage3_26[24],stage3_25[29],stage3_24[36]}
   );
   gpc1163_5 gpc3637 (
      {stage2_26[12], stage2_26[13], stage2_26[14]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage2_28[0]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[0],stage3_28[2],stage3_27[16],stage3_26[25]}
   );
   gpc606_5 gpc3638 (
      {stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20]},
      {stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6]},
      {stage3_30[1],stage3_29[1],stage3_28[3],stage3_27[17],stage3_26[26]}
   );
   gpc606_5 gpc3639 (
      {stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24], stage2_26[25], stage2_26[26]},
      {stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12]},
      {stage3_30[2],stage3_29[2],stage3_28[4],stage3_27[18],stage3_26[27]}
   );
   gpc606_5 gpc3640 (
      {stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18]},
      {stage3_30[3],stage3_29[3],stage3_28[5],stage3_27[19],stage3_26[28]}
   );
   gpc606_5 gpc3641 (
      {stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23], stage2_28[24]},
      {stage3_30[4],stage3_29[4],stage3_28[6],stage3_27[20],stage3_26[29]}
   );
   gpc606_5 gpc3642 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43], stage2_26[44]},
      {stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28], stage2_28[29], stage2_28[30]},
      {stage3_30[5],stage3_29[5],stage3_28[7],stage3_27[21],stage3_26[30]}
   );
   gpc606_5 gpc3643 (
      {stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48], stage2_26[49], stage2_26[50]},
      {stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35], stage2_28[36]},
      {stage3_30[6],stage3_29[6],stage3_28[8],stage3_27[22],stage3_26[31]}
   );
   gpc606_5 gpc3644 (
      {stage2_26[51], stage2_26[52], stage2_26[53], stage2_26[54], stage2_26[55], stage2_26[56]},
      {stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42]},
      {stage3_30[7],stage3_29[7],stage3_28[9],stage3_27[23],stage3_26[32]}
   );
   gpc606_5 gpc3645 (
      {stage2_26[57], stage2_26[58], stage2_26[59], stage2_26[60], stage2_26[61], stage2_26[62]},
      {stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage3_30[8],stage3_29[8],stage3_28[10],stage3_27[24],stage3_26[33]}
   );
   gpc606_5 gpc3646 (
      {stage2_26[63], stage2_26[64], stage2_26[65], stage2_26[66], stage2_26[67], stage2_26[68]},
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53], stage2_28[54]},
      {stage3_30[9],stage3_29[9],stage3_28[11],stage3_27[25],stage3_26[34]}
   );
   gpc606_5 gpc3647 (
      {stage2_26[69], stage2_26[70], stage2_26[71], stage2_26[72], stage2_26[73], stage2_26[74]},
      {stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58], stage2_28[59], stage2_28[60]},
      {stage3_30[10],stage3_29[10],stage3_28[12],stage3_27[26],stage3_26[35]}
   );
   gpc606_5 gpc3648 (
      {stage2_26[75], stage2_26[76], stage2_26[77], stage2_26[78], stage2_26[79], stage2_26[80]},
      {stage2_28[61], stage2_28[62], stage2_28[63], stage2_28[64], stage2_28[65], stage2_28[66]},
      {stage3_30[11],stage3_29[11],stage3_28[13],stage3_27[27],stage3_26[36]}
   );
   gpc606_5 gpc3649 (
      {stage2_26[81], stage2_26[82], stage2_26[83], stage2_26[84], stage2_26[85], stage2_26[86]},
      {stage2_28[67], stage2_28[68], stage2_28[69], stage2_28[70], stage2_28[71], stage2_28[72]},
      {stage3_30[12],stage3_29[12],stage3_28[14],stage3_27[28],stage3_26[37]}
   );
   gpc606_5 gpc3650 (
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6]},
      {stage3_31[0],stage3_30[13],stage3_29[13],stage3_28[15],stage3_27[29]}
   );
   gpc615_5 gpc3651 (
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16]},
      {stage2_28[73]},
      {stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11], stage2_29[12]},
      {stage3_31[1],stage3_30[14],stage3_29[14],stage3_28[16],stage3_27[30]}
   );
   gpc615_5 gpc3652 (
      {stage2_27[17], stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21]},
      {stage2_28[74]},
      {stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17], stage2_29[18]},
      {stage3_31[2],stage3_30[15],stage3_29[15],stage3_28[17],stage3_27[31]}
   );
   gpc615_5 gpc3653 (
      {stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26]},
      {stage2_28[75]},
      {stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23], stage2_29[24]},
      {stage3_31[3],stage3_30[16],stage3_29[16],stage3_28[18],stage3_27[32]}
   );
   gpc615_5 gpc3654 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31]},
      {stage2_28[76]},
      {stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29], stage2_29[30]},
      {stage3_31[4],stage3_30[17],stage3_29[17],stage3_28[19],stage3_27[33]}
   );
   gpc615_5 gpc3655 (
      {stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36]},
      {stage2_28[77]},
      {stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35], stage2_29[36]},
      {stage3_31[5],stage3_30[18],stage3_29[18],stage3_28[20],stage3_27[34]}
   );
   gpc615_5 gpc3656 (
      {stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_28[78]},
      {stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41], stage2_29[42]},
      {stage3_31[6],stage3_30[19],stage3_29[19],stage3_28[21],stage3_27[35]}
   );
   gpc615_5 gpc3657 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46]},
      {stage2_28[79]},
      {stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47], stage2_29[48]},
      {stage3_31[7],stage3_30[20],stage3_29[20],stage3_28[22],stage3_27[36]}
   );
   gpc615_5 gpc3658 (
      {stage2_27[47], stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51]},
      {stage2_28[80]},
      {stage2_29[49], stage2_29[50], stage2_29[51], stage2_29[52], stage2_29[53], stage2_29[54]},
      {stage3_31[8],stage3_30[21],stage3_29[21],stage3_28[23],stage3_27[37]}
   );
   gpc615_5 gpc3659 (
      {stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[81]},
      {stage2_29[55], stage2_29[56], stage2_29[57], stage2_29[58], stage2_29[59], stage2_29[60]},
      {stage3_31[9],stage3_30[22],stage3_29[22],stage3_28[24],stage3_27[38]}
   );
   gpc615_5 gpc3660 (
      {stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61]},
      {stage2_28[82]},
      {stage2_29[61], stage2_29[62], stage2_29[63], stage2_29[64], stage2_29[65], stage2_29[66]},
      {stage3_31[10],stage3_30[23],stage3_29[23],stage3_28[25],stage3_27[39]}
   );
   gpc615_5 gpc3661 (
      {stage2_27[62], stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66]},
      {stage2_28[83]},
      {stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70], stage2_29[71], stage2_29[72]},
      {stage3_31[11],stage3_30[24],stage3_29[24],stage3_28[26],stage3_27[40]}
   );
   gpc615_5 gpc3662 (
      {stage2_27[67], stage2_27[68], stage2_27[69], stage2_27[70], stage2_27[71]},
      {stage2_28[84]},
      {stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76], stage2_29[77], stage2_29[78]},
      {stage3_31[12],stage3_30[25],stage3_29[25],stage3_28[27],stage3_27[41]}
   );
   gpc606_5 gpc3663 (
      {stage2_28[85], stage2_28[86], stage2_28[87], stage2_28[88], stage2_28[89], stage2_28[90]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[13],stage3_30[26],stage3_29[26],stage3_28[28]}
   );
   gpc606_5 gpc3664 (
      {stage2_28[91], stage2_28[92], stage2_28[93], stage2_28[94], stage2_28[95], stage2_28[96]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[14],stage3_30[27],stage3_29[27],stage3_28[29]}
   );
   gpc606_5 gpc3665 (
      {stage2_28[97], stage2_28[98], stage2_28[99], stage2_28[100], stage2_28[101], stage2_28[102]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[15],stage3_30[28],stage3_29[28],stage3_28[30]}
   );
   gpc606_5 gpc3666 (
      {stage2_28[103], stage2_28[104], stage2_28[105], stage2_28[106], stage2_28[107], stage2_28[108]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[16],stage3_30[29],stage3_29[29],stage3_28[31]}
   );
   gpc606_5 gpc3667 (
      {stage2_28[109], stage2_28[110], stage2_28[111], stage2_28[112], stage2_28[113], stage2_28[114]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[17],stage3_30[30],stage3_29[30],stage3_28[32]}
   );
   gpc606_5 gpc3668 (
      {stage2_28[115], stage2_28[116], stage2_28[117], stage2_28[118], stage2_28[119], stage2_28[120]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[18],stage3_30[31],stage3_29[31],stage3_28[33]}
   );
   gpc606_5 gpc3669 (
      {stage2_28[121], stage2_28[122], stage2_28[123], stage2_28[124], stage2_28[125], stage2_28[126]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[19],stage3_30[32],stage3_29[32],stage3_28[34]}
   );
   gpc606_5 gpc3670 (
      {stage2_28[127], stage2_28[128], stage2_28[129], stage2_28[130], stage2_28[131], stage2_28[132]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[20],stage3_30[33],stage3_29[33],stage3_28[35]}
   );
   gpc606_5 gpc3671 (
      {stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82], stage2_29[83], stage2_29[84]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[8],stage3_31[21],stage3_30[34],stage3_29[34]}
   );
   gpc606_5 gpc3672 (
      {stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88], stage2_29[89], stage2_29[90]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[9],stage3_31[22],stage3_30[35],stage3_29[35]}
   );
   gpc606_5 gpc3673 (
      {stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94], stage2_29[95], stage2_29[96]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[10],stage3_31[23],stage3_30[36],stage3_29[36]}
   );
   gpc606_5 gpc3674 (
      {stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100], stage2_29[101], stage2_29[102]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[11],stage3_31[24],stage3_30[37],stage3_29[37]}
   );
   gpc606_5 gpc3675 (
      {stage2_29[103], stage2_29[104], stage2_29[105], stage2_29[106], stage2_29[107], stage2_29[108]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[12],stage3_31[25],stage3_30[38],stage3_29[38]}
   );
   gpc606_5 gpc3676 (
      {stage2_29[109], stage2_29[110], stage2_29[111], stage2_29[112], stage2_29[113], stage2_29[114]},
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35]},
      {stage3_33[5],stage3_32[13],stage3_31[26],stage3_30[39],stage3_29[39]}
   );
   gpc606_5 gpc3677 (
      {stage2_29[115], stage2_29[116], stage2_29[117], stage2_29[118], stage2_29[119], stage2_29[120]},
      {stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41]},
      {stage3_33[6],stage3_32[14],stage3_31[27],stage3_30[40],stage3_29[40]}
   );
   gpc606_5 gpc3678 (
      {stage2_29[121], stage2_29[122], stage2_29[123], stage2_29[124], stage2_29[125], stage2_29[126]},
      {stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46], stage2_31[47]},
      {stage3_33[7],stage3_32[15],stage3_31[28],stage3_30[41],stage3_29[41]}
   );
   gpc606_5 gpc3679 (
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[8],stage3_32[16],stage3_31[29],stage3_30[42]}
   );
   gpc606_5 gpc3680 (
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[9],stage3_32[17],stage3_31[30],stage3_30[43]}
   );
   gpc606_5 gpc3681 (
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[10],stage3_32[18],stage3_31[31],stage3_30[44]}
   );
   gpc615_5 gpc3682 (
      {stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[3],stage3_33[11],stage3_32[19],stage3_31[32]}
   );
   gpc615_5 gpc3683 (
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57]},
      {stage2_32[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[4],stage3_33[12],stage3_32[20],stage3_31[33]}
   );
   gpc615_5 gpc3684 (
      {stage2_31[58], stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62]},
      {stage2_32[20]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[5],stage3_33[13],stage3_32[21],stage3_31[34]}
   );
   gpc615_5 gpc3685 (
      {stage2_31[63], stage2_31[64], stage2_31[65], stage2_31[66], stage2_31[67]},
      {stage2_32[21]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[6],stage3_33[14],stage3_32[22],stage3_31[35]}
   );
   gpc615_5 gpc3686 (
      {stage2_31[68], stage2_31[69], stage2_31[70], stage2_31[71], stage2_31[72]},
      {stage2_32[22]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[7],stage3_33[15],stage3_32[23],stage3_31[36]}
   );
   gpc615_5 gpc3687 (
      {stage2_31[73], stage2_31[74], stage2_31[75], stage2_31[76], stage2_31[77]},
      {stage2_32[23]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[8],stage3_33[16],stage3_32[24],stage3_31[37]}
   );
   gpc615_5 gpc3688 (
      {stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_32[24]},
      {stage2_33[36], stage2_33[37], stage2_33[38], stage2_33[39], stage2_33[40], stage2_33[41]},
      {stage3_35[6],stage3_34[9],stage3_33[17],stage3_32[25],stage3_31[38]}
   );
   gpc606_5 gpc3689 (
      {stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[7],stage3_34[10],stage3_33[18],stage3_32[26]}
   );
   gpc615_5 gpc3690 (
      {stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage2_33[42]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[8],stage3_34[11],stage3_33[19],stage3_32[27]}
   );
   gpc615_5 gpc3691 (
      {stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40]},
      {stage2_33[43]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[9],stage3_34[12],stage3_33[20],stage3_32[28]}
   );
   gpc615_5 gpc3692 (
      {stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44], stage2_32[45]},
      {stage2_33[44]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[10],stage3_34[13],stage3_33[21],stage3_32[29]}
   );
   gpc606_5 gpc3693 (
      {stage2_33[45], stage2_33[46], stage2_33[47], stage2_33[48], stage2_33[49], stage2_33[50]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[4],stage3_35[11],stage3_34[14],stage3_33[22]}
   );
   gpc606_5 gpc3694 (
      {stage2_33[51], stage2_33[52], stage2_33[53], stage2_33[54], stage2_33[55], stage2_33[56]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[5],stage3_35[12],stage3_34[15],stage3_33[23]}
   );
   gpc1_1 gpc3695 (
      {stage2_1[48]},
      {stage3_1[18]}
   );
   gpc1_1 gpc3696 (
      {stage2_1[49]},
      {stage3_1[19]}
   );
   gpc1_1 gpc3697 (
      {stage2_1[50]},
      {stage3_1[20]}
   );
   gpc1_1 gpc3698 (
      {stage2_1[51]},
      {stage3_1[21]}
   );
   gpc1_1 gpc3699 (
      {stage2_1[52]},
      {stage3_1[22]}
   );
   gpc1_1 gpc3700 (
      {stage2_1[53]},
      {stage3_1[23]}
   );
   gpc1_1 gpc3701 (
      {stage2_1[54]},
      {stage3_1[24]}
   );
   gpc1_1 gpc3702 (
      {stage2_1[55]},
      {stage3_1[25]}
   );
   gpc1_1 gpc3703 (
      {stage2_2[81]},
      {stage3_2[22]}
   );
   gpc1_1 gpc3704 (
      {stage2_2[82]},
      {stage3_2[23]}
   );
   gpc1_1 gpc3705 (
      {stage2_2[83]},
      {stage3_2[24]}
   );
   gpc1_1 gpc3706 (
      {stage2_2[84]},
      {stage3_2[25]}
   );
   gpc1_1 gpc3707 (
      {stage2_2[85]},
      {stage3_2[26]}
   );
   gpc1_1 gpc3708 (
      {stage2_2[86]},
      {stage3_2[27]}
   );
   gpc1_1 gpc3709 (
      {stage2_2[87]},
      {stage3_2[28]}
   );
   gpc1_1 gpc3710 (
      {stage2_2[88]},
      {stage3_2[29]}
   );
   gpc1_1 gpc3711 (
      {stage2_2[89]},
      {stage3_2[30]}
   );
   gpc1_1 gpc3712 (
      {stage2_2[90]},
      {stage3_2[31]}
   );
   gpc1_1 gpc3713 (
      {stage2_2[91]},
      {stage3_2[32]}
   );
   gpc1_1 gpc3714 (
      {stage2_2[92]},
      {stage3_2[33]}
   );
   gpc1_1 gpc3715 (
      {stage2_2[93]},
      {stage3_2[34]}
   );
   gpc1_1 gpc3716 (
      {stage2_2[94]},
      {stage3_2[35]}
   );
   gpc1_1 gpc3717 (
      {stage2_4[114]},
      {stage3_4[42]}
   );
   gpc1_1 gpc3718 (
      {stage2_4[115]},
      {stage3_4[43]}
   );
   gpc1_1 gpc3719 (
      {stage2_4[116]},
      {stage3_4[44]}
   );
   gpc1_1 gpc3720 (
      {stage2_4[117]},
      {stage3_4[45]}
   );
   gpc1_1 gpc3721 (
      {stage2_4[118]},
      {stage3_4[46]}
   );
   gpc1_1 gpc3722 (
      {stage2_5[72]},
      {stage3_5[37]}
   );
   gpc1_1 gpc3723 (
      {stage2_5[73]},
      {stage3_5[38]}
   );
   gpc1_1 gpc3724 (
      {stage2_5[74]},
      {stage3_5[39]}
   );
   gpc1_1 gpc3725 (
      {stage2_5[75]},
      {stage3_5[40]}
   );
   gpc1_1 gpc3726 (
      {stage2_5[76]},
      {stage3_5[41]}
   );
   gpc1_1 gpc3727 (
      {stage2_5[77]},
      {stage3_5[42]}
   );
   gpc1_1 gpc3728 (
      {stage2_5[78]},
      {stage3_5[43]}
   );
   gpc1_1 gpc3729 (
      {stage2_5[79]},
      {stage3_5[44]}
   );
   gpc1_1 gpc3730 (
      {stage2_5[80]},
      {stage3_5[45]}
   );
   gpc1_1 gpc3731 (
      {stage2_5[81]},
      {stage3_5[46]}
   );
   gpc1_1 gpc3732 (
      {stage2_5[82]},
      {stage3_5[47]}
   );
   gpc1_1 gpc3733 (
      {stage2_5[83]},
      {stage3_5[48]}
   );
   gpc1_1 gpc3734 (
      {stage2_5[84]},
      {stage3_5[49]}
   );
   gpc1_1 gpc3735 (
      {stage2_5[85]},
      {stage3_5[50]}
   );
   gpc1_1 gpc3736 (
      {stage2_5[86]},
      {stage3_5[51]}
   );
   gpc1_1 gpc3737 (
      {stage2_5[87]},
      {stage3_5[52]}
   );
   gpc1_1 gpc3738 (
      {stage2_5[88]},
      {stage3_5[53]}
   );
   gpc1_1 gpc3739 (
      {stage2_5[89]},
      {stage3_5[54]}
   );
   gpc1_1 gpc3740 (
      {stage2_5[90]},
      {stage3_5[55]}
   );
   gpc1_1 gpc3741 (
      {stage2_5[91]},
      {stage3_5[56]}
   );
   gpc1_1 gpc3742 (
      {stage2_5[92]},
      {stage3_5[57]}
   );
   gpc1_1 gpc3743 (
      {stage2_5[93]},
      {stage3_5[58]}
   );
   gpc1_1 gpc3744 (
      {stage2_6[89]},
      {stage3_6[31]}
   );
   gpc1_1 gpc3745 (
      {stage2_6[90]},
      {stage3_6[32]}
   );
   gpc1_1 gpc3746 (
      {stage2_6[91]},
      {stage3_6[33]}
   );
   gpc1_1 gpc3747 (
      {stage2_6[92]},
      {stage3_6[34]}
   );
   gpc1_1 gpc3748 (
      {stage2_6[93]},
      {stage3_6[35]}
   );
   gpc1_1 gpc3749 (
      {stage2_6[94]},
      {stage3_6[36]}
   );
   gpc1_1 gpc3750 (
      {stage2_6[95]},
      {stage3_6[37]}
   );
   gpc1_1 gpc3751 (
      {stage2_7[102]},
      {stage3_7[40]}
   );
   gpc1_1 gpc3752 (
      {stage2_7[103]},
      {stage3_7[41]}
   );
   gpc1_1 gpc3753 (
      {stage2_7[104]},
      {stage3_7[42]}
   );
   gpc1_1 gpc3754 (
      {stage2_7[105]},
      {stage3_7[43]}
   );
   gpc1_1 gpc3755 (
      {stage2_7[106]},
      {stage3_7[44]}
   );
   gpc1_1 gpc3756 (
      {stage2_7[107]},
      {stage3_7[45]}
   );
   gpc1_1 gpc3757 (
      {stage2_7[108]},
      {stage3_7[46]}
   );
   gpc1_1 gpc3758 (
      {stage2_8[43]},
      {stage3_8[38]}
   );
   gpc1_1 gpc3759 (
      {stage2_8[44]},
      {stage3_8[39]}
   );
   gpc1_1 gpc3760 (
      {stage2_8[45]},
      {stage3_8[40]}
   );
   gpc1_1 gpc3761 (
      {stage2_8[46]},
      {stage3_8[41]}
   );
   gpc1_1 gpc3762 (
      {stage2_8[47]},
      {stage3_8[42]}
   );
   gpc1_1 gpc3763 (
      {stage2_8[48]},
      {stage3_8[43]}
   );
   gpc1_1 gpc3764 (
      {stage2_8[49]},
      {stage3_8[44]}
   );
   gpc1_1 gpc3765 (
      {stage2_8[50]},
      {stage3_8[45]}
   );
   gpc1_1 gpc3766 (
      {stage2_8[51]},
      {stage3_8[46]}
   );
   gpc1_1 gpc3767 (
      {stage2_8[52]},
      {stage3_8[47]}
   );
   gpc1_1 gpc3768 (
      {stage2_8[53]},
      {stage3_8[48]}
   );
   gpc1_1 gpc3769 (
      {stage2_8[54]},
      {stage3_8[49]}
   );
   gpc1_1 gpc3770 (
      {stage2_8[55]},
      {stage3_8[50]}
   );
   gpc1_1 gpc3771 (
      {stage2_8[56]},
      {stage3_8[51]}
   );
   gpc1_1 gpc3772 (
      {stage2_8[57]},
      {stage3_8[52]}
   );
   gpc1_1 gpc3773 (
      {stage2_8[58]},
      {stage3_8[53]}
   );
   gpc1_1 gpc3774 (
      {stage2_8[59]},
      {stage3_8[54]}
   );
   gpc1_1 gpc3775 (
      {stage2_8[60]},
      {stage3_8[55]}
   );
   gpc1_1 gpc3776 (
      {stage2_8[61]},
      {stage3_8[56]}
   );
   gpc1_1 gpc3777 (
      {stage2_8[62]},
      {stage3_8[57]}
   );
   gpc1_1 gpc3778 (
      {stage2_8[63]},
      {stage3_8[58]}
   );
   gpc1_1 gpc3779 (
      {stage2_8[64]},
      {stage3_8[59]}
   );
   gpc1_1 gpc3780 (
      {stage2_8[65]},
      {stage3_8[60]}
   );
   gpc1_1 gpc3781 (
      {stage2_8[66]},
      {stage3_8[61]}
   );
   gpc1_1 gpc3782 (
      {stage2_8[67]},
      {stage3_8[62]}
   );
   gpc1_1 gpc3783 (
      {stage2_8[68]},
      {stage3_8[63]}
   );
   gpc1_1 gpc3784 (
      {stage2_8[69]},
      {stage3_8[64]}
   );
   gpc1_1 gpc3785 (
      {stage2_8[70]},
      {stage3_8[65]}
   );
   gpc1_1 gpc3786 (
      {stage2_8[71]},
      {stage3_8[66]}
   );
   gpc1_1 gpc3787 (
      {stage2_8[72]},
      {stage3_8[67]}
   );
   gpc1_1 gpc3788 (
      {stage2_8[73]},
      {stage3_8[68]}
   );
   gpc1_1 gpc3789 (
      {stage2_8[74]},
      {stage3_8[69]}
   );
   gpc1_1 gpc3790 (
      {stage2_8[75]},
      {stage3_8[70]}
   );
   gpc1_1 gpc3791 (
      {stage2_8[76]},
      {stage3_8[71]}
   );
   gpc1_1 gpc3792 (
      {stage2_8[77]},
      {stage3_8[72]}
   );
   gpc1_1 gpc3793 (
      {stage2_8[78]},
      {stage3_8[73]}
   );
   gpc1_1 gpc3794 (
      {stage2_8[79]},
      {stage3_8[74]}
   );
   gpc1_1 gpc3795 (
      {stage2_8[80]},
      {stage3_8[75]}
   );
   gpc1_1 gpc3796 (
      {stage2_8[81]},
      {stage3_8[76]}
   );
   gpc1_1 gpc3797 (
      {stage2_8[82]},
      {stage3_8[77]}
   );
   gpc1_1 gpc3798 (
      {stage2_8[83]},
      {stage3_8[78]}
   );
   gpc1_1 gpc3799 (
      {stage2_8[84]},
      {stage3_8[79]}
   );
   gpc1_1 gpc3800 (
      {stage2_8[85]},
      {stage3_8[80]}
   );
   gpc1_1 gpc3801 (
      {stage2_8[86]},
      {stage3_8[81]}
   );
   gpc1_1 gpc3802 (
      {stage2_8[87]},
      {stage3_8[82]}
   );
   gpc1_1 gpc3803 (
      {stage2_8[88]},
      {stage3_8[83]}
   );
   gpc1_1 gpc3804 (
      {stage2_8[89]},
      {stage3_8[84]}
   );
   gpc1_1 gpc3805 (
      {stage2_8[90]},
      {stage3_8[85]}
   );
   gpc1_1 gpc3806 (
      {stage2_8[91]},
      {stage3_8[86]}
   );
   gpc1_1 gpc3807 (
      {stage2_8[92]},
      {stage3_8[87]}
   );
   gpc1_1 gpc3808 (
      {stage2_8[93]},
      {stage3_8[88]}
   );
   gpc1_1 gpc3809 (
      {stage2_8[94]},
      {stage3_8[89]}
   );
   gpc1_1 gpc3810 (
      {stage2_8[95]},
      {stage3_8[90]}
   );
   gpc1_1 gpc3811 (
      {stage2_8[96]},
      {stage3_8[91]}
   );
   gpc1_1 gpc3812 (
      {stage2_8[97]},
      {stage3_8[92]}
   );
   gpc1_1 gpc3813 (
      {stage2_9[83]},
      {stage3_9[25]}
   );
   gpc1_1 gpc3814 (
      {stage2_9[84]},
      {stage3_9[26]}
   );
   gpc1_1 gpc3815 (
      {stage2_9[85]},
      {stage3_9[27]}
   );
   gpc1_1 gpc3816 (
      {stage2_9[86]},
      {stage3_9[28]}
   );
   gpc1_1 gpc3817 (
      {stage2_9[87]},
      {stage3_9[29]}
   );
   gpc1_1 gpc3818 (
      {stage2_9[88]},
      {stage3_9[30]}
   );
   gpc1_1 gpc3819 (
      {stage2_9[89]},
      {stage3_9[31]}
   );
   gpc1_1 gpc3820 (
      {stage2_9[90]},
      {stage3_9[32]}
   );
   gpc1_1 gpc3821 (
      {stage2_9[91]},
      {stage3_9[33]}
   );
   gpc1_1 gpc3822 (
      {stage2_9[92]},
      {stage3_9[34]}
   );
   gpc1_1 gpc3823 (
      {stage2_9[93]},
      {stage3_9[35]}
   );
   gpc1_1 gpc3824 (
      {stage2_9[94]},
      {stage3_9[36]}
   );
   gpc1_1 gpc3825 (
      {stage2_9[95]},
      {stage3_9[37]}
   );
   gpc1_1 gpc3826 (
      {stage2_9[96]},
      {stage3_9[38]}
   );
   gpc1_1 gpc3827 (
      {stage2_9[97]},
      {stage3_9[39]}
   );
   gpc1_1 gpc3828 (
      {stage2_9[98]},
      {stage3_9[40]}
   );
   gpc1_1 gpc3829 (
      {stage2_9[99]},
      {stage3_9[41]}
   );
   gpc1_1 gpc3830 (
      {stage2_9[100]},
      {stage3_9[42]}
   );
   gpc1_1 gpc3831 (
      {stage2_9[101]},
      {stage3_9[43]}
   );
   gpc1_1 gpc3832 (
      {stage2_9[102]},
      {stage3_9[44]}
   );
   gpc1_1 gpc3833 (
      {stage2_9[103]},
      {stage3_9[45]}
   );
   gpc1_1 gpc3834 (
      {stage2_9[104]},
      {stage3_9[46]}
   );
   gpc1_1 gpc3835 (
      {stage2_9[105]},
      {stage3_9[47]}
   );
   gpc1_1 gpc3836 (
      {stage2_9[106]},
      {stage3_9[48]}
   );
   gpc1_1 gpc3837 (
      {stage2_9[107]},
      {stage3_9[49]}
   );
   gpc1_1 gpc3838 (
      {stage2_10[87]},
      {stage3_10[30]}
   );
   gpc1_1 gpc3839 (
      {stage2_10[88]},
      {stage3_10[31]}
   );
   gpc1_1 gpc3840 (
      {stage2_10[89]},
      {stage3_10[32]}
   );
   gpc1_1 gpc3841 (
      {stage2_10[90]},
      {stage3_10[33]}
   );
   gpc1_1 gpc3842 (
      {stage2_10[91]},
      {stage3_10[34]}
   );
   gpc1_1 gpc3843 (
      {stage2_10[92]},
      {stage3_10[35]}
   );
   gpc1_1 gpc3844 (
      {stage2_10[93]},
      {stage3_10[36]}
   );
   gpc1_1 gpc3845 (
      {stage2_10[94]},
      {stage3_10[37]}
   );
   gpc1_1 gpc3846 (
      {stage2_11[110]},
      {stage3_11[49]}
   );
   gpc1_1 gpc3847 (
      {stage2_11[111]},
      {stage3_11[50]}
   );
   gpc1_1 gpc3848 (
      {stage2_11[112]},
      {stage3_11[51]}
   );
   gpc1_1 gpc3849 (
      {stage2_11[113]},
      {stage3_11[52]}
   );
   gpc1_1 gpc3850 (
      {stage2_11[114]},
      {stage3_11[53]}
   );
   gpc1_1 gpc3851 (
      {stage2_11[115]},
      {stage3_11[54]}
   );
   gpc1_1 gpc3852 (
      {stage2_12[92]},
      {stage3_12[37]}
   );
   gpc1_1 gpc3853 (
      {stage2_12[93]},
      {stage3_12[38]}
   );
   gpc1_1 gpc3854 (
      {stage2_12[94]},
      {stage3_12[39]}
   );
   gpc1_1 gpc3855 (
      {stage2_12[95]},
      {stage3_12[40]}
   );
   gpc1_1 gpc3856 (
      {stage2_12[96]},
      {stage3_12[41]}
   );
   gpc1_1 gpc3857 (
      {stage2_12[97]},
      {stage3_12[42]}
   );
   gpc1_1 gpc3858 (
      {stage2_12[98]},
      {stage3_12[43]}
   );
   gpc1_1 gpc3859 (
      {stage2_12[99]},
      {stage3_12[44]}
   );
   gpc1_1 gpc3860 (
      {stage2_12[100]},
      {stage3_12[45]}
   );
   gpc1_1 gpc3861 (
      {stage2_12[101]},
      {stage3_12[46]}
   );
   gpc1_1 gpc3862 (
      {stage2_13[120]},
      {stage3_13[33]}
   );
   gpc1_1 gpc3863 (
      {stage2_13[121]},
      {stage3_13[34]}
   );
   gpc1_1 gpc3864 (
      {stage2_13[122]},
      {stage3_13[35]}
   );
   gpc1_1 gpc3865 (
      {stage2_13[123]},
      {stage3_13[36]}
   );
   gpc1_1 gpc3866 (
      {stage2_14[56]},
      {stage3_14[42]}
   );
   gpc1_1 gpc3867 (
      {stage2_14[57]},
      {stage3_14[43]}
   );
   gpc1_1 gpc3868 (
      {stage2_14[58]},
      {stage3_14[44]}
   );
   gpc1_1 gpc3869 (
      {stage2_14[59]},
      {stage3_14[45]}
   );
   gpc1_1 gpc3870 (
      {stage2_14[60]},
      {stage3_14[46]}
   );
   gpc1_1 gpc3871 (
      {stage2_14[61]},
      {stage3_14[47]}
   );
   gpc1_1 gpc3872 (
      {stage2_14[62]},
      {stage3_14[48]}
   );
   gpc1_1 gpc3873 (
      {stage2_14[63]},
      {stage3_14[49]}
   );
   gpc1_1 gpc3874 (
      {stage2_14[64]},
      {stage3_14[50]}
   );
   gpc1_1 gpc3875 (
      {stage2_14[65]},
      {stage3_14[51]}
   );
   gpc1_1 gpc3876 (
      {stage2_14[66]},
      {stage3_14[52]}
   );
   gpc1_1 gpc3877 (
      {stage2_14[67]},
      {stage3_14[53]}
   );
   gpc1_1 gpc3878 (
      {stage2_14[68]},
      {stage3_14[54]}
   );
   gpc1_1 gpc3879 (
      {stage2_14[69]},
      {stage3_14[55]}
   );
   gpc1_1 gpc3880 (
      {stage2_15[70]},
      {stage3_15[43]}
   );
   gpc1_1 gpc3881 (
      {stage2_15[71]},
      {stage3_15[44]}
   );
   gpc1_1 gpc3882 (
      {stage2_15[72]},
      {stage3_15[45]}
   );
   gpc1_1 gpc3883 (
      {stage2_15[73]},
      {stage3_15[46]}
   );
   gpc1_1 gpc3884 (
      {stage2_15[74]},
      {stage3_15[47]}
   );
   gpc1_1 gpc3885 (
      {stage2_15[75]},
      {stage3_15[48]}
   );
   gpc1_1 gpc3886 (
      {stage2_15[76]},
      {stage3_15[49]}
   );
   gpc1_1 gpc3887 (
      {stage2_15[77]},
      {stage3_15[50]}
   );
   gpc1_1 gpc3888 (
      {stage2_15[78]},
      {stage3_15[51]}
   );
   gpc1_1 gpc3889 (
      {stage2_15[79]},
      {stage3_15[52]}
   );
   gpc1_1 gpc3890 (
      {stage2_15[80]},
      {stage3_15[53]}
   );
   gpc1_1 gpc3891 (
      {stage2_15[81]},
      {stage3_15[54]}
   );
   gpc1_1 gpc3892 (
      {stage2_15[82]},
      {stage3_15[55]}
   );
   gpc1_1 gpc3893 (
      {stage2_15[83]},
      {stage3_15[56]}
   );
   gpc1_1 gpc3894 (
      {stage2_15[84]},
      {stage3_15[57]}
   );
   gpc1_1 gpc3895 (
      {stage2_15[85]},
      {stage3_15[58]}
   );
   gpc1_1 gpc3896 (
      {stage2_15[86]},
      {stage3_15[59]}
   );
   gpc1_1 gpc3897 (
      {stage2_15[87]},
      {stage3_15[60]}
   );
   gpc1_1 gpc3898 (
      {stage2_15[88]},
      {stage3_15[61]}
   );
   gpc1_1 gpc3899 (
      {stage2_15[89]},
      {stage3_15[62]}
   );
   gpc1_1 gpc3900 (
      {stage2_15[90]},
      {stage3_15[63]}
   );
   gpc1_1 gpc3901 (
      {stage2_15[91]},
      {stage3_15[64]}
   );
   gpc1_1 gpc3902 (
      {stage2_15[92]},
      {stage3_15[65]}
   );
   gpc1_1 gpc3903 (
      {stage2_15[93]},
      {stage3_15[66]}
   );
   gpc1_1 gpc3904 (
      {stage2_15[94]},
      {stage3_15[67]}
   );
   gpc1_1 gpc3905 (
      {stage2_15[95]},
      {stage3_15[68]}
   );
   gpc1_1 gpc3906 (
      {stage2_15[96]},
      {stage3_15[69]}
   );
   gpc1_1 gpc3907 (
      {stage2_15[97]},
      {stage3_15[70]}
   );
   gpc1_1 gpc3908 (
      {stage2_16[83]},
      {stage3_16[25]}
   );
   gpc1_1 gpc3909 (
      {stage2_16[84]},
      {stage3_16[26]}
   );
   gpc1_1 gpc3910 (
      {stage2_16[85]},
      {stage3_16[27]}
   );
   gpc1_1 gpc3911 (
      {stage2_16[86]},
      {stage3_16[28]}
   );
   gpc1_1 gpc3912 (
      {stage2_16[87]},
      {stage3_16[29]}
   );
   gpc1_1 gpc3913 (
      {stage2_16[88]},
      {stage3_16[30]}
   );
   gpc1_1 gpc3914 (
      {stage2_16[89]},
      {stage3_16[31]}
   );
   gpc1_1 gpc3915 (
      {stage2_16[90]},
      {stage3_16[32]}
   );
   gpc1_1 gpc3916 (
      {stage2_16[91]},
      {stage3_16[33]}
   );
   gpc1_1 gpc3917 (
      {stage2_16[92]},
      {stage3_16[34]}
   );
   gpc1_1 gpc3918 (
      {stage2_16[93]},
      {stage3_16[35]}
   );
   gpc1_1 gpc3919 (
      {stage2_16[94]},
      {stage3_16[36]}
   );
   gpc1_1 gpc3920 (
      {stage2_16[95]},
      {stage3_16[37]}
   );
   gpc1_1 gpc3921 (
      {stage2_16[96]},
      {stage3_16[38]}
   );
   gpc1_1 gpc3922 (
      {stage2_16[97]},
      {stage3_16[39]}
   );
   gpc1_1 gpc3923 (
      {stage2_16[98]},
      {stage3_16[40]}
   );
   gpc1_1 gpc3924 (
      {stage2_16[99]},
      {stage3_16[41]}
   );
   gpc1_1 gpc3925 (
      {stage2_16[100]},
      {stage3_16[42]}
   );
   gpc1_1 gpc3926 (
      {stage2_16[101]},
      {stage3_16[43]}
   );
   gpc1_1 gpc3927 (
      {stage2_16[102]},
      {stage3_16[44]}
   );
   gpc1_1 gpc3928 (
      {stage2_16[103]},
      {stage3_16[45]}
   );
   gpc1_1 gpc3929 (
      {stage2_16[104]},
      {stage3_16[46]}
   );
   gpc1_1 gpc3930 (
      {stage2_16[105]},
      {stage3_16[47]}
   );
   gpc1_1 gpc3931 (
      {stage2_16[106]},
      {stage3_16[48]}
   );
   gpc1_1 gpc3932 (
      {stage2_16[107]},
      {stage3_16[49]}
   );
   gpc1_1 gpc3933 (
      {stage2_16[108]},
      {stage3_16[50]}
   );
   gpc1_1 gpc3934 (
      {stage2_16[109]},
      {stage3_16[51]}
   );
   gpc1_1 gpc3935 (
      {stage2_16[110]},
      {stage3_16[52]}
   );
   gpc1_1 gpc3936 (
      {stage2_16[111]},
      {stage3_16[53]}
   );
   gpc1_1 gpc3937 (
      {stage2_16[112]},
      {stage3_16[54]}
   );
   gpc1_1 gpc3938 (
      {stage2_16[113]},
      {stage3_16[55]}
   );
   gpc1_1 gpc3939 (
      {stage2_16[114]},
      {stage3_16[56]}
   );
   gpc1_1 gpc3940 (
      {stage2_16[115]},
      {stage3_16[57]}
   );
   gpc1_1 gpc3941 (
      {stage2_16[116]},
      {stage3_16[58]}
   );
   gpc1_1 gpc3942 (
      {stage2_16[117]},
      {stage3_16[59]}
   );
   gpc1_1 gpc3943 (
      {stage2_16[118]},
      {stage3_16[60]}
   );
   gpc1_1 gpc3944 (
      {stage2_16[119]},
      {stage3_16[61]}
   );
   gpc1_1 gpc3945 (
      {stage2_16[120]},
      {stage3_16[62]}
   );
   gpc1_1 gpc3946 (
      {stage2_16[121]},
      {stage3_16[63]}
   );
   gpc1_1 gpc3947 (
      {stage2_16[122]},
      {stage3_16[64]}
   );
   gpc1_1 gpc3948 (
      {stage2_16[123]},
      {stage3_16[65]}
   );
   gpc1_1 gpc3949 (
      {stage2_16[124]},
      {stage3_16[66]}
   );
   gpc1_1 gpc3950 (
      {stage2_17[75]},
      {stage3_17[24]}
   );
   gpc1_1 gpc3951 (
      {stage2_17[76]},
      {stage3_17[25]}
   );
   gpc1_1 gpc3952 (
      {stage2_17[77]},
      {stage3_17[26]}
   );
   gpc1_1 gpc3953 (
      {stage2_17[78]},
      {stage3_17[27]}
   );
   gpc1_1 gpc3954 (
      {stage2_17[79]},
      {stage3_17[28]}
   );
   gpc1_1 gpc3955 (
      {stage2_17[80]},
      {stage3_17[29]}
   );
   gpc1_1 gpc3956 (
      {stage2_17[81]},
      {stage3_17[30]}
   );
   gpc1_1 gpc3957 (
      {stage2_17[82]},
      {stage3_17[31]}
   );
   gpc1_1 gpc3958 (
      {stage2_17[83]},
      {stage3_17[32]}
   );
   gpc1_1 gpc3959 (
      {stage2_17[84]},
      {stage3_17[33]}
   );
   gpc1_1 gpc3960 (
      {stage2_17[85]},
      {stage3_17[34]}
   );
   gpc1_1 gpc3961 (
      {stage2_17[86]},
      {stage3_17[35]}
   );
   gpc1_1 gpc3962 (
      {stage2_17[87]},
      {stage3_17[36]}
   );
   gpc1_1 gpc3963 (
      {stage2_17[88]},
      {stage3_17[37]}
   );
   gpc1_1 gpc3964 (
      {stage2_17[89]},
      {stage3_17[38]}
   );
   gpc1_1 gpc3965 (
      {stage2_17[90]},
      {stage3_17[39]}
   );
   gpc1_1 gpc3966 (
      {stage2_17[91]},
      {stage3_17[40]}
   );
   gpc1_1 gpc3967 (
      {stage2_17[92]},
      {stage3_17[41]}
   );
   gpc1_1 gpc3968 (
      {stage2_17[93]},
      {stage3_17[42]}
   );
   gpc1_1 gpc3969 (
      {stage2_17[94]},
      {stage3_17[43]}
   );
   gpc1_1 gpc3970 (
      {stage2_17[95]},
      {stage3_17[44]}
   );
   gpc1_1 gpc3971 (
      {stage2_17[96]},
      {stage3_17[45]}
   );
   gpc1_1 gpc3972 (
      {stage2_17[97]},
      {stage3_17[46]}
   );
   gpc1_1 gpc3973 (
      {stage2_17[98]},
      {stage3_17[47]}
   );
   gpc1_1 gpc3974 (
      {stage2_17[99]},
      {stage3_17[48]}
   );
   gpc1_1 gpc3975 (
      {stage2_17[100]},
      {stage3_17[49]}
   );
   gpc1_1 gpc3976 (
      {stage2_17[101]},
      {stage3_17[50]}
   );
   gpc1_1 gpc3977 (
      {stage2_17[102]},
      {stage3_17[51]}
   );
   gpc1_1 gpc3978 (
      {stage2_17[103]},
      {stage3_17[52]}
   );
   gpc1_1 gpc3979 (
      {stage2_17[104]},
      {stage3_17[53]}
   );
   gpc1_1 gpc3980 (
      {stage2_17[105]},
      {stage3_17[54]}
   );
   gpc1_1 gpc3981 (
      {stage2_17[106]},
      {stage3_17[55]}
   );
   gpc1_1 gpc3982 (
      {stage2_17[107]},
      {stage3_17[56]}
   );
   gpc1_1 gpc3983 (
      {stage2_17[108]},
      {stage3_17[57]}
   );
   gpc1_1 gpc3984 (
      {stage2_17[109]},
      {stage3_17[58]}
   );
   gpc1_1 gpc3985 (
      {stage2_17[110]},
      {stage3_17[59]}
   );
   gpc1_1 gpc3986 (
      {stage2_17[111]},
      {stage3_17[60]}
   );
   gpc1_1 gpc3987 (
      {stage2_17[112]},
      {stage3_17[61]}
   );
   gpc1_1 gpc3988 (
      {stage2_17[113]},
      {stage3_17[62]}
   );
   gpc1_1 gpc3989 (
      {stage2_17[114]},
      {stage3_17[63]}
   );
   gpc1_1 gpc3990 (
      {stage2_17[115]},
      {stage3_17[64]}
   );
   gpc1_1 gpc3991 (
      {stage2_17[116]},
      {stage3_17[65]}
   );
   gpc1_1 gpc3992 (
      {stage2_17[117]},
      {stage3_17[66]}
   );
   gpc1_1 gpc3993 (
      {stage2_17[118]},
      {stage3_17[67]}
   );
   gpc1_1 gpc3994 (
      {stage2_17[119]},
      {stage3_17[68]}
   );
   gpc1_1 gpc3995 (
      {stage2_17[120]},
      {stage3_17[69]}
   );
   gpc1_1 gpc3996 (
      {stage2_17[121]},
      {stage3_17[70]}
   );
   gpc1_1 gpc3997 (
      {stage2_17[122]},
      {stage3_17[71]}
   );
   gpc1_1 gpc3998 (
      {stage2_17[123]},
      {stage3_17[72]}
   );
   gpc1_1 gpc3999 (
      {stage2_17[124]},
      {stage3_17[73]}
   );
   gpc1_1 gpc4000 (
      {stage2_17[125]},
      {stage3_17[74]}
   );
   gpc1_1 gpc4001 (
      {stage2_17[126]},
      {stage3_17[75]}
   );
   gpc1_1 gpc4002 (
      {stage2_17[127]},
      {stage3_17[76]}
   );
   gpc1_1 gpc4003 (
      {stage2_19[64]},
      {stage3_19[36]}
   );
   gpc1_1 gpc4004 (
      {stage2_19[65]},
      {stage3_19[37]}
   );
   gpc1_1 gpc4005 (
      {stage2_19[66]},
      {stage3_19[38]}
   );
   gpc1_1 gpc4006 (
      {stage2_19[67]},
      {stage3_19[39]}
   );
   gpc1_1 gpc4007 (
      {stage2_19[68]},
      {stage3_19[40]}
   );
   gpc1_1 gpc4008 (
      {stage2_19[69]},
      {stage3_19[41]}
   );
   gpc1_1 gpc4009 (
      {stage2_19[70]},
      {stage3_19[42]}
   );
   gpc1_1 gpc4010 (
      {stage2_19[71]},
      {stage3_19[43]}
   );
   gpc1_1 gpc4011 (
      {stage2_19[72]},
      {stage3_19[44]}
   );
   gpc1_1 gpc4012 (
      {stage2_19[73]},
      {stage3_19[45]}
   );
   gpc1_1 gpc4013 (
      {stage2_19[74]},
      {stage3_19[46]}
   );
   gpc1_1 gpc4014 (
      {stage2_19[75]},
      {stage3_19[47]}
   );
   gpc1_1 gpc4015 (
      {stage2_19[76]},
      {stage3_19[48]}
   );
   gpc1_1 gpc4016 (
      {stage2_19[77]},
      {stage3_19[49]}
   );
   gpc1_1 gpc4017 (
      {stage2_19[78]},
      {stage3_19[50]}
   );
   gpc1_1 gpc4018 (
      {stage2_19[79]},
      {stage3_19[51]}
   );
   gpc1_1 gpc4019 (
      {stage2_19[80]},
      {stage3_19[52]}
   );
   gpc1_1 gpc4020 (
      {stage2_19[81]},
      {stage3_19[53]}
   );
   gpc1_1 gpc4021 (
      {stage2_19[82]},
      {stage3_19[54]}
   );
   gpc1_1 gpc4022 (
      {stage2_19[83]},
      {stage3_19[55]}
   );
   gpc1_1 gpc4023 (
      {stage2_19[84]},
      {stage3_19[56]}
   );
   gpc1_1 gpc4024 (
      {stage2_19[85]},
      {stage3_19[57]}
   );
   gpc1_1 gpc4025 (
      {stage2_19[86]},
      {stage3_19[58]}
   );
   gpc1_1 gpc4026 (
      {stage2_19[87]},
      {stage3_19[59]}
   );
   gpc1_1 gpc4027 (
      {stage2_19[88]},
      {stage3_19[60]}
   );
   gpc1_1 gpc4028 (
      {stage2_19[89]},
      {stage3_19[61]}
   );
   gpc1_1 gpc4029 (
      {stage2_19[90]},
      {stage3_19[62]}
   );
   gpc1_1 gpc4030 (
      {stage2_19[91]},
      {stage3_19[63]}
   );
   gpc1_1 gpc4031 (
      {stage2_19[92]},
      {stage3_19[64]}
   );
   gpc1_1 gpc4032 (
      {stage2_19[93]},
      {stage3_19[65]}
   );
   gpc1_1 gpc4033 (
      {stage2_19[94]},
      {stage3_19[66]}
   );
   gpc1_1 gpc4034 (
      {stage2_19[95]},
      {stage3_19[67]}
   );
   gpc1_1 gpc4035 (
      {stage2_19[96]},
      {stage3_19[68]}
   );
   gpc1_1 gpc4036 (
      {stage2_19[97]},
      {stage3_19[69]}
   );
   gpc1_1 gpc4037 (
      {stage2_21[96]},
      {stage3_21[34]}
   );
   gpc1_1 gpc4038 (
      {stage2_21[97]},
      {stage3_21[35]}
   );
   gpc1_1 gpc4039 (
      {stage2_21[98]},
      {stage3_21[36]}
   );
   gpc1_1 gpc4040 (
      {stage2_21[99]},
      {stage3_21[37]}
   );
   gpc1_1 gpc4041 (
      {stage2_21[100]},
      {stage3_21[38]}
   );
   gpc1_1 gpc4042 (
      {stage2_21[101]},
      {stage3_21[39]}
   );
   gpc1_1 gpc4043 (
      {stage2_21[102]},
      {stage3_21[40]}
   );
   gpc1_1 gpc4044 (
      {stage2_21[103]},
      {stage3_21[41]}
   );
   gpc1_1 gpc4045 (
      {stage2_21[104]},
      {stage3_21[42]}
   );
   gpc1_1 gpc4046 (
      {stage2_21[105]},
      {stage3_21[43]}
   );
   gpc1_1 gpc4047 (
      {stage2_21[106]},
      {stage3_21[44]}
   );
   gpc1_1 gpc4048 (
      {stage2_21[107]},
      {stage3_21[45]}
   );
   gpc1_1 gpc4049 (
      {stage2_21[108]},
      {stage3_21[46]}
   );
   gpc1_1 gpc4050 (
      {stage2_21[109]},
      {stage3_21[47]}
   );
   gpc1_1 gpc4051 (
      {stage2_21[110]},
      {stage3_21[48]}
   );
   gpc1_1 gpc4052 (
      {stage2_21[111]},
      {stage3_21[49]}
   );
   gpc1_1 gpc4053 (
      {stage2_21[112]},
      {stage3_21[50]}
   );
   gpc1_1 gpc4054 (
      {stage2_21[113]},
      {stage3_21[51]}
   );
   gpc1_1 gpc4055 (
      {stage2_21[114]},
      {stage3_21[52]}
   );
   gpc1_1 gpc4056 (
      {stage2_21[115]},
      {stage3_21[53]}
   );
   gpc1_1 gpc4057 (
      {stage2_21[116]},
      {stage3_21[54]}
   );
   gpc1_1 gpc4058 (
      {stage2_21[117]},
      {stage3_21[55]}
   );
   gpc1_1 gpc4059 (
      {stage2_21[118]},
      {stage3_21[56]}
   );
   gpc1_1 gpc4060 (
      {stage2_21[119]},
      {stage3_21[57]}
   );
   gpc1_1 gpc4061 (
      {stage2_21[120]},
      {stage3_21[58]}
   );
   gpc1_1 gpc4062 (
      {stage2_21[121]},
      {stage3_21[59]}
   );
   gpc1_1 gpc4063 (
      {stage2_21[122]},
      {stage3_21[60]}
   );
   gpc1_1 gpc4064 (
      {stage2_21[123]},
      {stage3_21[61]}
   );
   gpc1_1 gpc4065 (
      {stage2_21[124]},
      {stage3_21[62]}
   );
   gpc1_1 gpc4066 (
      {stage2_22[87]},
      {stage3_22[43]}
   );
   gpc1_1 gpc4067 (
      {stage2_22[88]},
      {stage3_22[44]}
   );
   gpc1_1 gpc4068 (
      {stage2_22[89]},
      {stage3_22[45]}
   );
   gpc1_1 gpc4069 (
      {stage2_22[90]},
      {stage3_22[46]}
   );
   gpc1_1 gpc4070 (
      {stage2_22[91]},
      {stage3_22[47]}
   );
   gpc1_1 gpc4071 (
      {stage2_22[92]},
      {stage3_22[48]}
   );
   gpc1_1 gpc4072 (
      {stage2_22[93]},
      {stage3_22[49]}
   );
   gpc1_1 gpc4073 (
      {stage2_22[94]},
      {stage3_22[50]}
   );
   gpc1_1 gpc4074 (
      {stage2_24[66]},
      {stage3_24[37]}
   );
   gpc1_1 gpc4075 (
      {stage2_24[67]},
      {stage3_24[38]}
   );
   gpc1_1 gpc4076 (
      {stage2_24[68]},
      {stage3_24[39]}
   );
   gpc1_1 gpc4077 (
      {stage2_24[69]},
      {stage3_24[40]}
   );
   gpc1_1 gpc4078 (
      {stage2_24[70]},
      {stage3_24[41]}
   );
   gpc1_1 gpc4079 (
      {stage2_24[71]},
      {stage3_24[42]}
   );
   gpc1_1 gpc4080 (
      {stage2_24[72]},
      {stage3_24[43]}
   );
   gpc1_1 gpc4081 (
      {stage2_24[73]},
      {stage3_24[44]}
   );
   gpc1_1 gpc4082 (
      {stage2_24[74]},
      {stage3_24[45]}
   );
   gpc1_1 gpc4083 (
      {stage2_24[75]},
      {stage3_24[46]}
   );
   gpc1_1 gpc4084 (
      {stage2_24[76]},
      {stage3_24[47]}
   );
   gpc1_1 gpc4085 (
      {stage2_24[77]},
      {stage3_24[48]}
   );
   gpc1_1 gpc4086 (
      {stage2_24[78]},
      {stage3_24[49]}
   );
   gpc1_1 gpc4087 (
      {stage2_24[79]},
      {stage3_24[50]}
   );
   gpc1_1 gpc4088 (
      {stage2_24[80]},
      {stage3_24[51]}
   );
   gpc1_1 gpc4089 (
      {stage2_24[81]},
      {stage3_24[52]}
   );
   gpc1_1 gpc4090 (
      {stage2_24[82]},
      {stage3_24[53]}
   );
   gpc1_1 gpc4091 (
      {stage2_24[83]},
      {stage3_24[54]}
   );
   gpc1_1 gpc4092 (
      {stage2_24[84]},
      {stage3_24[55]}
   );
   gpc1_1 gpc4093 (
      {stage2_24[85]},
      {stage3_24[56]}
   );
   gpc1_1 gpc4094 (
      {stage2_24[86]},
      {stage3_24[57]}
   );
   gpc1_1 gpc4095 (
      {stage2_24[87]},
      {stage3_24[58]}
   );
   gpc1_1 gpc4096 (
      {stage2_24[88]},
      {stage3_24[59]}
   );
   gpc1_1 gpc4097 (
      {stage2_24[89]},
      {stage3_24[60]}
   );
   gpc1_1 gpc4098 (
      {stage2_25[84]},
      {stage3_25[30]}
   );
   gpc1_1 gpc4099 (
      {stage2_25[85]},
      {stage3_25[31]}
   );
   gpc1_1 gpc4100 (
      {stage2_25[86]},
      {stage3_25[32]}
   );
   gpc1_1 gpc4101 (
      {stage2_25[87]},
      {stage3_25[33]}
   );
   gpc1_1 gpc4102 (
      {stage2_25[88]},
      {stage3_25[34]}
   );
   gpc1_1 gpc4103 (
      {stage2_25[89]},
      {stage3_25[35]}
   );
   gpc1_1 gpc4104 (
      {stage2_25[90]},
      {stage3_25[36]}
   );
   gpc1_1 gpc4105 (
      {stage2_25[91]},
      {stage3_25[37]}
   );
   gpc1_1 gpc4106 (
      {stage2_25[92]},
      {stage3_25[38]}
   );
   gpc1_1 gpc4107 (
      {stage2_25[93]},
      {stage3_25[39]}
   );
   gpc1_1 gpc4108 (
      {stage2_25[94]},
      {stage3_25[40]}
   );
   gpc1_1 gpc4109 (
      {stage2_25[95]},
      {stage3_25[41]}
   );
   gpc1_1 gpc4110 (
      {stage2_25[96]},
      {stage3_25[42]}
   );
   gpc1_1 gpc4111 (
      {stage2_25[97]},
      {stage3_25[43]}
   );
   gpc1_1 gpc4112 (
      {stage2_25[98]},
      {stage3_25[44]}
   );
   gpc1_1 gpc4113 (
      {stage2_25[99]},
      {stage3_25[45]}
   );
   gpc1_1 gpc4114 (
      {stage2_25[100]},
      {stage3_25[46]}
   );
   gpc1_1 gpc4115 (
      {stage2_25[101]},
      {stage3_25[47]}
   );
   gpc1_1 gpc4116 (
      {stage2_25[102]},
      {stage3_25[48]}
   );
   gpc1_1 gpc4117 (
      {stage2_26[87]},
      {stage3_26[38]}
   );
   gpc1_1 gpc4118 (
      {stage2_26[88]},
      {stage3_26[39]}
   );
   gpc1_1 gpc4119 (
      {stage2_26[89]},
      {stage3_26[40]}
   );
   gpc1_1 gpc4120 (
      {stage2_26[90]},
      {stage3_26[41]}
   );
   gpc1_1 gpc4121 (
      {stage2_26[91]},
      {stage3_26[42]}
   );
   gpc1_1 gpc4122 (
      {stage2_26[92]},
      {stage3_26[43]}
   );
   gpc1_1 gpc4123 (
      {stage2_26[93]},
      {stage3_26[44]}
   );
   gpc1_1 gpc4124 (
      {stage2_26[94]},
      {stage3_26[45]}
   );
   gpc1_1 gpc4125 (
      {stage2_26[95]},
      {stage3_26[46]}
   );
   gpc1_1 gpc4126 (
      {stage2_26[96]},
      {stage3_26[47]}
   );
   gpc1_1 gpc4127 (
      {stage2_26[97]},
      {stage3_26[48]}
   );
   gpc1_1 gpc4128 (
      {stage2_26[98]},
      {stage3_26[49]}
   );
   gpc1_1 gpc4129 (
      {stage2_26[99]},
      {stage3_26[50]}
   );
   gpc1_1 gpc4130 (
      {stage2_27[72]},
      {stage3_27[42]}
   );
   gpc1_1 gpc4131 (
      {stage2_27[73]},
      {stage3_27[43]}
   );
   gpc1_1 gpc4132 (
      {stage2_27[74]},
      {stage3_27[44]}
   );
   gpc1_1 gpc4133 (
      {stage2_27[75]},
      {stage3_27[45]}
   );
   gpc1_1 gpc4134 (
      {stage2_27[76]},
      {stage3_27[46]}
   );
   gpc1_1 gpc4135 (
      {stage2_27[77]},
      {stage3_27[47]}
   );
   gpc1_1 gpc4136 (
      {stage2_27[78]},
      {stage3_27[48]}
   );
   gpc1_1 gpc4137 (
      {stage2_27[79]},
      {stage3_27[49]}
   );
   gpc1_1 gpc4138 (
      {stage2_27[80]},
      {stage3_27[50]}
   );
   gpc1_1 gpc4139 (
      {stage2_27[81]},
      {stage3_27[51]}
   );
   gpc1_1 gpc4140 (
      {stage2_27[82]},
      {stage3_27[52]}
   );
   gpc1_1 gpc4141 (
      {stage2_27[83]},
      {stage3_27[53]}
   );
   gpc1_1 gpc4142 (
      {stage2_27[84]},
      {stage3_27[54]}
   );
   gpc1_1 gpc4143 (
      {stage2_28[133]},
      {stage3_28[36]}
   );
   gpc1_1 gpc4144 (
      {stage2_28[134]},
      {stage3_28[37]}
   );
   gpc1_1 gpc4145 (
      {stage2_28[135]},
      {stage3_28[38]}
   );
   gpc1_1 gpc4146 (
      {stage2_28[136]},
      {stage3_28[39]}
   );
   gpc1_1 gpc4147 (
      {stage2_28[137]},
      {stage3_28[40]}
   );
   gpc1_1 gpc4148 (
      {stage2_28[138]},
      {stage3_28[41]}
   );
   gpc1_1 gpc4149 (
      {stage2_28[139]},
      {stage3_28[42]}
   );
   gpc1_1 gpc4150 (
      {stage2_28[140]},
      {stage3_28[43]}
   );
   gpc1_1 gpc4151 (
      {stage2_28[141]},
      {stage3_28[44]}
   );
   gpc1_1 gpc4152 (
      {stage2_28[142]},
      {stage3_28[45]}
   );
   gpc1_1 gpc4153 (
      {stage2_28[143]},
      {stage3_28[46]}
   );
   gpc1_1 gpc4154 (
      {stage2_28[144]},
      {stage3_28[47]}
   );
   gpc1_1 gpc4155 (
      {stage2_28[145]},
      {stage3_28[48]}
   );
   gpc1_1 gpc4156 (
      {stage2_28[146]},
      {stage3_28[49]}
   );
   gpc1_1 gpc4157 (
      {stage2_28[147]},
      {stage3_28[50]}
   );
   gpc1_1 gpc4158 (
      {stage2_28[148]},
      {stage3_28[51]}
   );
   gpc1_1 gpc4159 (
      {stage2_28[149]},
      {stage3_28[52]}
   );
   gpc1_1 gpc4160 (
      {stage2_28[150]},
      {stage3_28[53]}
   );
   gpc1_1 gpc4161 (
      {stage2_28[151]},
      {stage3_28[54]}
   );
   gpc1_1 gpc4162 (
      {stage2_28[152]},
      {stage3_28[55]}
   );
   gpc1_1 gpc4163 (
      {stage2_28[153]},
      {stage3_28[56]}
   );
   gpc1_1 gpc4164 (
      {stage2_28[154]},
      {stage3_28[57]}
   );
   gpc1_1 gpc4165 (
      {stage2_28[155]},
      {stage3_28[58]}
   );
   gpc1_1 gpc4166 (
      {stage2_28[156]},
      {stage3_28[59]}
   );
   gpc1_1 gpc4167 (
      {stage2_28[157]},
      {stage3_28[60]}
   );
   gpc1_1 gpc4168 (
      {stage2_28[158]},
      {stage3_28[61]}
   );
   gpc1_1 gpc4169 (
      {stage2_28[159]},
      {stage3_28[62]}
   );
   gpc1_1 gpc4170 (
      {stage2_28[160]},
      {stage3_28[63]}
   );
   gpc1_1 gpc4171 (
      {stage2_28[161]},
      {stage3_28[64]}
   );
   gpc1_1 gpc4172 (
      {stage2_28[162]},
      {stage3_28[65]}
   );
   gpc1_1 gpc4173 (
      {stage2_28[163]},
      {stage3_28[66]}
   );
   gpc1_1 gpc4174 (
      {stage2_28[164]},
      {stage3_28[67]}
   );
   gpc1_1 gpc4175 (
      {stage2_28[165]},
      {stage3_28[68]}
   );
   gpc1_1 gpc4176 (
      {stage2_28[166]},
      {stage3_28[69]}
   );
   gpc1_1 gpc4177 (
      {stage2_28[167]},
      {stage3_28[70]}
   );
   gpc1_1 gpc4178 (
      {stage2_28[168]},
      {stage3_28[71]}
   );
   gpc1_1 gpc4179 (
      {stage2_28[169]},
      {stage3_28[72]}
   );
   gpc1_1 gpc4180 (
      {stage2_28[170]},
      {stage3_28[73]}
   );
   gpc1_1 gpc4181 (
      {stage2_29[127]},
      {stage3_29[42]}
   );
   gpc1_1 gpc4182 (
      {stage2_29[128]},
      {stage3_29[43]}
   );
   gpc1_1 gpc4183 (
      {stage2_29[129]},
      {stage3_29[44]}
   );
   gpc1_1 gpc4184 (
      {stage2_29[130]},
      {stage3_29[45]}
   );
   gpc1_1 gpc4185 (
      {stage2_29[131]},
      {stage3_29[46]}
   );
   gpc1_1 gpc4186 (
      {stage2_29[132]},
      {stage3_29[47]}
   );
   gpc1_1 gpc4187 (
      {stage2_29[133]},
      {stage3_29[48]}
   );
   gpc1_1 gpc4188 (
      {stage2_29[134]},
      {stage3_29[49]}
   );
   gpc1_1 gpc4189 (
      {stage2_29[135]},
      {stage3_29[50]}
   );
   gpc1_1 gpc4190 (
      {stage2_29[136]},
      {stage3_29[51]}
   );
   gpc1_1 gpc4191 (
      {stage2_29[137]},
      {stage3_29[52]}
   );
   gpc1_1 gpc4192 (
      {stage2_29[138]},
      {stage3_29[53]}
   );
   gpc1_1 gpc4193 (
      {stage2_29[139]},
      {stage3_29[54]}
   );
   gpc1_1 gpc4194 (
      {stage2_29[140]},
      {stage3_29[55]}
   );
   gpc1_1 gpc4195 (
      {stage2_29[141]},
      {stage3_29[56]}
   );
   gpc1_1 gpc4196 (
      {stage2_29[142]},
      {stage3_29[57]}
   );
   gpc1_1 gpc4197 (
      {stage2_30[66]},
      {stage3_30[45]}
   );
   gpc1_1 gpc4198 (
      {stage2_30[67]},
      {stage3_30[46]}
   );
   gpc1_1 gpc4199 (
      {stage2_30[68]},
      {stage3_30[47]}
   );
   gpc1_1 gpc4200 (
      {stage2_30[69]},
      {stage3_30[48]}
   );
   gpc1_1 gpc4201 (
      {stage2_30[70]},
      {stage3_30[49]}
   );
   gpc1_1 gpc4202 (
      {stage2_30[71]},
      {stage3_30[50]}
   );
   gpc1_1 gpc4203 (
      {stage2_30[72]},
      {stage3_30[51]}
   );
   gpc1_1 gpc4204 (
      {stage2_30[73]},
      {stage3_30[52]}
   );
   gpc1_1 gpc4205 (
      {stage2_30[74]},
      {stage3_30[53]}
   );
   gpc1_1 gpc4206 (
      {stage2_30[75]},
      {stage3_30[54]}
   );
   gpc1_1 gpc4207 (
      {stage2_30[76]},
      {stage3_30[55]}
   );
   gpc1_1 gpc4208 (
      {stage2_30[77]},
      {stage3_30[56]}
   );
   gpc1_1 gpc4209 (
      {stage2_30[78]},
      {stage3_30[57]}
   );
   gpc1_1 gpc4210 (
      {stage2_30[79]},
      {stage3_30[58]}
   );
   gpc1_1 gpc4211 (
      {stage2_30[80]},
      {stage3_30[59]}
   );
   gpc1_1 gpc4212 (
      {stage2_30[81]},
      {stage3_30[60]}
   );
   gpc1_1 gpc4213 (
      {stage2_30[82]},
      {stage3_30[61]}
   );
   gpc1_1 gpc4214 (
      {stage2_30[83]},
      {stage3_30[62]}
   );
   gpc1_1 gpc4215 (
      {stage2_30[84]},
      {stage3_30[63]}
   );
   gpc1_1 gpc4216 (
      {stage2_30[85]},
      {stage3_30[64]}
   );
   gpc1_1 gpc4217 (
      {stage2_30[86]},
      {stage3_30[65]}
   );
   gpc1_1 gpc4218 (
      {stage2_30[87]},
      {stage3_30[66]}
   );
   gpc1_1 gpc4219 (
      {stage2_30[88]},
      {stage3_30[67]}
   );
   gpc1_1 gpc4220 (
      {stage2_30[89]},
      {stage3_30[68]}
   );
   gpc1_1 gpc4221 (
      {stage2_30[90]},
      {stage3_30[69]}
   );
   gpc1_1 gpc4222 (
      {stage2_30[91]},
      {stage3_30[70]}
   );
   gpc1_1 gpc4223 (
      {stage2_31[83]},
      {stage3_31[39]}
   );
   gpc1_1 gpc4224 (
      {stage2_31[84]},
      {stage3_31[40]}
   );
   gpc1_1 gpc4225 (
      {stage2_31[85]},
      {stage3_31[41]}
   );
   gpc1_1 gpc4226 (
      {stage2_31[86]},
      {stage3_31[42]}
   );
   gpc1_1 gpc4227 (
      {stage2_31[87]},
      {stage3_31[43]}
   );
   gpc1_1 gpc4228 (
      {stage2_31[88]},
      {stage3_31[44]}
   );
   gpc1_1 gpc4229 (
      {stage2_31[89]},
      {stage3_31[45]}
   );
   gpc1_1 gpc4230 (
      {stage2_31[90]},
      {stage3_31[46]}
   );
   gpc1_1 gpc4231 (
      {stage2_31[91]},
      {stage3_31[47]}
   );
   gpc1_1 gpc4232 (
      {stage2_31[92]},
      {stage3_31[48]}
   );
   gpc1_1 gpc4233 (
      {stage2_31[93]},
      {stage3_31[49]}
   );
   gpc1_1 gpc4234 (
      {stage2_31[94]},
      {stage3_31[50]}
   );
   gpc1_1 gpc4235 (
      {stage2_31[95]},
      {stage3_31[51]}
   );
   gpc1_1 gpc4236 (
      {stage2_31[96]},
      {stage3_31[52]}
   );
   gpc1_1 gpc4237 (
      {stage2_31[97]},
      {stage3_31[53]}
   );
   gpc1_1 gpc4238 (
      {stage2_31[98]},
      {stage3_31[54]}
   );
   gpc1_1 gpc4239 (
      {stage2_31[99]},
      {stage3_31[55]}
   );
   gpc1_1 gpc4240 (
      {stage2_31[100]},
      {stage3_31[56]}
   );
   gpc1_1 gpc4241 (
      {stage2_31[101]},
      {stage3_31[57]}
   );
   gpc1_1 gpc4242 (
      {stage2_32[46]},
      {stage3_32[30]}
   );
   gpc1_1 gpc4243 (
      {stage2_32[47]},
      {stage3_32[31]}
   );
   gpc1_1 gpc4244 (
      {stage2_32[48]},
      {stage3_32[32]}
   );
   gpc1_1 gpc4245 (
      {stage2_32[49]},
      {stage3_32[33]}
   );
   gpc1_1 gpc4246 (
      {stage2_32[50]},
      {stage3_32[34]}
   );
   gpc1_1 gpc4247 (
      {stage2_32[51]},
      {stage3_32[35]}
   );
   gpc1_1 gpc4248 (
      {stage2_32[52]},
      {stage3_32[36]}
   );
   gpc1_1 gpc4249 (
      {stage2_32[53]},
      {stage3_32[37]}
   );
   gpc1_1 gpc4250 (
      {stage2_32[54]},
      {stage3_32[38]}
   );
   gpc1_1 gpc4251 (
      {stage2_32[55]},
      {stage3_32[39]}
   );
   gpc1_1 gpc4252 (
      {stage2_32[56]},
      {stage3_32[40]}
   );
   gpc1_1 gpc4253 (
      {stage2_32[57]},
      {stage3_32[41]}
   );
   gpc1_1 gpc4254 (
      {stage2_32[58]},
      {stage3_32[42]}
   );
   gpc1_1 gpc4255 (
      {stage2_32[59]},
      {stage3_32[43]}
   );
   gpc1_1 gpc4256 (
      {stage2_32[60]},
      {stage3_32[44]}
   );
   gpc1_1 gpc4257 (
      {stage2_32[61]},
      {stage3_32[45]}
   );
   gpc1_1 gpc4258 (
      {stage2_32[62]},
      {stage3_32[46]}
   );
   gpc1_1 gpc4259 (
      {stage2_32[63]},
      {stage3_32[47]}
   );
   gpc1_1 gpc4260 (
      {stage2_32[64]},
      {stage3_32[48]}
   );
   gpc1_1 gpc4261 (
      {stage2_32[65]},
      {stage3_32[49]}
   );
   gpc1_1 gpc4262 (
      {stage2_32[66]},
      {stage3_32[50]}
   );
   gpc1_1 gpc4263 (
      {stage2_32[67]},
      {stage3_32[51]}
   );
   gpc1_1 gpc4264 (
      {stage2_32[68]},
      {stage3_32[52]}
   );
   gpc1_1 gpc4265 (
      {stage2_32[69]},
      {stage3_32[53]}
   );
   gpc1_1 gpc4266 (
      {stage2_32[70]},
      {stage3_32[54]}
   );
   gpc1_1 gpc4267 (
      {stage2_32[71]},
      {stage3_32[55]}
   );
   gpc1_1 gpc4268 (
      {stage2_32[72]},
      {stage3_32[56]}
   );
   gpc1_1 gpc4269 (
      {stage2_32[73]},
      {stage3_32[57]}
   );
   gpc1_1 gpc4270 (
      {stage2_33[57]},
      {stage3_33[24]}
   );
   gpc1_1 gpc4271 (
      {stage2_33[58]},
      {stage3_33[25]}
   );
   gpc1_1 gpc4272 (
      {stage2_33[59]},
      {stage3_33[26]}
   );
   gpc1_1 gpc4273 (
      {stage2_34[24]},
      {stage3_34[16]}
   );
   gpc1_1 gpc4274 (
      {stage2_34[25]},
      {stage3_34[17]}
   );
   gpc1_1 gpc4275 (
      {stage2_34[26]},
      {stage3_34[18]}
   );
   gpc1_1 gpc4276 (
      {stage2_34[27]},
      {stage3_34[19]}
   );
   gpc1_1 gpc4277 (
      {stage2_34[28]},
      {stage3_34[20]}
   );
   gpc1_1 gpc4278 (
      {stage2_34[29]},
      {stage3_34[21]}
   );
   gpc1_1 gpc4279 (
      {stage2_34[30]},
      {stage3_34[22]}
   );
   gpc1_1 gpc4280 (
      {stage2_34[31]},
      {stage3_34[23]}
   );
   gpc1_1 gpc4281 (
      {stage2_34[32]},
      {stage3_34[24]}
   );
   gpc1_1 gpc4282 (
      {stage2_34[33]},
      {stage3_34[25]}
   );
   gpc1_1 gpc4283 (
      {stage2_34[34]},
      {stage3_34[26]}
   );
   gpc606_5 gpc4284 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc4285 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc4286 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc4287 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc4288 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[4],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc4289 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[5],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc4290 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27], stage3_4[28], stage3_4[29]},
      {stage4_6[4],stage4_5[6],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc606_5 gpc4291 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[5],stage4_5[7]}
   );
   gpc606_5 gpc4292 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[1],stage4_7[1],stage4_6[6],stage4_5[8]}
   );
   gpc606_5 gpc4293 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[2],stage4_7[2],stage4_6[7],stage4_5[9]}
   );
   gpc606_5 gpc4294 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[3],stage4_7[3],stage4_6[8],stage4_5[10]}
   );
   gpc615_5 gpc4295 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[24]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[4],stage4_8[4],stage4_7[4],stage4_6[9]}
   );
   gpc615_5 gpc4296 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[25]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[5],stage4_8[5],stage4_7[5],stage4_6[10]}
   );
   gpc615_5 gpc4297 (
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14]},
      {stage3_7[26]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[6],stage4_8[6],stage4_7[6],stage4_6[11]}
   );
   gpc615_5 gpc4298 (
      {stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18], stage3_6[19]},
      {stage3_7[27]},
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22], stage3_8[23]},
      {stage4_10[3],stage4_9[7],stage4_8[7],stage4_7[7],stage4_6[12]}
   );
   gpc615_5 gpc4299 (
      {stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23], stage3_6[24]},
      {stage3_7[28]},
      {stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28], stage3_8[29]},
      {stage4_10[4],stage4_9[8],stage4_8[8],stage4_7[8],stage4_6[13]}
   );
   gpc615_5 gpc4300 (
      {stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage3_7[29]},
      {stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34], stage3_8[35]},
      {stage4_10[5],stage4_9[9],stage4_8[9],stage4_7[9],stage4_6[14]}
   );
   gpc615_5 gpc4301 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[36]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[6],stage4_9[10],stage4_8[10],stage4_7[10]}
   );
   gpc615_5 gpc4302 (
      {stage3_7[35], stage3_7[36], stage3_7[37], stage3_7[38], stage3_7[39]},
      {stage3_8[37]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[7],stage4_9[11],stage4_8[11],stage4_7[11]}
   );
   gpc615_5 gpc4303 (
      {stage3_7[40], stage3_7[41], stage3_7[42], stage3_7[43], stage3_7[44]},
      {stage3_8[38]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[8],stage4_9[12],stage4_8[12],stage4_7[12]}
   );
   gpc117_4 gpc4304 (
      {stage3_8[39], stage3_8[40], stage3_8[41], stage3_8[42], stage3_8[43], stage3_8[44], stage3_8[45]},
      {stage3_9[18]},
      {stage3_10[0]},
      {stage4_11[3],stage4_10[9],stage4_9[13],stage4_8[13]}
   );
   gpc117_4 gpc4305 (
      {stage3_8[46], stage3_8[47], stage3_8[48], stage3_8[49], stage3_8[50], stage3_8[51], stage3_8[52]},
      {stage3_9[19]},
      {stage3_10[1]},
      {stage4_11[4],stage4_10[10],stage4_9[14],stage4_8[14]}
   );
   gpc606_5 gpc4306 (
      {stage3_8[53], stage3_8[54], stage3_8[55], stage3_8[56], stage3_8[57], stage3_8[58]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[0],stage4_11[5],stage4_10[11],stage4_9[15],stage4_8[15]}
   );
   gpc606_5 gpc4307 (
      {stage3_8[59], stage3_8[60], stage3_8[61], stage3_8[62], stage3_8[63], stage3_8[64]},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[6],stage4_10[12],stage4_9[16],stage4_8[16]}
   );
   gpc615_5 gpc4308 (
      {stage3_8[65], stage3_8[66], stage3_8[67], stage3_8[68], stage3_8[69]},
      {stage3_9[20]},
      {stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage4_12[2],stage4_11[7],stage4_10[13],stage4_9[17],stage4_8[17]}
   );
   gpc615_5 gpc4309 (
      {stage3_8[70], stage3_8[71], stage3_8[72], stage3_8[73], stage3_8[74]},
      {stage3_9[21]},
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage4_12[3],stage4_11[8],stage4_10[14],stage4_9[18],stage4_8[18]}
   );
   gpc615_5 gpc4310 (
      {stage3_8[75], stage3_8[76], stage3_8[77], stage3_8[78], stage3_8[79]},
      {stage3_9[22]},
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage4_12[4],stage4_11[9],stage4_10[15],stage4_9[19],stage4_8[19]}
   );
   gpc615_5 gpc4311 (
      {stage3_8[80], stage3_8[81], stage3_8[82], stage3_8[83], stage3_8[84]},
      {stage3_9[23]},
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage4_12[5],stage4_11[10],stage4_10[16],stage4_9[20],stage4_8[20]}
   );
   gpc606_5 gpc4312 (
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[6],stage4_11[11],stage4_10[17],stage4_9[21]}
   );
   gpc1163_5 gpc4313 (
      {stage3_11[6], stage3_11[7], stage3_11[8]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[7],stage4_11[12]}
   );
   gpc1163_5 gpc4314 (
      {stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_13[1]},
      {stage3_14[1]},
      {stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[8],stage4_11[13]}
   );
   gpc1163_5 gpc4315 (
      {stage3_11[12], stage3_11[13], stage3_11[14]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_13[2]},
      {stage3_14[2]},
      {stage4_15[2],stage4_14[2],stage4_13[3],stage4_12[9],stage4_11[14]}
   );
   gpc1163_5 gpc4316 (
      {stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_13[3]},
      {stage3_14[3]},
      {stage4_15[3],stage4_14[3],stage4_13[4],stage4_12[10],stage4_11[15]}
   );
   gpc1163_5 gpc4317 (
      {stage3_11[18], stage3_11[19], stage3_11[20]},
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_13[4]},
      {stage3_14[4]},
      {stage4_15[4],stage4_14[4],stage4_13[5],stage4_12[11],stage4_11[16]}
   );
   gpc615_5 gpc4318 (
      {stage3_11[21], stage3_11[22], stage3_11[23], stage3_11[24], stage3_11[25]},
      {stage3_12[30]},
      {stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage4_15[5],stage4_14[5],stage4_13[6],stage4_12[12],stage4_11[17]}
   );
   gpc615_5 gpc4319 (
      {stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29], stage3_11[30]},
      {stage3_12[31]},
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16]},
      {stage4_15[6],stage4_14[6],stage4_13[7],stage4_12[13],stage4_11[18]}
   );
   gpc606_5 gpc4320 (
      {stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35], stage3_12[36], stage3_12[37]},
      {stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10]},
      {stage4_16[0],stage4_15[7],stage4_14[7],stage4_13[8],stage4_12[14]}
   );
   gpc606_5 gpc4321 (
      {stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[8],stage4_14[8],stage4_13[9]}
   );
   gpc606_5 gpc4322 (
      {stage3_13[23], stage3_13[24], stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[9],stage4_14[9],stage4_13[10]}
   );
   gpc615_5 gpc4323 (
      {stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15]},
      {stage3_15[12]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[10],stage4_14[10]}
   );
   gpc615_5 gpc4324 (
      {stage3_14[16], stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20]},
      {stage3_15[13]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[11],stage4_14[11]}
   );
   gpc615_5 gpc4325 (
      {stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24], stage3_14[25]},
      {stage3_15[14]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[12],stage4_14[12]}
   );
   gpc615_5 gpc4326 (
      {stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[15]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[13],stage4_14[13]}
   );
   gpc615_5 gpc4327 (
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35]},
      {stage3_15[16]},
      {stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29]},
      {stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[14],stage4_14[14]}
   );
   gpc1163_5 gpc4328 (
      {stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[5],stage4_17[7],stage4_16[8],stage4_15[15]}
   );
   gpc615_5 gpc4329 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[36]},
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6]},
      {stage4_19[1],stage4_18[6],stage4_17[8],stage4_16[9],stage4_15[16]}
   );
   gpc615_5 gpc4330 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[37]},
      {stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11], stage3_17[12]},
      {stage4_19[2],stage4_18[7],stage4_17[9],stage4_16[10],stage4_15[17]}
   );
   gpc615_5 gpc4331 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[38]},
      {stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17], stage3_17[18]},
      {stage4_19[3],stage4_18[8],stage4_17[10],stage4_16[11],stage4_15[18]}
   );
   gpc615_5 gpc4332 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[39]},
      {stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23], stage3_17[24]},
      {stage4_19[4],stage4_18[9],stage4_17[11],stage4_16[12],stage4_15[19]}
   );
   gpc615_5 gpc4333 (
      {stage3_15[40], stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44]},
      {stage3_16[40]},
      {stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29], stage3_17[30]},
      {stage4_19[5],stage4_18[10],stage4_17[12],stage4_16[13],stage4_15[20]}
   );
   gpc615_5 gpc4334 (
      {stage3_15[45], stage3_15[46], stage3_15[47], stage3_15[48], stage3_15[49]},
      {stage3_16[41]},
      {stage3_17[31], stage3_17[32], stage3_17[33], stage3_17[34], stage3_17[35], stage3_17[36]},
      {stage4_19[6],stage4_18[11],stage4_17[13],stage4_16[14],stage4_15[21]}
   );
   gpc615_5 gpc4335 (
      {stage3_15[50], stage3_15[51], stage3_15[52], stage3_15[53], stage3_15[54]},
      {stage3_16[42]},
      {stage3_17[37], stage3_17[38], stage3_17[39], stage3_17[40], stage3_17[41], stage3_17[42]},
      {stage4_19[7],stage4_18[12],stage4_17[14],stage4_16[15],stage4_15[22]}
   );
   gpc606_5 gpc4336 (
      {stage3_16[43], stage3_16[44], stage3_16[45], stage3_16[46], stage3_16[47], stage3_16[48]},
      {stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5], stage3_18[6]},
      {stage4_20[0],stage4_19[8],stage4_18[13],stage4_17[15],stage4_16[16]}
   );
   gpc606_5 gpc4337 (
      {stage3_16[49], stage3_16[50], stage3_16[51], stage3_16[52], stage3_16[53], stage3_16[54]},
      {stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage4_20[1],stage4_19[9],stage4_18[14],stage4_17[16],stage4_16[17]}
   );
   gpc606_5 gpc4338 (
      {stage3_16[55], stage3_16[56], stage3_16[57], stage3_16[58], stage3_16[59], stage3_16[60]},
      {stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17], stage3_18[18]},
      {stage4_20[2],stage4_19[10],stage4_18[15],stage4_17[17],stage4_16[18]}
   );
   gpc606_5 gpc4339 (
      {stage3_16[61], stage3_16[62], stage3_16[63], stage3_16[64], stage3_16[65], stage3_16[66]},
      {stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24]},
      {stage4_20[3],stage4_19[11],stage4_18[16],stage4_17[18],stage4_16[19]}
   );
   gpc606_5 gpc4340 (
      {stage3_17[43], stage3_17[44], stage3_17[45], stage3_17[46], stage3_17[47], stage3_17[48]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[4],stage4_19[12],stage4_18[17],stage4_17[19]}
   );
   gpc606_5 gpc4341 (
      {stage3_17[49], stage3_17[50], stage3_17[51], stage3_17[52], stage3_17[53], stage3_17[54]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[5],stage4_19[13],stage4_18[18],stage4_17[20]}
   );
   gpc615_5 gpc4342 (
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16]},
      {stage3_20[0]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[2],stage4_20[6],stage4_19[14]}
   );
   gpc615_5 gpc4343 (
      {stage3_19[17], stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21]},
      {stage3_20[1]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[3],stage4_20[7],stage4_19[15]}
   );
   gpc615_5 gpc4344 (
      {stage3_19[22], stage3_19[23], stage3_19[24], stage3_19[25], stage3_19[26]},
      {stage3_20[2]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[4],stage4_20[8],stage4_19[16]}
   );
   gpc615_5 gpc4345 (
      {stage3_19[27], stage3_19[28], stage3_19[29], stage3_19[30], stage3_19[31]},
      {stage3_20[3]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[3],stage4_21[5],stage4_20[9],stage4_19[17]}
   );
   gpc615_5 gpc4346 (
      {stage3_19[32], stage3_19[33], stage3_19[34], stage3_19[35], stage3_19[36]},
      {stage3_20[4]},
      {stage3_21[24], stage3_21[25], stage3_21[26], stage3_21[27], stage3_21[28], stage3_21[29]},
      {stage4_23[4],stage4_22[4],stage4_21[6],stage4_20[10],stage4_19[18]}
   );
   gpc615_5 gpc4347 (
      {stage3_19[37], stage3_19[38], stage3_19[39], stage3_19[40], stage3_19[41]},
      {stage3_20[5]},
      {stage3_21[30], stage3_21[31], stage3_21[32], stage3_21[33], stage3_21[34], stage3_21[35]},
      {stage4_23[5],stage4_22[5],stage4_21[7],stage4_20[11],stage4_19[19]}
   );
   gpc615_5 gpc4348 (
      {stage3_19[42], stage3_19[43], stage3_19[44], stage3_19[45], stage3_19[46]},
      {stage3_20[6]},
      {stage3_21[36], stage3_21[37], stage3_21[38], stage3_21[39], stage3_21[40], stage3_21[41]},
      {stage4_23[6],stage4_22[6],stage4_21[8],stage4_20[12],stage4_19[20]}
   );
   gpc615_5 gpc4349 (
      {stage3_19[47], stage3_19[48], stage3_19[49], stage3_19[50], stage3_19[51]},
      {stage3_20[7]},
      {stage3_21[42], stage3_21[43], stage3_21[44], stage3_21[45], stage3_21[46], stage3_21[47]},
      {stage4_23[7],stage4_22[7],stage4_21[9],stage4_20[13],stage4_19[21]}
   );
   gpc1325_5 gpc4350 (
      {stage3_19[52], stage3_19[53], stage3_19[54], stage3_19[55], stage3_19[56]},
      {stage3_20[8], stage3_20[9]},
      {stage3_21[48], stage3_21[49], stage3_21[50]},
      {stage3_22[0]},
      {stage4_23[8],stage4_22[8],stage4_21[10],stage4_20[14],stage4_19[22]}
   );
   gpc1325_5 gpc4351 (
      {stage3_19[57], stage3_19[58], stage3_19[59], stage3_19[60], stage3_19[61]},
      {stage3_20[10], stage3_20[11]},
      {stage3_21[51], stage3_21[52], stage3_21[53]},
      {stage3_22[1]},
      {stage4_23[9],stage4_22[9],stage4_21[11],stage4_20[15],stage4_19[23]}
   );
   gpc606_5 gpc4352 (
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6], stage3_22[7]},
      {stage4_24[0],stage4_23[10],stage4_22[10],stage4_21[12],stage4_20[16]}
   );
   gpc606_5 gpc4353 (
      {stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23]},
      {stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11], stage3_22[12], stage3_22[13]},
      {stage4_24[1],stage4_23[11],stage4_22[11],stage4_21[13],stage4_20[17]}
   );
   gpc606_5 gpc4354 (
      {stage3_20[24], stage3_20[25], stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29]},
      {stage3_22[14], stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage4_24[2],stage4_23[12],stage4_22[12],stage4_21[14],stage4_20[18]}
   );
   gpc606_5 gpc4355 (
      {stage3_21[54], stage3_21[55], stage3_21[56], stage3_21[57], stage3_21[58], stage3_21[59]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[3],stage4_23[13],stage4_22[13],stage4_21[15]}
   );
   gpc207_4 gpc4356 (
      {stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24], stage3_22[25], stage3_22[26]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[1],stage4_24[4],stage4_23[14],stage4_22[14]}
   );
   gpc615_5 gpc4357 (
      {stage3_22[27], stage3_22[28], stage3_22[29], stage3_22[30], stage3_22[31]},
      {stage3_23[6]},
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7]},
      {stage4_26[0],stage4_25[2],stage4_24[5],stage4_23[15],stage4_22[15]}
   );
   gpc615_5 gpc4358 (
      {stage3_22[32], stage3_22[33], stage3_22[34], stage3_22[35], stage3_22[36]},
      {stage3_23[7]},
      {stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11], stage3_24[12], stage3_24[13]},
      {stage4_26[1],stage4_25[3],stage4_24[6],stage4_23[16],stage4_22[16]}
   );
   gpc606_5 gpc4359 (
      {stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12], stage3_23[13]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[4],stage4_24[7],stage4_23[17]}
   );
   gpc615_5 gpc4360 (
      {stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17], stage3_23[18]},
      {stage3_24[14]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[5],stage4_24[8],stage4_23[18]}
   );
   gpc615_5 gpc4361 (
      {stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23]},
      {stage3_24[15]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[4],stage4_25[6],stage4_24[9],stage4_23[19]}
   );
   gpc615_5 gpc4362 (
      {stage3_23[24], stage3_23[25], stage3_23[26], stage3_23[27], stage3_23[28]},
      {stage3_24[16]},
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage4_27[3],stage4_26[5],stage4_25[7],stage4_24[10],stage4_23[20]}
   );
   gpc606_5 gpc4363 (
      {stage3_24[17], stage3_24[18], stage3_24[19], stage3_24[20], stage3_24[21], stage3_24[22]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[4],stage4_26[6],stage4_25[8],stage4_24[11]}
   );
   gpc606_5 gpc4364 (
      {stage3_24[23], stage3_24[24], stage3_24[25], stage3_24[26], stage3_24[27], stage3_24[28]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[1],stage4_27[5],stage4_26[7],stage4_25[9],stage4_24[12]}
   );
   gpc606_5 gpc4365 (
      {stage3_24[29], stage3_24[30], stage3_24[31], stage3_24[32], stage3_24[33], stage3_24[34]},
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage4_28[2],stage4_27[6],stage4_26[8],stage4_25[10],stage4_24[13]}
   );
   gpc606_5 gpc4366 (
      {stage3_24[35], stage3_24[36], stage3_24[37], stage3_24[38], stage3_24[39], stage3_24[40]},
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage4_28[3],stage4_27[7],stage4_26[9],stage4_25[11],stage4_24[14]}
   );
   gpc606_5 gpc4367 (
      {stage3_24[41], stage3_24[42], stage3_24[43], stage3_24[44], stage3_24[45], stage3_24[46]},
      {stage3_26[24], stage3_26[25], stage3_26[26], stage3_26[27], stage3_26[28], stage3_26[29]},
      {stage4_28[4],stage4_27[8],stage4_26[10],stage4_25[12],stage4_24[15]}
   );
   gpc606_5 gpc4368 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28], stage3_25[29]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[5],stage4_27[9],stage4_26[11],stage4_25[13]}
   );
   gpc606_5 gpc4369 (
      {stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33], stage3_25[34], stage3_25[35]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[6],stage4_27[10],stage4_26[12],stage4_25[14]}
   );
   gpc606_5 gpc4370 (
      {stage3_25[36], stage3_25[37], stage3_25[38], stage3_25[39], stage3_25[40], stage3_25[41]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[7],stage4_27[11],stage4_26[13],stage4_25[15]}
   );
   gpc615_5 gpc4371 (
      {stage3_25[42], stage3_25[43], stage3_25[44], stage3_25[45], stage3_25[46]},
      {stage3_26[30]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[8],stage4_27[12],stage4_26[14],stage4_25[16]}
   );
   gpc615_5 gpc4372 (
      {stage3_26[31], stage3_26[32], stage3_26[33], stage3_26[34], stage3_26[35]},
      {stage3_27[24]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[4],stage4_28[9],stage4_27[13],stage4_26[15]}
   );
   gpc615_5 gpc4373 (
      {stage3_26[36], stage3_26[37], stage3_26[38], stage3_26[39], stage3_26[40]},
      {stage3_27[25]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage4_30[1],stage4_29[5],stage4_28[10],stage4_27[14],stage4_26[16]}
   );
   gpc615_5 gpc4374 (
      {stage3_26[41], stage3_26[42], stage3_26[43], stage3_26[44], stage3_26[45]},
      {stage3_27[26]},
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17]},
      {stage4_30[2],stage4_29[6],stage4_28[11],stage4_27[15],stage4_26[17]}
   );
   gpc606_5 gpc4375 (
      {stage3_27[27], stage3_27[28], stage3_27[29], stage3_27[30], stage3_27[31], stage3_27[32]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[3],stage4_29[7],stage4_28[12],stage4_27[16]}
   );
   gpc615_5 gpc4376 (
      {stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36], stage3_27[37]},
      {stage3_28[18]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[4],stage4_29[8],stage4_28[13],stage4_27[17]}
   );
   gpc615_5 gpc4377 (
      {stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41], stage3_27[42]},
      {stage3_28[19]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[5],stage4_29[9],stage4_28[14],stage4_27[18]}
   );
   gpc615_5 gpc4378 (
      {stage3_27[43], stage3_27[44], stage3_27[45], stage3_27[46], stage3_27[47]},
      {stage3_28[20]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[6],stage4_29[10],stage4_28[15],stage4_27[19]}
   );
   gpc606_5 gpc4379 (
      {stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[4],stage4_30[7],stage4_29[11],stage4_28[16]}
   );
   gpc606_5 gpc4380 (
      {stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30], stage3_28[31], stage3_28[32]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[5],stage4_30[8],stage4_29[12],stage4_28[17]}
   );
   gpc606_5 gpc4381 (
      {stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36], stage3_28[37], stage3_28[38]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[6],stage4_30[9],stage4_29[13],stage4_28[18]}
   );
   gpc606_5 gpc4382 (
      {stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42], stage3_28[43], stage3_28[44]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[7],stage4_30[10],stage4_29[14],stage4_28[19]}
   );
   gpc606_5 gpc4383 (
      {stage3_28[45], stage3_28[46], stage3_28[47], stage3_28[48], stage3_28[49], stage3_28[50]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage4_32[4],stage4_31[8],stage4_30[11],stage4_29[15],stage4_28[20]}
   );
   gpc606_5 gpc4384 (
      {stage3_28[51], stage3_28[52], stage3_28[53], stage3_28[54], stage3_28[55], stage3_28[56]},
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage4_32[5],stage4_31[9],stage4_30[12],stage4_29[16],stage4_28[21]}
   );
   gpc606_5 gpc4385 (
      {stage3_28[57], stage3_28[58], stage3_28[59], stage3_28[60], stage3_28[61], stage3_28[62]},
      {stage3_30[36], stage3_30[37], stage3_30[38], stage3_30[39], stage3_30[40], stage3_30[41]},
      {stage4_32[6],stage4_31[10],stage4_30[13],stage4_29[17],stage4_28[22]}
   );
   gpc606_5 gpc4386 (
      {stage3_28[63], stage3_28[64], stage3_28[65], stage3_28[66], stage3_28[67], stage3_28[68]},
      {stage3_30[42], stage3_30[43], stage3_30[44], stage3_30[45], stage3_30[46], stage3_30[47]},
      {stage4_32[7],stage4_31[11],stage4_30[14],stage4_29[18],stage4_28[23]}
   );
   gpc606_5 gpc4387 (
      {stage3_28[69], stage3_28[70], stage3_28[71], stage3_28[72], stage3_28[73], 1'b0},
      {stage3_30[48], stage3_30[49], stage3_30[50], stage3_30[51], stage3_30[52], stage3_30[53]},
      {stage4_32[8],stage4_31[12],stage4_30[15],stage4_29[19],stage4_28[24]}
   );
   gpc606_5 gpc4388 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[9],stage4_31[13],stage4_30[16],stage4_29[20]}
   );
   gpc606_5 gpc4389 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], stage3_29[35]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[10],stage4_31[14],stage4_30[17],stage4_29[21]}
   );
   gpc606_5 gpc4390 (
      {stage3_29[36], stage3_29[37], stage3_29[38], stage3_29[39], stage3_29[40], stage3_29[41]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[11],stage4_31[15],stage4_30[18],stage4_29[22]}
   );
   gpc606_5 gpc4391 (
      {stage3_29[42], stage3_29[43], stage3_29[44], stage3_29[45], stage3_29[46], stage3_29[47]},
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23]},
      {stage4_33[3],stage4_32[12],stage4_31[16],stage4_30[19],stage4_29[23]}
   );
   gpc615_5 gpc4392 (
      {stage3_29[48], stage3_29[49], stage3_29[50], stage3_29[51], stage3_29[52]},
      {stage3_30[54]},
      {stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage4_33[4],stage4_32[13],stage4_31[17],stage4_30[20],stage4_29[24]}
   );
   gpc615_5 gpc4393 (
      {stage3_29[53], stage3_29[54], stage3_29[55], stage3_29[56], stage3_29[57]},
      {stage3_30[55]},
      {stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33], stage3_31[34], stage3_31[35]},
      {stage4_33[5],stage4_32[14],stage4_31[18],stage4_30[21],stage4_29[25]}
   );
   gpc606_5 gpc4394 (
      {stage3_30[56], stage3_30[57], stage3_30[58], stage3_30[59], stage3_30[60], stage3_30[61]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[6],stage4_32[15],stage4_31[19],stage4_30[22]}
   );
   gpc606_5 gpc4395 (
      {stage3_30[62], stage3_30[63], stage3_30[64], stage3_30[65], stage3_30[66], stage3_30[67]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[7],stage4_32[16],stage4_31[20],stage4_30[23]}
   );
   gpc615_5 gpc4396 (
      {stage3_31[36], stage3_31[37], stage3_31[38], stage3_31[39], stage3_31[40]},
      {stage3_32[12]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[8],stage4_32[17],stage4_31[21]}
   );
   gpc615_5 gpc4397 (
      {stage3_31[41], stage3_31[42], stage3_31[43], stage3_31[44], stage3_31[45]},
      {stage3_32[13]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[3],stage4_33[9],stage4_32[18],stage4_31[22]}
   );
   gpc615_5 gpc4398 (
      {stage3_31[46], stage3_31[47], stage3_31[48], stage3_31[49], stage3_31[50]},
      {stage3_32[14]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[4],stage4_33[10],stage4_32[19],stage4_31[23]}
   );
   gpc606_5 gpc4399 (
      {stage3_32[15], stage3_32[16], stage3_32[17], stage3_32[18], stage3_32[19], stage3_32[20]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[3],stage4_34[5],stage4_33[11],stage4_32[20]}
   );
   gpc606_5 gpc4400 (
      {stage3_32[21], stage3_32[22], stage3_32[23], stage3_32[24], stage3_32[25], stage3_32[26]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[4],stage4_34[6],stage4_33[12],stage4_32[21]}
   );
   gpc606_5 gpc4401 (
      {stage3_32[27], stage3_32[28], stage3_32[29], stage3_32[30], stage3_32[31], stage3_32[32]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[5],stage4_34[7],stage4_33[13],stage4_32[22]}
   );
   gpc606_5 gpc4402 (
      {stage3_32[33], stage3_32[34], stage3_32[35], stage3_32[36], stage3_32[37], stage3_32[38]},
      {stage3_34[18], stage3_34[19], stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23]},
      {stage4_36[3],stage4_35[6],stage4_34[8],stage4_33[14],stage4_32[23]}
   );
   gpc606_5 gpc4403 (
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[4],stage4_35[7],stage4_34[9],stage4_33[15]}
   );
   gpc1_1 gpc4404 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc4405 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc4406 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4407 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc4408 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc4409 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc4410 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc4411 (
      {stage3_0[7]},
      {stage4_0[7]}
   );
   gpc1_1 gpc4412 (
      {stage3_0[8]},
      {stage4_0[8]}
   );
   gpc1_1 gpc4413 (
      {stage3_0[9]},
      {stage4_0[9]}
   );
   gpc1_1 gpc4414 (
      {stage3_0[10]},
      {stage4_0[10]}
   );
   gpc1_1 gpc4415 (
      {stage3_1[12]},
      {stage4_1[2]}
   );
   gpc1_1 gpc4416 (
      {stage3_1[13]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4417 (
      {stage3_1[14]},
      {stage4_1[4]}
   );
   gpc1_1 gpc4418 (
      {stage3_1[15]},
      {stage4_1[5]}
   );
   gpc1_1 gpc4419 (
      {stage3_1[16]},
      {stage4_1[6]}
   );
   gpc1_1 gpc4420 (
      {stage3_1[17]},
      {stage4_1[7]}
   );
   gpc1_1 gpc4421 (
      {stage3_1[18]},
      {stage4_1[8]}
   );
   gpc1_1 gpc4422 (
      {stage3_1[19]},
      {stage4_1[9]}
   );
   gpc1_1 gpc4423 (
      {stage3_1[20]},
      {stage4_1[10]}
   );
   gpc1_1 gpc4424 (
      {stage3_1[21]},
      {stage4_1[11]}
   );
   gpc1_1 gpc4425 (
      {stage3_1[22]},
      {stage4_1[12]}
   );
   gpc1_1 gpc4426 (
      {stage3_1[23]},
      {stage4_1[13]}
   );
   gpc1_1 gpc4427 (
      {stage3_1[24]},
      {stage4_1[14]}
   );
   gpc1_1 gpc4428 (
      {stage3_1[25]},
      {stage4_1[15]}
   );
   gpc1_1 gpc4429 (
      {stage3_2[30]},
      {stage4_2[7]}
   );
   gpc1_1 gpc4430 (
      {stage3_2[31]},
      {stage4_2[8]}
   );
   gpc1_1 gpc4431 (
      {stage3_2[32]},
      {stage4_2[9]}
   );
   gpc1_1 gpc4432 (
      {stage3_2[33]},
      {stage4_2[10]}
   );
   gpc1_1 gpc4433 (
      {stage3_2[34]},
      {stage4_2[11]}
   );
   gpc1_1 gpc4434 (
      {stage3_2[35]},
      {stage4_2[12]}
   );
   gpc1_1 gpc4435 (
      {stage3_3[12]},
      {stage4_3[7]}
   );
   gpc1_1 gpc4436 (
      {stage3_3[13]},
      {stage4_3[8]}
   );
   gpc1_1 gpc4437 (
      {stage3_3[14]},
      {stage4_3[9]}
   );
   gpc1_1 gpc4438 (
      {stage3_3[15]},
      {stage4_3[10]}
   );
   gpc1_1 gpc4439 (
      {stage3_3[16]},
      {stage4_3[11]}
   );
   gpc1_1 gpc4440 (
      {stage3_3[17]},
      {stage4_3[12]}
   );
   gpc1_1 gpc4441 (
      {stage3_3[18]},
      {stage4_3[13]}
   );
   gpc1_1 gpc4442 (
      {stage3_3[19]},
      {stage4_3[14]}
   );
   gpc1_1 gpc4443 (
      {stage3_3[20]},
      {stage4_3[15]}
   );
   gpc1_1 gpc4444 (
      {stage3_3[21]},
      {stage4_3[16]}
   );
   gpc1_1 gpc4445 (
      {stage3_3[22]},
      {stage4_3[17]}
   );
   gpc1_1 gpc4446 (
      {stage3_3[23]},
      {stage4_3[18]}
   );
   gpc1_1 gpc4447 (
      {stage3_3[24]},
      {stage4_3[19]}
   );
   gpc1_1 gpc4448 (
      {stage3_3[25]},
      {stage4_3[20]}
   );
   gpc1_1 gpc4449 (
      {stage3_3[26]},
      {stage4_3[21]}
   );
   gpc1_1 gpc4450 (
      {stage3_3[27]},
      {stage4_3[22]}
   );
   gpc1_1 gpc4451 (
      {stage3_4[30]},
      {stage4_4[7]}
   );
   gpc1_1 gpc4452 (
      {stage3_4[31]},
      {stage4_4[8]}
   );
   gpc1_1 gpc4453 (
      {stage3_4[32]},
      {stage4_4[9]}
   );
   gpc1_1 gpc4454 (
      {stage3_4[33]},
      {stage4_4[10]}
   );
   gpc1_1 gpc4455 (
      {stage3_4[34]},
      {stage4_4[11]}
   );
   gpc1_1 gpc4456 (
      {stage3_4[35]},
      {stage4_4[12]}
   );
   gpc1_1 gpc4457 (
      {stage3_4[36]},
      {stage4_4[13]}
   );
   gpc1_1 gpc4458 (
      {stage3_4[37]},
      {stage4_4[14]}
   );
   gpc1_1 gpc4459 (
      {stage3_4[38]},
      {stage4_4[15]}
   );
   gpc1_1 gpc4460 (
      {stage3_4[39]},
      {stage4_4[16]}
   );
   gpc1_1 gpc4461 (
      {stage3_4[40]},
      {stage4_4[17]}
   );
   gpc1_1 gpc4462 (
      {stage3_4[41]},
      {stage4_4[18]}
   );
   gpc1_1 gpc4463 (
      {stage3_4[42]},
      {stage4_4[19]}
   );
   gpc1_1 gpc4464 (
      {stage3_4[43]},
      {stage4_4[20]}
   );
   gpc1_1 gpc4465 (
      {stage3_4[44]},
      {stage4_4[21]}
   );
   gpc1_1 gpc4466 (
      {stage3_4[45]},
      {stage4_4[22]}
   );
   gpc1_1 gpc4467 (
      {stage3_4[46]},
      {stage4_4[23]}
   );
   gpc1_1 gpc4468 (
      {stage3_5[24]},
      {stage4_5[11]}
   );
   gpc1_1 gpc4469 (
      {stage3_5[25]},
      {stage4_5[12]}
   );
   gpc1_1 gpc4470 (
      {stage3_5[26]},
      {stage4_5[13]}
   );
   gpc1_1 gpc4471 (
      {stage3_5[27]},
      {stage4_5[14]}
   );
   gpc1_1 gpc4472 (
      {stage3_5[28]},
      {stage4_5[15]}
   );
   gpc1_1 gpc4473 (
      {stage3_5[29]},
      {stage4_5[16]}
   );
   gpc1_1 gpc4474 (
      {stage3_5[30]},
      {stage4_5[17]}
   );
   gpc1_1 gpc4475 (
      {stage3_5[31]},
      {stage4_5[18]}
   );
   gpc1_1 gpc4476 (
      {stage3_5[32]},
      {stage4_5[19]}
   );
   gpc1_1 gpc4477 (
      {stage3_5[33]},
      {stage4_5[20]}
   );
   gpc1_1 gpc4478 (
      {stage3_5[34]},
      {stage4_5[21]}
   );
   gpc1_1 gpc4479 (
      {stage3_5[35]},
      {stage4_5[22]}
   );
   gpc1_1 gpc4480 (
      {stage3_5[36]},
      {stage4_5[23]}
   );
   gpc1_1 gpc4481 (
      {stage3_5[37]},
      {stage4_5[24]}
   );
   gpc1_1 gpc4482 (
      {stage3_5[38]},
      {stage4_5[25]}
   );
   gpc1_1 gpc4483 (
      {stage3_5[39]},
      {stage4_5[26]}
   );
   gpc1_1 gpc4484 (
      {stage3_5[40]},
      {stage4_5[27]}
   );
   gpc1_1 gpc4485 (
      {stage3_5[41]},
      {stage4_5[28]}
   );
   gpc1_1 gpc4486 (
      {stage3_5[42]},
      {stage4_5[29]}
   );
   gpc1_1 gpc4487 (
      {stage3_5[43]},
      {stage4_5[30]}
   );
   gpc1_1 gpc4488 (
      {stage3_5[44]},
      {stage4_5[31]}
   );
   gpc1_1 gpc4489 (
      {stage3_5[45]},
      {stage4_5[32]}
   );
   gpc1_1 gpc4490 (
      {stage3_5[46]},
      {stage4_5[33]}
   );
   gpc1_1 gpc4491 (
      {stage3_5[47]},
      {stage4_5[34]}
   );
   gpc1_1 gpc4492 (
      {stage3_5[48]},
      {stage4_5[35]}
   );
   gpc1_1 gpc4493 (
      {stage3_5[49]},
      {stage4_5[36]}
   );
   gpc1_1 gpc4494 (
      {stage3_5[50]},
      {stage4_5[37]}
   );
   gpc1_1 gpc4495 (
      {stage3_5[51]},
      {stage4_5[38]}
   );
   gpc1_1 gpc4496 (
      {stage3_5[52]},
      {stage4_5[39]}
   );
   gpc1_1 gpc4497 (
      {stage3_5[53]},
      {stage4_5[40]}
   );
   gpc1_1 gpc4498 (
      {stage3_5[54]},
      {stage4_5[41]}
   );
   gpc1_1 gpc4499 (
      {stage3_5[55]},
      {stage4_5[42]}
   );
   gpc1_1 gpc4500 (
      {stage3_5[56]},
      {stage4_5[43]}
   );
   gpc1_1 gpc4501 (
      {stage3_5[57]},
      {stage4_5[44]}
   );
   gpc1_1 gpc4502 (
      {stage3_5[58]},
      {stage4_5[45]}
   );
   gpc1_1 gpc4503 (
      {stage3_6[30]},
      {stage4_6[15]}
   );
   gpc1_1 gpc4504 (
      {stage3_6[31]},
      {stage4_6[16]}
   );
   gpc1_1 gpc4505 (
      {stage3_6[32]},
      {stage4_6[17]}
   );
   gpc1_1 gpc4506 (
      {stage3_6[33]},
      {stage4_6[18]}
   );
   gpc1_1 gpc4507 (
      {stage3_6[34]},
      {stage4_6[19]}
   );
   gpc1_1 gpc4508 (
      {stage3_6[35]},
      {stage4_6[20]}
   );
   gpc1_1 gpc4509 (
      {stage3_6[36]},
      {stage4_6[21]}
   );
   gpc1_1 gpc4510 (
      {stage3_6[37]},
      {stage4_6[22]}
   );
   gpc1_1 gpc4511 (
      {stage3_7[45]},
      {stage4_7[13]}
   );
   gpc1_1 gpc4512 (
      {stage3_7[46]},
      {stage4_7[14]}
   );
   gpc1_1 gpc4513 (
      {stage3_8[85]},
      {stage4_8[21]}
   );
   gpc1_1 gpc4514 (
      {stage3_8[86]},
      {stage4_8[22]}
   );
   gpc1_1 gpc4515 (
      {stage3_8[87]},
      {stage4_8[23]}
   );
   gpc1_1 gpc4516 (
      {stage3_8[88]},
      {stage4_8[24]}
   );
   gpc1_1 gpc4517 (
      {stage3_8[89]},
      {stage4_8[25]}
   );
   gpc1_1 gpc4518 (
      {stage3_8[90]},
      {stage4_8[26]}
   );
   gpc1_1 gpc4519 (
      {stage3_8[91]},
      {stage4_8[27]}
   );
   gpc1_1 gpc4520 (
      {stage3_8[92]},
      {stage4_8[28]}
   );
   gpc1_1 gpc4521 (
      {stage3_9[30]},
      {stage4_9[22]}
   );
   gpc1_1 gpc4522 (
      {stage3_9[31]},
      {stage4_9[23]}
   );
   gpc1_1 gpc4523 (
      {stage3_9[32]},
      {stage4_9[24]}
   );
   gpc1_1 gpc4524 (
      {stage3_9[33]},
      {stage4_9[25]}
   );
   gpc1_1 gpc4525 (
      {stage3_9[34]},
      {stage4_9[26]}
   );
   gpc1_1 gpc4526 (
      {stage3_9[35]},
      {stage4_9[27]}
   );
   gpc1_1 gpc4527 (
      {stage3_9[36]},
      {stage4_9[28]}
   );
   gpc1_1 gpc4528 (
      {stage3_9[37]},
      {stage4_9[29]}
   );
   gpc1_1 gpc4529 (
      {stage3_9[38]},
      {stage4_9[30]}
   );
   gpc1_1 gpc4530 (
      {stage3_9[39]},
      {stage4_9[31]}
   );
   gpc1_1 gpc4531 (
      {stage3_9[40]},
      {stage4_9[32]}
   );
   gpc1_1 gpc4532 (
      {stage3_9[41]},
      {stage4_9[33]}
   );
   gpc1_1 gpc4533 (
      {stage3_9[42]},
      {stage4_9[34]}
   );
   gpc1_1 gpc4534 (
      {stage3_9[43]},
      {stage4_9[35]}
   );
   gpc1_1 gpc4535 (
      {stage3_9[44]},
      {stage4_9[36]}
   );
   gpc1_1 gpc4536 (
      {stage3_9[45]},
      {stage4_9[37]}
   );
   gpc1_1 gpc4537 (
      {stage3_9[46]},
      {stage4_9[38]}
   );
   gpc1_1 gpc4538 (
      {stage3_9[47]},
      {stage4_9[39]}
   );
   gpc1_1 gpc4539 (
      {stage3_9[48]},
      {stage4_9[40]}
   );
   gpc1_1 gpc4540 (
      {stage3_9[49]},
      {stage4_9[41]}
   );
   gpc1_1 gpc4541 (
      {stage3_11[31]},
      {stage4_11[19]}
   );
   gpc1_1 gpc4542 (
      {stage3_11[32]},
      {stage4_11[20]}
   );
   gpc1_1 gpc4543 (
      {stage3_11[33]},
      {stage4_11[21]}
   );
   gpc1_1 gpc4544 (
      {stage3_11[34]},
      {stage4_11[22]}
   );
   gpc1_1 gpc4545 (
      {stage3_11[35]},
      {stage4_11[23]}
   );
   gpc1_1 gpc4546 (
      {stage3_11[36]},
      {stage4_11[24]}
   );
   gpc1_1 gpc4547 (
      {stage3_11[37]},
      {stage4_11[25]}
   );
   gpc1_1 gpc4548 (
      {stage3_11[38]},
      {stage4_11[26]}
   );
   gpc1_1 gpc4549 (
      {stage3_11[39]},
      {stage4_11[27]}
   );
   gpc1_1 gpc4550 (
      {stage3_11[40]},
      {stage4_11[28]}
   );
   gpc1_1 gpc4551 (
      {stage3_11[41]},
      {stage4_11[29]}
   );
   gpc1_1 gpc4552 (
      {stage3_11[42]},
      {stage4_11[30]}
   );
   gpc1_1 gpc4553 (
      {stage3_11[43]},
      {stage4_11[31]}
   );
   gpc1_1 gpc4554 (
      {stage3_11[44]},
      {stage4_11[32]}
   );
   gpc1_1 gpc4555 (
      {stage3_11[45]},
      {stage4_11[33]}
   );
   gpc1_1 gpc4556 (
      {stage3_11[46]},
      {stage4_11[34]}
   );
   gpc1_1 gpc4557 (
      {stage3_11[47]},
      {stage4_11[35]}
   );
   gpc1_1 gpc4558 (
      {stage3_11[48]},
      {stage4_11[36]}
   );
   gpc1_1 gpc4559 (
      {stage3_11[49]},
      {stage4_11[37]}
   );
   gpc1_1 gpc4560 (
      {stage3_11[50]},
      {stage4_11[38]}
   );
   gpc1_1 gpc4561 (
      {stage3_11[51]},
      {stage4_11[39]}
   );
   gpc1_1 gpc4562 (
      {stage3_11[52]},
      {stage4_11[40]}
   );
   gpc1_1 gpc4563 (
      {stage3_11[53]},
      {stage4_11[41]}
   );
   gpc1_1 gpc4564 (
      {stage3_11[54]},
      {stage4_11[42]}
   );
   gpc1_1 gpc4565 (
      {stage3_12[38]},
      {stage4_12[15]}
   );
   gpc1_1 gpc4566 (
      {stage3_12[39]},
      {stage4_12[16]}
   );
   gpc1_1 gpc4567 (
      {stage3_12[40]},
      {stage4_12[17]}
   );
   gpc1_1 gpc4568 (
      {stage3_12[41]},
      {stage4_12[18]}
   );
   gpc1_1 gpc4569 (
      {stage3_12[42]},
      {stage4_12[19]}
   );
   gpc1_1 gpc4570 (
      {stage3_12[43]},
      {stage4_12[20]}
   );
   gpc1_1 gpc4571 (
      {stage3_12[44]},
      {stage4_12[21]}
   );
   gpc1_1 gpc4572 (
      {stage3_12[45]},
      {stage4_12[22]}
   );
   gpc1_1 gpc4573 (
      {stage3_12[46]},
      {stage4_12[23]}
   );
   gpc1_1 gpc4574 (
      {stage3_13[29]},
      {stage4_13[11]}
   );
   gpc1_1 gpc4575 (
      {stage3_13[30]},
      {stage4_13[12]}
   );
   gpc1_1 gpc4576 (
      {stage3_13[31]},
      {stage4_13[13]}
   );
   gpc1_1 gpc4577 (
      {stage3_13[32]},
      {stage4_13[14]}
   );
   gpc1_1 gpc4578 (
      {stage3_13[33]},
      {stage4_13[15]}
   );
   gpc1_1 gpc4579 (
      {stage3_13[34]},
      {stage4_13[16]}
   );
   gpc1_1 gpc4580 (
      {stage3_13[35]},
      {stage4_13[17]}
   );
   gpc1_1 gpc4581 (
      {stage3_13[36]},
      {stage4_13[18]}
   );
   gpc1_1 gpc4582 (
      {stage3_14[36]},
      {stage4_14[15]}
   );
   gpc1_1 gpc4583 (
      {stage3_14[37]},
      {stage4_14[16]}
   );
   gpc1_1 gpc4584 (
      {stage3_14[38]},
      {stage4_14[17]}
   );
   gpc1_1 gpc4585 (
      {stage3_14[39]},
      {stage4_14[18]}
   );
   gpc1_1 gpc4586 (
      {stage3_14[40]},
      {stage4_14[19]}
   );
   gpc1_1 gpc4587 (
      {stage3_14[41]},
      {stage4_14[20]}
   );
   gpc1_1 gpc4588 (
      {stage3_14[42]},
      {stage4_14[21]}
   );
   gpc1_1 gpc4589 (
      {stage3_14[43]},
      {stage4_14[22]}
   );
   gpc1_1 gpc4590 (
      {stage3_14[44]},
      {stage4_14[23]}
   );
   gpc1_1 gpc4591 (
      {stage3_14[45]},
      {stage4_14[24]}
   );
   gpc1_1 gpc4592 (
      {stage3_14[46]},
      {stage4_14[25]}
   );
   gpc1_1 gpc4593 (
      {stage3_14[47]},
      {stage4_14[26]}
   );
   gpc1_1 gpc4594 (
      {stage3_14[48]},
      {stage4_14[27]}
   );
   gpc1_1 gpc4595 (
      {stage3_14[49]},
      {stage4_14[28]}
   );
   gpc1_1 gpc4596 (
      {stage3_14[50]},
      {stage4_14[29]}
   );
   gpc1_1 gpc4597 (
      {stage3_14[51]},
      {stage4_14[30]}
   );
   gpc1_1 gpc4598 (
      {stage3_14[52]},
      {stage4_14[31]}
   );
   gpc1_1 gpc4599 (
      {stage3_14[53]},
      {stage4_14[32]}
   );
   gpc1_1 gpc4600 (
      {stage3_14[54]},
      {stage4_14[33]}
   );
   gpc1_1 gpc4601 (
      {stage3_14[55]},
      {stage4_14[34]}
   );
   gpc1_1 gpc4602 (
      {stage3_15[55]},
      {stage4_15[23]}
   );
   gpc1_1 gpc4603 (
      {stage3_15[56]},
      {stage4_15[24]}
   );
   gpc1_1 gpc4604 (
      {stage3_15[57]},
      {stage4_15[25]}
   );
   gpc1_1 gpc4605 (
      {stage3_15[58]},
      {stage4_15[26]}
   );
   gpc1_1 gpc4606 (
      {stage3_15[59]},
      {stage4_15[27]}
   );
   gpc1_1 gpc4607 (
      {stage3_15[60]},
      {stage4_15[28]}
   );
   gpc1_1 gpc4608 (
      {stage3_15[61]},
      {stage4_15[29]}
   );
   gpc1_1 gpc4609 (
      {stage3_15[62]},
      {stage4_15[30]}
   );
   gpc1_1 gpc4610 (
      {stage3_15[63]},
      {stage4_15[31]}
   );
   gpc1_1 gpc4611 (
      {stage3_15[64]},
      {stage4_15[32]}
   );
   gpc1_1 gpc4612 (
      {stage3_15[65]},
      {stage4_15[33]}
   );
   gpc1_1 gpc4613 (
      {stage3_15[66]},
      {stage4_15[34]}
   );
   gpc1_1 gpc4614 (
      {stage3_15[67]},
      {stage4_15[35]}
   );
   gpc1_1 gpc4615 (
      {stage3_15[68]},
      {stage4_15[36]}
   );
   gpc1_1 gpc4616 (
      {stage3_15[69]},
      {stage4_15[37]}
   );
   gpc1_1 gpc4617 (
      {stage3_15[70]},
      {stage4_15[38]}
   );
   gpc1_1 gpc4618 (
      {stage3_17[55]},
      {stage4_17[21]}
   );
   gpc1_1 gpc4619 (
      {stage3_17[56]},
      {stage4_17[22]}
   );
   gpc1_1 gpc4620 (
      {stage3_17[57]},
      {stage4_17[23]}
   );
   gpc1_1 gpc4621 (
      {stage3_17[58]},
      {stage4_17[24]}
   );
   gpc1_1 gpc4622 (
      {stage3_17[59]},
      {stage4_17[25]}
   );
   gpc1_1 gpc4623 (
      {stage3_17[60]},
      {stage4_17[26]}
   );
   gpc1_1 gpc4624 (
      {stage3_17[61]},
      {stage4_17[27]}
   );
   gpc1_1 gpc4625 (
      {stage3_17[62]},
      {stage4_17[28]}
   );
   gpc1_1 gpc4626 (
      {stage3_17[63]},
      {stage4_17[29]}
   );
   gpc1_1 gpc4627 (
      {stage3_17[64]},
      {stage4_17[30]}
   );
   gpc1_1 gpc4628 (
      {stage3_17[65]},
      {stage4_17[31]}
   );
   gpc1_1 gpc4629 (
      {stage3_17[66]},
      {stage4_17[32]}
   );
   gpc1_1 gpc4630 (
      {stage3_17[67]},
      {stage4_17[33]}
   );
   gpc1_1 gpc4631 (
      {stage3_17[68]},
      {stage4_17[34]}
   );
   gpc1_1 gpc4632 (
      {stage3_17[69]},
      {stage4_17[35]}
   );
   gpc1_1 gpc4633 (
      {stage3_17[70]},
      {stage4_17[36]}
   );
   gpc1_1 gpc4634 (
      {stage3_17[71]},
      {stage4_17[37]}
   );
   gpc1_1 gpc4635 (
      {stage3_17[72]},
      {stage4_17[38]}
   );
   gpc1_1 gpc4636 (
      {stage3_17[73]},
      {stage4_17[39]}
   );
   gpc1_1 gpc4637 (
      {stage3_17[74]},
      {stage4_17[40]}
   );
   gpc1_1 gpc4638 (
      {stage3_17[75]},
      {stage4_17[41]}
   );
   gpc1_1 gpc4639 (
      {stage3_17[76]},
      {stage4_17[42]}
   );
   gpc1_1 gpc4640 (
      {stage3_18[25]},
      {stage4_18[19]}
   );
   gpc1_1 gpc4641 (
      {stage3_18[26]},
      {stage4_18[20]}
   );
   gpc1_1 gpc4642 (
      {stage3_18[27]},
      {stage4_18[21]}
   );
   gpc1_1 gpc4643 (
      {stage3_18[28]},
      {stage4_18[22]}
   );
   gpc1_1 gpc4644 (
      {stage3_18[29]},
      {stage4_18[23]}
   );
   gpc1_1 gpc4645 (
      {stage3_18[30]},
      {stage4_18[24]}
   );
   gpc1_1 gpc4646 (
      {stage3_18[31]},
      {stage4_18[25]}
   );
   gpc1_1 gpc4647 (
      {stage3_18[32]},
      {stage4_18[26]}
   );
   gpc1_1 gpc4648 (
      {stage3_18[33]},
      {stage4_18[27]}
   );
   gpc1_1 gpc4649 (
      {stage3_18[34]},
      {stage4_18[28]}
   );
   gpc1_1 gpc4650 (
      {stage3_19[62]},
      {stage4_19[24]}
   );
   gpc1_1 gpc4651 (
      {stage3_19[63]},
      {stage4_19[25]}
   );
   gpc1_1 gpc4652 (
      {stage3_19[64]},
      {stage4_19[26]}
   );
   gpc1_1 gpc4653 (
      {stage3_19[65]},
      {stage4_19[27]}
   );
   gpc1_1 gpc4654 (
      {stage3_19[66]},
      {stage4_19[28]}
   );
   gpc1_1 gpc4655 (
      {stage3_19[67]},
      {stage4_19[29]}
   );
   gpc1_1 gpc4656 (
      {stage3_19[68]},
      {stage4_19[30]}
   );
   gpc1_1 gpc4657 (
      {stage3_19[69]},
      {stage4_19[31]}
   );
   gpc1_1 gpc4658 (
      {stage3_21[60]},
      {stage4_21[16]}
   );
   gpc1_1 gpc4659 (
      {stage3_21[61]},
      {stage4_21[17]}
   );
   gpc1_1 gpc4660 (
      {stage3_21[62]},
      {stage4_21[18]}
   );
   gpc1_1 gpc4661 (
      {stage3_22[37]},
      {stage4_22[17]}
   );
   gpc1_1 gpc4662 (
      {stage3_22[38]},
      {stage4_22[18]}
   );
   gpc1_1 gpc4663 (
      {stage3_22[39]},
      {stage4_22[19]}
   );
   gpc1_1 gpc4664 (
      {stage3_22[40]},
      {stage4_22[20]}
   );
   gpc1_1 gpc4665 (
      {stage3_22[41]},
      {stage4_22[21]}
   );
   gpc1_1 gpc4666 (
      {stage3_22[42]},
      {stage4_22[22]}
   );
   gpc1_1 gpc4667 (
      {stage3_22[43]},
      {stage4_22[23]}
   );
   gpc1_1 gpc4668 (
      {stage3_22[44]},
      {stage4_22[24]}
   );
   gpc1_1 gpc4669 (
      {stage3_22[45]},
      {stage4_22[25]}
   );
   gpc1_1 gpc4670 (
      {stage3_22[46]},
      {stage4_22[26]}
   );
   gpc1_1 gpc4671 (
      {stage3_22[47]},
      {stage4_22[27]}
   );
   gpc1_1 gpc4672 (
      {stage3_22[48]},
      {stage4_22[28]}
   );
   gpc1_1 gpc4673 (
      {stage3_22[49]},
      {stage4_22[29]}
   );
   gpc1_1 gpc4674 (
      {stage3_22[50]},
      {stage4_22[30]}
   );
   gpc1_1 gpc4675 (
      {stage3_23[29]},
      {stage4_23[21]}
   );
   gpc1_1 gpc4676 (
      {stage3_23[30]},
      {stage4_23[22]}
   );
   gpc1_1 gpc4677 (
      {stage3_23[31]},
      {stage4_23[23]}
   );
   gpc1_1 gpc4678 (
      {stage3_23[32]},
      {stage4_23[24]}
   );
   gpc1_1 gpc4679 (
      {stage3_23[33]},
      {stage4_23[25]}
   );
   gpc1_1 gpc4680 (
      {stage3_23[34]},
      {stage4_23[26]}
   );
   gpc1_1 gpc4681 (
      {stage3_23[35]},
      {stage4_23[27]}
   );
   gpc1_1 gpc4682 (
      {stage3_23[36]},
      {stage4_23[28]}
   );
   gpc1_1 gpc4683 (
      {stage3_23[37]},
      {stage4_23[29]}
   );
   gpc1_1 gpc4684 (
      {stage3_23[38]},
      {stage4_23[30]}
   );
   gpc1_1 gpc4685 (
      {stage3_23[39]},
      {stage4_23[31]}
   );
   gpc1_1 gpc4686 (
      {stage3_23[40]},
      {stage4_23[32]}
   );
   gpc1_1 gpc4687 (
      {stage3_23[41]},
      {stage4_23[33]}
   );
   gpc1_1 gpc4688 (
      {stage3_23[42]},
      {stage4_23[34]}
   );
   gpc1_1 gpc4689 (
      {stage3_23[43]},
      {stage4_23[35]}
   );
   gpc1_1 gpc4690 (
      {stage3_23[44]},
      {stage4_23[36]}
   );
   gpc1_1 gpc4691 (
      {stage3_23[45]},
      {stage4_23[37]}
   );
   gpc1_1 gpc4692 (
      {stage3_24[47]},
      {stage4_24[16]}
   );
   gpc1_1 gpc4693 (
      {stage3_24[48]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4694 (
      {stage3_24[49]},
      {stage4_24[18]}
   );
   gpc1_1 gpc4695 (
      {stage3_24[50]},
      {stage4_24[19]}
   );
   gpc1_1 gpc4696 (
      {stage3_24[51]},
      {stage4_24[20]}
   );
   gpc1_1 gpc4697 (
      {stage3_24[52]},
      {stage4_24[21]}
   );
   gpc1_1 gpc4698 (
      {stage3_24[53]},
      {stage4_24[22]}
   );
   gpc1_1 gpc4699 (
      {stage3_24[54]},
      {stage4_24[23]}
   );
   gpc1_1 gpc4700 (
      {stage3_24[55]},
      {stage4_24[24]}
   );
   gpc1_1 gpc4701 (
      {stage3_24[56]},
      {stage4_24[25]}
   );
   gpc1_1 gpc4702 (
      {stage3_24[57]},
      {stage4_24[26]}
   );
   gpc1_1 gpc4703 (
      {stage3_24[58]},
      {stage4_24[27]}
   );
   gpc1_1 gpc4704 (
      {stage3_24[59]},
      {stage4_24[28]}
   );
   gpc1_1 gpc4705 (
      {stage3_24[60]},
      {stage4_24[29]}
   );
   gpc1_1 gpc4706 (
      {stage3_25[47]},
      {stage4_25[17]}
   );
   gpc1_1 gpc4707 (
      {stage3_25[48]},
      {stage4_25[18]}
   );
   gpc1_1 gpc4708 (
      {stage3_26[46]},
      {stage4_26[18]}
   );
   gpc1_1 gpc4709 (
      {stage3_26[47]},
      {stage4_26[19]}
   );
   gpc1_1 gpc4710 (
      {stage3_26[48]},
      {stage4_26[20]}
   );
   gpc1_1 gpc4711 (
      {stage3_26[49]},
      {stage4_26[21]}
   );
   gpc1_1 gpc4712 (
      {stage3_26[50]},
      {stage4_26[22]}
   );
   gpc1_1 gpc4713 (
      {stage3_27[48]},
      {stage4_27[20]}
   );
   gpc1_1 gpc4714 (
      {stage3_27[49]},
      {stage4_27[21]}
   );
   gpc1_1 gpc4715 (
      {stage3_27[50]},
      {stage4_27[22]}
   );
   gpc1_1 gpc4716 (
      {stage3_27[51]},
      {stage4_27[23]}
   );
   gpc1_1 gpc4717 (
      {stage3_27[52]},
      {stage4_27[24]}
   );
   gpc1_1 gpc4718 (
      {stage3_27[53]},
      {stage4_27[25]}
   );
   gpc1_1 gpc4719 (
      {stage3_27[54]},
      {stage4_27[26]}
   );
   gpc1_1 gpc4720 (
      {stage3_30[68]},
      {stage4_30[24]}
   );
   gpc1_1 gpc4721 (
      {stage3_30[69]},
      {stage4_30[25]}
   );
   gpc1_1 gpc4722 (
      {stage3_30[70]},
      {stage4_30[26]}
   );
   gpc1_1 gpc4723 (
      {stage3_31[51]},
      {stage4_31[24]}
   );
   gpc1_1 gpc4724 (
      {stage3_31[52]},
      {stage4_31[25]}
   );
   gpc1_1 gpc4725 (
      {stage3_31[53]},
      {stage4_31[26]}
   );
   gpc1_1 gpc4726 (
      {stage3_31[54]},
      {stage4_31[27]}
   );
   gpc1_1 gpc4727 (
      {stage3_31[55]},
      {stage4_31[28]}
   );
   gpc1_1 gpc4728 (
      {stage3_31[56]},
      {stage4_31[29]}
   );
   gpc1_1 gpc4729 (
      {stage3_31[57]},
      {stage4_31[30]}
   );
   gpc1_1 gpc4730 (
      {stage3_32[39]},
      {stage4_32[24]}
   );
   gpc1_1 gpc4731 (
      {stage3_32[40]},
      {stage4_32[25]}
   );
   gpc1_1 gpc4732 (
      {stage3_32[41]},
      {stage4_32[26]}
   );
   gpc1_1 gpc4733 (
      {stage3_32[42]},
      {stage4_32[27]}
   );
   gpc1_1 gpc4734 (
      {stage3_32[43]},
      {stage4_32[28]}
   );
   gpc1_1 gpc4735 (
      {stage3_32[44]},
      {stage4_32[29]}
   );
   gpc1_1 gpc4736 (
      {stage3_32[45]},
      {stage4_32[30]}
   );
   gpc1_1 gpc4737 (
      {stage3_32[46]},
      {stage4_32[31]}
   );
   gpc1_1 gpc4738 (
      {stage3_32[47]},
      {stage4_32[32]}
   );
   gpc1_1 gpc4739 (
      {stage3_32[48]},
      {stage4_32[33]}
   );
   gpc1_1 gpc4740 (
      {stage3_32[49]},
      {stage4_32[34]}
   );
   gpc1_1 gpc4741 (
      {stage3_32[50]},
      {stage4_32[35]}
   );
   gpc1_1 gpc4742 (
      {stage3_32[51]},
      {stage4_32[36]}
   );
   gpc1_1 gpc4743 (
      {stage3_32[52]},
      {stage4_32[37]}
   );
   gpc1_1 gpc4744 (
      {stage3_32[53]},
      {stage4_32[38]}
   );
   gpc1_1 gpc4745 (
      {stage3_32[54]},
      {stage4_32[39]}
   );
   gpc1_1 gpc4746 (
      {stage3_32[55]},
      {stage4_32[40]}
   );
   gpc1_1 gpc4747 (
      {stage3_32[56]},
      {stage4_32[41]}
   );
   gpc1_1 gpc4748 (
      {stage3_32[57]},
      {stage4_32[42]}
   );
   gpc1_1 gpc4749 (
      {stage3_33[24]},
      {stage4_33[16]}
   );
   gpc1_1 gpc4750 (
      {stage3_33[25]},
      {stage4_33[17]}
   );
   gpc1_1 gpc4751 (
      {stage3_33[26]},
      {stage4_33[18]}
   );
   gpc1_1 gpc4752 (
      {stage3_34[24]},
      {stage4_34[10]}
   );
   gpc1_1 gpc4753 (
      {stage3_34[25]},
      {stage4_34[11]}
   );
   gpc1_1 gpc4754 (
      {stage3_34[26]},
      {stage4_34[12]}
   );
   gpc1_1 gpc4755 (
      {stage3_35[6]},
      {stage4_35[8]}
   );
   gpc1_1 gpc4756 (
      {stage3_35[7]},
      {stage4_35[9]}
   );
   gpc1_1 gpc4757 (
      {stage3_35[8]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4758 (
      {stage3_35[9]},
      {stage4_35[11]}
   );
   gpc1_1 gpc4759 (
      {stage3_35[10]},
      {stage4_35[12]}
   );
   gpc1_1 gpc4760 (
      {stage3_35[11]},
      {stage4_35[13]}
   );
   gpc1_1 gpc4761 (
      {stage3_35[12]},
      {stage4_35[14]}
   );
   gpc1_1 gpc4762 (
      {stage3_36[0]},
      {stage4_36[5]}
   );
   gpc1_1 gpc4763 (
      {stage3_36[1]},
      {stage4_36[6]}
   );
   gpc1_1 gpc4764 (
      {stage3_36[2]},
      {stage4_36[7]}
   );
   gpc1_1 gpc4765 (
      {stage3_36[3]},
      {stage4_36[8]}
   );
   gpc1_1 gpc4766 (
      {stage3_36[4]},
      {stage4_36[9]}
   );
   gpc1_1 gpc4767 (
      {stage3_36[5]},
      {stage4_36[10]}
   );
   gpc1_1 gpc4768 (
      {stage3_37[0]},
      {stage4_37[1]}
   );
   gpc1_1 gpc4769 (
      {stage3_37[1]},
      {stage4_37[2]}
   );
   gpc606_5 gpc4770 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc615_5 gpc4771 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[6]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[1],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc615_5 gpc4772 (
      {stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[6]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[1],stage5_5[2],stage5_4[2],stage5_3[2]}
   );
   gpc615_5 gpc4773 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16]},
      {stage4_4[7]},
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage5_7[1],stage5_6[2],stage5_5[3],stage5_4[3],stage5_3[3]}
   );
   gpc615_5 gpc4774 (
      {stage4_3[17], stage4_3[18], stage4_3[19], stage4_3[20], stage4_3[21]},
      {stage4_4[8]},
      {stage4_5[12], stage4_5[13], stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17]},
      {stage5_7[2],stage5_6[3],stage5_5[4],stage5_4[4],stage5_3[4]}
   );
   gpc606_5 gpc4775 (
      {stage4_4[9], stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[3],stage5_6[4],stage5_5[5],stage5_4[5]}
   );
   gpc606_5 gpc4776 (
      {stage4_4[15], stage4_4[16], stage4_4[17], stage4_4[18], stage4_4[19], stage4_4[20]},
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11]},
      {stage5_8[1],stage5_7[4],stage5_6[5],stage5_5[6],stage5_4[6]}
   );
   gpc7_3 gpc4777 (
      {stage4_5[18], stage4_5[19], stage4_5[20], stage4_5[21], stage4_5[22], stage4_5[23], stage4_5[24]},
      {stage5_7[5],stage5_6[6],stage5_5[7]}
   );
   gpc7_3 gpc4778 (
      {stage4_5[25], stage4_5[26], stage4_5[27], stage4_5[28], stage4_5[29], stage4_5[30], stage4_5[31]},
      {stage5_7[6],stage5_6[7],stage5_5[8]}
   );
   gpc7_3 gpc4779 (
      {stage4_5[32], stage4_5[33], stage4_5[34], stage4_5[35], stage4_5[36], stage4_5[37], stage4_5[38]},
      {stage5_7[7],stage5_6[8],stage5_5[9]}
   );
   gpc7_3 gpc4780 (
      {stage4_5[39], stage4_5[40], stage4_5[41], stage4_5[42], stage4_5[43], stage4_5[44], stage4_5[45]},
      {stage5_7[8],stage5_6[9],stage5_5[10]}
   );
   gpc615_5 gpc4781 (
      {stage4_6[12], stage4_6[13], stage4_6[14], stage4_6[15], stage4_6[16]},
      {stage4_7[0]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[2],stage5_7[9],stage5_6[10]}
   );
   gpc615_5 gpc4782 (
      {stage4_6[17], stage4_6[18], stage4_6[19], stage4_6[20], stage4_6[21]},
      {stage4_7[1]},
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage5_10[1],stage5_9[1],stage5_8[3],stage5_7[10],stage5_6[11]}
   );
   gpc1163_5 gpc4783 (
      {stage4_7[2], stage4_7[3], stage4_7[4]},
      {stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17]},
      {stage4_9[0]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[4],stage5_7[11]}
   );
   gpc623_5 gpc4784 (
      {stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[18], stage4_8[19]},
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[5],stage5_7[12]}
   );
   gpc606_5 gpc4785 (
      {stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24], stage4_8[25]},
      {stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6]},
      {stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[4],stage5_8[6]}
   );
   gpc606_5 gpc4786 (
      {stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[5]}
   );
   gpc606_5 gpc4787 (
      {stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16], stage4_9[17], stage4_9[18]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[6]}
   );
   gpc606_5 gpc4788 (
      {stage4_9[19], stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23], stage4_9[24]},
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage5_13[2],stage5_12[3],stage5_11[5],stage5_10[7],stage5_9[7]}
   );
   gpc606_5 gpc4789 (
      {stage4_9[25], stage4_9[26], stage4_9[27], stage4_9[28], stage4_9[29], stage4_9[30]},
      {stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21], stage4_11[22], stage4_11[23]},
      {stage5_13[3],stage5_12[4],stage5_11[6],stage5_10[8],stage5_9[8]}
   );
   gpc606_5 gpc4790 (
      {stage4_9[31], stage4_9[32], stage4_9[33], stage4_9[34], stage4_9[35], stage4_9[36]},
      {stage4_11[24], stage4_11[25], stage4_11[26], stage4_11[27], stage4_11[28], stage4_11[29]},
      {stage5_13[4],stage5_12[5],stage5_11[7],stage5_10[9],stage5_9[9]}
   );
   gpc615_5 gpc4791 (
      {stage4_9[37], stage4_9[38], stage4_9[39], stage4_9[40], stage4_9[41]},
      {stage4_10[7]},
      {stage4_11[30], stage4_11[31], stage4_11[32], stage4_11[33], stage4_11[34], stage4_11[35]},
      {stage5_13[5],stage5_12[6],stage5_11[8],stage5_10[10],stage5_9[10]}
   );
   gpc615_5 gpc4792 (
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12]},
      {stage4_11[36]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[6],stage5_12[7],stage5_11[9],stage5_10[11]}
   );
   gpc615_5 gpc4793 (
      {stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17]},
      {stage4_11[37]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[7],stage5_12[8],stage5_11[10],stage5_10[12]}
   );
   gpc606_5 gpc4794 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[8],stage5_12[9]}
   );
   gpc606_5 gpc4795 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[1],stage5_14[3],stage5_13[9],stage5_12[10]}
   );
   gpc1163_5 gpc4796 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16], stage4_14[17]},
      {stage4_15[0]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[2],stage5_15[2],stage5_14[4],stage5_13[10]}
   );
   gpc1163_5 gpc4797 (
      {stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_14[18], stage4_14[19], stage4_14[20], stage4_14[21], stage4_14[22], stage4_14[23]},
      {stage4_15[1]},
      {stage4_16[1]},
      {stage5_17[1],stage5_16[3],stage5_15[3],stage5_14[5],stage5_13[11]}
   );
   gpc1163_5 gpc4798 (
      {stage4_13[6], stage4_13[7], stage4_13[8]},
      {stage4_14[24], stage4_14[25], stage4_14[26], stage4_14[27], stage4_14[28], stage4_14[29]},
      {stage4_15[2]},
      {stage4_16[2]},
      {stage5_17[2],stage5_16[4],stage5_15[4],stage5_14[6],stage5_13[12]}
   );
   gpc606_5 gpc4799 (
      {stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13], stage4_13[14]},
      {stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6], stage4_15[7], stage4_15[8]},
      {stage5_17[3],stage5_16[5],stage5_15[5],stage5_14[7],stage5_13[13]}
   );
   gpc606_5 gpc4800 (
      {stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], 1'b0, 1'b0},
      {stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12], stage4_15[13], stage4_15[14]},
      {stage5_17[4],stage5_16[6],stage5_15[6],stage5_14[8],stage5_13[14]}
   );
   gpc135_4 gpc4801 (
      {stage4_14[30], stage4_14[31], stage4_14[32], stage4_14[33], stage4_14[34]},
      {stage4_15[15], stage4_15[16], stage4_15[17]},
      {stage4_16[3]},
      {stage5_17[5],stage5_16[7],stage5_15[7],stage5_14[9]}
   );
   gpc615_5 gpc4802 (
      {stage4_15[18], stage4_15[19], stage4_15[20], stage4_15[21], stage4_15[22]},
      {stage4_16[4]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[6],stage5_16[8],stage5_15[8]}
   );
   gpc615_5 gpc4803 (
      {stage4_15[23], stage4_15[24], stage4_15[25], stage4_15[26], stage4_15[27]},
      {stage4_16[5]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[1],stage5_17[7],stage5_16[9],stage5_15[9]}
   );
   gpc615_5 gpc4804 (
      {stage4_15[28], stage4_15[29], stage4_15[30], stage4_15[31], stage4_15[32]},
      {stage4_16[6]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[2],stage5_17[8],stage5_16[10],stage5_15[10]}
   );
   gpc615_5 gpc4805 (
      {stage4_15[33], stage4_15[34], stage4_15[35], stage4_15[36], stage4_15[37]},
      {stage4_16[7]},
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], stage4_17[22], stage4_17[23]},
      {stage5_19[3],stage5_18[3],stage5_17[9],stage5_16[11],stage5_15[11]}
   );
   gpc606_5 gpc4806 (
      {stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12], stage4_16[13]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[4],stage5_18[4],stage5_17[10],stage5_16[12]}
   );
   gpc615_5 gpc4807 (
      {stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_17[24]},
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage5_20[1],stage5_19[5],stage5_18[5],stage5_17[11],stage5_16[13]}
   );
   gpc606_5 gpc4808 (
      {stage4_17[25], stage4_17[26], stage4_17[27], stage4_17[28], stage4_17[29], stage4_17[30]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[2],stage5_19[6],stage5_18[6],stage5_17[12]}
   );
   gpc606_5 gpc4809 (
      {stage4_17[31], stage4_17[32], stage4_17[33], stage4_17[34], stage4_17[35], stage4_17[36]},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[3],stage5_19[7],stage5_18[7],stage5_17[13]}
   );
   gpc606_5 gpc4810 (
      {stage4_17[37], stage4_17[38], stage4_17[39], stage4_17[40], stage4_17[41], stage4_17[42]},
      {stage4_19[12], stage4_19[13], stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17]},
      {stage5_21[2],stage5_20[4],stage5_19[8],stage5_18[8],stage5_17[14]}
   );
   gpc606_5 gpc4811 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[3],stage5_20[5],stage5_19[9],stage5_18[9]}
   );
   gpc615_5 gpc4812 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22]},
      {stage4_19[18]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[4],stage5_20[6],stage5_19[10],stage5_18[10]}
   );
   gpc615_5 gpc4813 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4]},
      {stage4_22[0]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[2],stage5_21[5]}
   );
   gpc615_5 gpc4814 (
      {stage4_21[5], stage4_21[6], stage4_21[7], stage4_21[8], stage4_21[9]},
      {stage4_22[1]},
      {stage4_23[6], stage4_23[7], stage4_23[8], stage4_23[9], stage4_23[10], stage4_23[11]},
      {stage5_25[1],stage5_24[1],stage5_23[1],stage5_22[3],stage5_21[6]}
   );
   gpc615_5 gpc4815 (
      {stage4_21[10], stage4_21[11], stage4_21[12], stage4_21[13], stage4_21[14]},
      {stage4_22[2]},
      {stage4_23[12], stage4_23[13], stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17]},
      {stage5_25[2],stage5_24[2],stage5_23[2],stage5_22[4],stage5_21[7]}
   );
   gpc615_5 gpc4816 (
      {stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18], 1'b0},
      {stage4_22[3]},
      {stage4_23[18], stage4_23[19], stage4_23[20], stage4_23[21], stage4_23[22], stage4_23[23]},
      {stage5_25[3],stage5_24[3],stage5_23[3],stage5_22[5],stage5_21[8]}
   );
   gpc615_5 gpc4817 (
      {stage4_22[4], stage4_22[5], stage4_22[6], stage4_22[7], stage4_22[8]},
      {stage4_23[24]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[4],stage5_24[4],stage5_23[4],stage5_22[6]}
   );
   gpc615_5 gpc4818 (
      {stage4_22[9], stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13]},
      {stage4_23[25]},
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage5_26[1],stage5_25[5],stage5_24[5],stage5_23[5],stage5_22[7]}
   );
   gpc615_5 gpc4819 (
      {stage4_22[14], stage4_22[15], stage4_22[16], stage4_22[17], stage4_22[18]},
      {stage4_23[26]},
      {stage4_24[12], stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17]},
      {stage5_26[2],stage5_25[6],stage5_24[6],stage5_23[6],stage5_22[8]}
   );
   gpc615_5 gpc4820 (
      {stage4_22[19], stage4_22[20], stage4_22[21], stage4_22[22], stage4_22[23]},
      {stage4_23[27]},
      {stage4_24[18], stage4_24[19], stage4_24[20], stage4_24[21], stage4_24[22], stage4_24[23]},
      {stage5_26[3],stage5_25[7],stage5_24[7],stage5_23[7],stage5_22[9]}
   );
   gpc615_5 gpc4821 (
      {stage4_23[28], stage4_23[29], stage4_23[30], stage4_23[31], stage4_23[32]},
      {stage4_24[24]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[4],stage5_25[8],stage5_24[8],stage5_23[8]}
   );
   gpc615_5 gpc4822 (
      {stage4_23[33], stage4_23[34], stage4_23[35], stage4_23[36], stage4_23[37]},
      {stage4_24[25]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[5],stage5_25[9],stage5_24[9],stage5_23[9]}
   );
   gpc606_5 gpc4823 (
      {stage4_25[12], stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], stage4_25[17]},
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage5_29[0],stage5_28[0],stage5_27[2],stage5_26[6],stage5_25[10]}
   );
   gpc615_5 gpc4824 (
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4]},
      {stage4_27[6]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[1],stage5_28[1],stage5_27[3],stage5_26[7]}
   );
   gpc615_5 gpc4825 (
      {stage4_26[5], stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9]},
      {stage4_27[7]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[2],stage5_28[2],stage5_27[4],stage5_26[8]}
   );
   gpc615_5 gpc4826 (
      {stage4_26[10], stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14]},
      {stage4_27[8]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[3],stage5_28[3],stage5_27[5],stage5_26[9]}
   );
   gpc615_5 gpc4827 (
      {stage4_26[15], stage4_26[16], stage4_26[17], stage4_26[18], stage4_26[19]},
      {stage4_27[9]},
      {stage4_28[18], stage4_28[19], stage4_28[20], stage4_28[21], stage4_28[22], stage4_28[23]},
      {stage5_30[3],stage5_29[4],stage5_28[4],stage5_27[6],stage5_26[10]}
   );
   gpc207_4 gpc4828 (
      {stage4_27[10], stage4_27[11], stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[4],stage5_29[5],stage5_28[5],stage5_27[7]}
   );
   gpc615_5 gpc4829 (
      {stage4_27[17], stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21]},
      {stage4_28[24]},
      {stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5], stage4_29[6], stage4_29[7]},
      {stage5_31[0],stage5_30[5],stage5_29[6],stage5_28[6],stage5_27[8]}
   );
   gpc615_5 gpc4830 (
      {stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[1],stage5_30[6],stage5_29[7]}
   );
   gpc615_5 gpc4831 (
      {stage4_29[13], stage4_29[14], stage4_29[15], stage4_29[16], stage4_29[17]},
      {stage4_30[1]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage5_33[1],stage5_32[1],stage5_31[2],stage5_30[7],stage5_29[8]}
   );
   gpc615_5 gpc4832 (
      {stage4_29[18], stage4_29[19], stage4_29[20], stage4_29[21], stage4_29[22]},
      {stage4_30[2]},
      {stage4_31[12], stage4_31[13], stage4_31[14], stage4_31[15], stage4_31[16], stage4_31[17]},
      {stage5_33[2],stage5_32[2],stage5_31[3],stage5_30[8],stage5_29[9]}
   );
   gpc615_5 gpc4833 (
      {stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6], stage4_30[7]},
      {stage4_31[18]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[3],stage5_32[3],stage5_31[4],stage5_30[9]}
   );
   gpc615_5 gpc4834 (
      {stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11], stage4_30[12]},
      {stage4_31[19]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[4],stage5_32[4],stage5_31[5],stage5_30[10]}
   );
   gpc615_5 gpc4835 (
      {stage4_30[13], stage4_30[14], stage4_30[15], stage4_30[16], stage4_30[17]},
      {stage4_31[20]},
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage5_34[2],stage5_33[5],stage5_32[5],stage5_31[6],stage5_30[11]}
   );
   gpc615_5 gpc4836 (
      {stage4_30[18], stage4_30[19], stage4_30[20], stage4_30[21], stage4_30[22]},
      {stage4_31[21]},
      {stage4_32[18], stage4_32[19], stage4_32[20], stage4_32[21], stage4_32[22], stage4_32[23]},
      {stage5_34[3],stage5_33[6],stage5_32[6],stage5_31[7],stage5_30[12]}
   );
   gpc615_5 gpc4837 (
      {stage4_31[22], stage4_31[23], stage4_31[24], stage4_31[25], stage4_31[26]},
      {stage4_32[24]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[4],stage5_33[7],stage5_32[7],stage5_31[8]}
   );
   gpc606_5 gpc4838 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[5],stage5_33[8]}
   );
   gpc606_5 gpc4839 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], stage4_33[17]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[1],stage5_35[2],stage5_34[6],stage5_33[9]}
   );
   gpc606_5 gpc4840 (
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage5_38[0],stage5_37[2],stage5_36[2],stage5_35[3],stage5_34[7]}
   );
   gpc606_5 gpc4841 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], 1'b0},
      {stage5_38[1],stage5_37[3],stage5_36[3],stage5_35[4],stage5_34[8]}
   );
   gpc1_1 gpc4842 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc4843 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4844 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc4845 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc4846 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc4847 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc4848 (
      {stage4_0[6]},
      {stage5_0[6]}
   );
   gpc1_1 gpc4849 (
      {stage4_0[7]},
      {stage5_0[7]}
   );
   gpc1_1 gpc4850 (
      {stage4_0[8]},
      {stage5_0[8]}
   );
   gpc1_1 gpc4851 (
      {stage4_0[9]},
      {stage5_0[9]}
   );
   gpc1_1 gpc4852 (
      {stage4_0[10]},
      {stage5_0[10]}
   );
   gpc1_1 gpc4853 (
      {stage4_1[6]},
      {stage5_1[1]}
   );
   gpc1_1 gpc4854 (
      {stage4_1[7]},
      {stage5_1[2]}
   );
   gpc1_1 gpc4855 (
      {stage4_1[8]},
      {stage5_1[3]}
   );
   gpc1_1 gpc4856 (
      {stage4_1[9]},
      {stage5_1[4]}
   );
   gpc1_1 gpc4857 (
      {stage4_1[10]},
      {stage5_1[5]}
   );
   gpc1_1 gpc4858 (
      {stage4_1[11]},
      {stage5_1[6]}
   );
   gpc1_1 gpc4859 (
      {stage4_1[12]},
      {stage5_1[7]}
   );
   gpc1_1 gpc4860 (
      {stage4_1[13]},
      {stage5_1[8]}
   );
   gpc1_1 gpc4861 (
      {stage4_1[14]},
      {stage5_1[9]}
   );
   gpc1_1 gpc4862 (
      {stage4_1[15]},
      {stage5_1[10]}
   );
   gpc1_1 gpc4863 (
      {stage4_2[5]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4864 (
      {stage4_2[6]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4865 (
      {stage4_2[7]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4866 (
      {stage4_2[8]},
      {stage5_2[5]}
   );
   gpc1_1 gpc4867 (
      {stage4_2[9]},
      {stage5_2[6]}
   );
   gpc1_1 gpc4868 (
      {stage4_2[10]},
      {stage5_2[7]}
   );
   gpc1_1 gpc4869 (
      {stage4_2[11]},
      {stage5_2[8]}
   );
   gpc1_1 gpc4870 (
      {stage4_2[12]},
      {stage5_2[9]}
   );
   gpc1_1 gpc4871 (
      {stage4_3[22]},
      {stage5_3[5]}
   );
   gpc1_1 gpc4872 (
      {stage4_4[21]},
      {stage5_4[7]}
   );
   gpc1_1 gpc4873 (
      {stage4_4[22]},
      {stage5_4[8]}
   );
   gpc1_1 gpc4874 (
      {stage4_4[23]},
      {stage5_4[9]}
   );
   gpc1_1 gpc4875 (
      {stage4_6[22]},
      {stage5_6[12]}
   );
   gpc1_1 gpc4876 (
      {stage4_7[8]},
      {stage5_7[13]}
   );
   gpc1_1 gpc4877 (
      {stage4_7[9]},
      {stage5_7[14]}
   );
   gpc1_1 gpc4878 (
      {stage4_7[10]},
      {stage5_7[15]}
   );
   gpc1_1 gpc4879 (
      {stage4_7[11]},
      {stage5_7[16]}
   );
   gpc1_1 gpc4880 (
      {stage4_7[12]},
      {stage5_7[17]}
   );
   gpc1_1 gpc4881 (
      {stage4_7[13]},
      {stage5_7[18]}
   );
   gpc1_1 gpc4882 (
      {stage4_7[14]},
      {stage5_7[19]}
   );
   gpc1_1 gpc4883 (
      {stage4_8[26]},
      {stage5_8[7]}
   );
   gpc1_1 gpc4884 (
      {stage4_8[27]},
      {stage5_8[8]}
   );
   gpc1_1 gpc4885 (
      {stage4_8[28]},
      {stage5_8[9]}
   );
   gpc1_1 gpc4886 (
      {stage4_11[38]},
      {stage5_11[11]}
   );
   gpc1_1 gpc4887 (
      {stage4_11[39]},
      {stage5_11[12]}
   );
   gpc1_1 gpc4888 (
      {stage4_11[40]},
      {stage5_11[13]}
   );
   gpc1_1 gpc4889 (
      {stage4_11[41]},
      {stage5_11[14]}
   );
   gpc1_1 gpc4890 (
      {stage4_11[42]},
      {stage5_11[15]}
   );
   gpc1_1 gpc4891 (
      {stage4_15[38]},
      {stage5_15[12]}
   );
   gpc1_1 gpc4892 (
      {stage4_16[19]},
      {stage5_16[14]}
   );
   gpc1_1 gpc4893 (
      {stage4_18[23]},
      {stage5_18[11]}
   );
   gpc1_1 gpc4894 (
      {stage4_18[24]},
      {stage5_18[12]}
   );
   gpc1_1 gpc4895 (
      {stage4_18[25]},
      {stage5_18[13]}
   );
   gpc1_1 gpc4896 (
      {stage4_18[26]},
      {stage5_18[14]}
   );
   gpc1_1 gpc4897 (
      {stage4_18[27]},
      {stage5_18[15]}
   );
   gpc1_1 gpc4898 (
      {stage4_18[28]},
      {stage5_18[16]}
   );
   gpc1_1 gpc4899 (
      {stage4_19[19]},
      {stage5_19[11]}
   );
   gpc1_1 gpc4900 (
      {stage4_19[20]},
      {stage5_19[12]}
   );
   gpc1_1 gpc4901 (
      {stage4_19[21]},
      {stage5_19[13]}
   );
   gpc1_1 gpc4902 (
      {stage4_19[22]},
      {stage5_19[14]}
   );
   gpc1_1 gpc4903 (
      {stage4_19[23]},
      {stage5_19[15]}
   );
   gpc1_1 gpc4904 (
      {stage4_19[24]},
      {stage5_19[16]}
   );
   gpc1_1 gpc4905 (
      {stage4_19[25]},
      {stage5_19[17]}
   );
   gpc1_1 gpc4906 (
      {stage4_19[26]},
      {stage5_19[18]}
   );
   gpc1_1 gpc4907 (
      {stage4_19[27]},
      {stage5_19[19]}
   );
   gpc1_1 gpc4908 (
      {stage4_19[28]},
      {stage5_19[20]}
   );
   gpc1_1 gpc4909 (
      {stage4_19[29]},
      {stage5_19[21]}
   );
   gpc1_1 gpc4910 (
      {stage4_19[30]},
      {stage5_19[22]}
   );
   gpc1_1 gpc4911 (
      {stage4_19[31]},
      {stage5_19[23]}
   );
   gpc1_1 gpc4912 (
      {stage4_20[12]},
      {stage5_20[7]}
   );
   gpc1_1 gpc4913 (
      {stage4_20[13]},
      {stage5_20[8]}
   );
   gpc1_1 gpc4914 (
      {stage4_20[14]},
      {stage5_20[9]}
   );
   gpc1_1 gpc4915 (
      {stage4_20[15]},
      {stage5_20[10]}
   );
   gpc1_1 gpc4916 (
      {stage4_20[16]},
      {stage5_20[11]}
   );
   gpc1_1 gpc4917 (
      {stage4_20[17]},
      {stage5_20[12]}
   );
   gpc1_1 gpc4918 (
      {stage4_20[18]},
      {stage5_20[13]}
   );
   gpc1_1 gpc4919 (
      {stage4_22[24]},
      {stage5_22[10]}
   );
   gpc1_1 gpc4920 (
      {stage4_22[25]},
      {stage5_22[11]}
   );
   gpc1_1 gpc4921 (
      {stage4_22[26]},
      {stage5_22[12]}
   );
   gpc1_1 gpc4922 (
      {stage4_22[27]},
      {stage5_22[13]}
   );
   gpc1_1 gpc4923 (
      {stage4_22[28]},
      {stage5_22[14]}
   );
   gpc1_1 gpc4924 (
      {stage4_22[29]},
      {stage5_22[15]}
   );
   gpc1_1 gpc4925 (
      {stage4_22[30]},
      {stage5_22[16]}
   );
   gpc1_1 gpc4926 (
      {stage4_24[26]},
      {stage5_24[10]}
   );
   gpc1_1 gpc4927 (
      {stage4_24[27]},
      {stage5_24[11]}
   );
   gpc1_1 gpc4928 (
      {stage4_24[28]},
      {stage5_24[12]}
   );
   gpc1_1 gpc4929 (
      {stage4_24[29]},
      {stage5_24[13]}
   );
   gpc1_1 gpc4930 (
      {stage4_25[18]},
      {stage5_25[11]}
   );
   gpc1_1 gpc4931 (
      {stage4_26[20]},
      {stage5_26[11]}
   );
   gpc1_1 gpc4932 (
      {stage4_26[21]},
      {stage5_26[12]}
   );
   gpc1_1 gpc4933 (
      {stage4_26[22]},
      {stage5_26[13]}
   );
   gpc1_1 gpc4934 (
      {stage4_27[22]},
      {stage5_27[9]}
   );
   gpc1_1 gpc4935 (
      {stage4_27[23]},
      {stage5_27[10]}
   );
   gpc1_1 gpc4936 (
      {stage4_27[24]},
      {stage5_27[11]}
   );
   gpc1_1 gpc4937 (
      {stage4_27[25]},
      {stage5_27[12]}
   );
   gpc1_1 gpc4938 (
      {stage4_27[26]},
      {stage5_27[13]}
   );
   gpc1_1 gpc4939 (
      {stage4_29[23]},
      {stage5_29[10]}
   );
   gpc1_1 gpc4940 (
      {stage4_29[24]},
      {stage5_29[11]}
   );
   gpc1_1 gpc4941 (
      {stage4_29[25]},
      {stage5_29[12]}
   );
   gpc1_1 gpc4942 (
      {stage4_30[23]},
      {stage5_30[13]}
   );
   gpc1_1 gpc4943 (
      {stage4_30[24]},
      {stage5_30[14]}
   );
   gpc1_1 gpc4944 (
      {stage4_30[25]},
      {stage5_30[15]}
   );
   gpc1_1 gpc4945 (
      {stage4_30[26]},
      {stage5_30[16]}
   );
   gpc1_1 gpc4946 (
      {stage4_31[27]},
      {stage5_31[9]}
   );
   gpc1_1 gpc4947 (
      {stage4_31[28]},
      {stage5_31[10]}
   );
   gpc1_1 gpc4948 (
      {stage4_31[29]},
      {stage5_31[11]}
   );
   gpc1_1 gpc4949 (
      {stage4_31[30]},
      {stage5_31[12]}
   );
   gpc1_1 gpc4950 (
      {stage4_32[25]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4951 (
      {stage4_32[26]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4952 (
      {stage4_32[27]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4953 (
      {stage4_32[28]},
      {stage5_32[11]}
   );
   gpc1_1 gpc4954 (
      {stage4_32[29]},
      {stage5_32[12]}
   );
   gpc1_1 gpc4955 (
      {stage4_32[30]},
      {stage5_32[13]}
   );
   gpc1_1 gpc4956 (
      {stage4_32[31]},
      {stage5_32[14]}
   );
   gpc1_1 gpc4957 (
      {stage4_32[32]},
      {stage5_32[15]}
   );
   gpc1_1 gpc4958 (
      {stage4_32[33]},
      {stage5_32[16]}
   );
   gpc1_1 gpc4959 (
      {stage4_32[34]},
      {stage5_32[17]}
   );
   gpc1_1 gpc4960 (
      {stage4_32[35]},
      {stage5_32[18]}
   );
   gpc1_1 gpc4961 (
      {stage4_32[36]},
      {stage5_32[19]}
   );
   gpc1_1 gpc4962 (
      {stage4_32[37]},
      {stage5_32[20]}
   );
   gpc1_1 gpc4963 (
      {stage4_32[38]},
      {stage5_32[21]}
   );
   gpc1_1 gpc4964 (
      {stage4_32[39]},
      {stage5_32[22]}
   );
   gpc1_1 gpc4965 (
      {stage4_32[40]},
      {stage5_32[23]}
   );
   gpc1_1 gpc4966 (
      {stage4_32[41]},
      {stage5_32[24]}
   );
   gpc1_1 gpc4967 (
      {stage4_32[42]},
      {stage5_32[25]}
   );
   gpc1_1 gpc4968 (
      {stage4_33[18]},
      {stage5_33[10]}
   );
   gpc1_1 gpc4969 (
      {stage4_34[12]},
      {stage5_34[9]}
   );
   gpc1_1 gpc4970 (
      {stage4_35[12]},
      {stage5_35[5]}
   );
   gpc1_1 gpc4971 (
      {stage4_35[13]},
      {stage5_35[6]}
   );
   gpc1_1 gpc4972 (
      {stage4_35[14]},
      {stage5_35[7]}
   );
   gpc1_1 gpc4973 (
      {stage4_37[0]},
      {stage5_37[4]}
   );
   gpc1_1 gpc4974 (
      {stage4_37[1]},
      {stage5_37[5]}
   );
   gpc1_1 gpc4975 (
      {stage4_37[2]},
      {stage5_37[6]}
   );
   gpc1343_5 gpc4976 (
      {stage5_0[0], stage5_0[1], stage5_0[2]},
      {stage5_1[0], stage5_1[1], stage5_1[2], stage5_1[3]},
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc1343_5 gpc4977 (
      {stage5_0[3], stage5_0[4], stage5_0[5]},
      {stage5_1[4], stage5_1[5], stage5_1[6], stage5_1[7]},
      {stage5_2[3], stage5_2[4], stage5_2[5]},
      {stage5_3[1]},
      {stage6_4[1],stage6_3[1],stage6_2[1],stage6_1[1],stage6_0[1]}
   );
   gpc117_4 gpc4978 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6]},
      {stage5_5[0]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[2]}
   );
   gpc1343_5 gpc4979 (
      {stage5_5[1], stage5_5[2], stage5_5[3]},
      {stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc4980 (
      {stage5_5[4], stage5_5[5], stage5_5[6]},
      {stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8]},
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[1]},
      {stage6_9[1],stage6_8[1],stage6_7[2],stage6_6[2],stage6_5[2]}
   );
   gpc1343_5 gpc4981 (
      {stage5_5[7], stage5_5[8], stage5_5[9]},
      {stage5_6[9], stage5_6[10], stage5_6[11], stage5_6[12]},
      {stage5_7[6], stage5_7[7], stage5_7[8]},
      {stage5_8[2]},
      {stage6_9[2],stage6_8[2],stage6_7[3],stage6_6[3],stage6_5[3]}
   );
   gpc606_5 gpc4982 (
      {stage5_7[9], stage5_7[10], stage5_7[11], stage5_7[12], stage5_7[13], stage5_7[14]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[3],stage6_8[3],stage6_7[4]}
   );
   gpc615_5 gpc4983 (
      {stage5_7[15], stage5_7[16], stage5_7[17], stage5_7[18], stage5_7[19]},
      {stage5_8[3]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], 1'b0},
      {stage6_11[1],stage6_10[1],stage6_9[4],stage6_8[4],stage6_7[5]}
   );
   gpc606_5 gpc4984 (
      {stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[2],stage6_10[2],stage6_9[5],stage6_8[5]}
   );
   gpc7_3 gpc4985 (
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11], stage5_10[12]},
      {stage6_12[1],stage6_11[3],stage6_10[3]}
   );
   gpc207_4 gpc4986 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6]},
      {stage5_13[0], stage5_13[1]},
      {stage6_14[0],stage6_13[0],stage6_12[2],stage6_11[4]}
   );
   gpc207_4 gpc4987 (
      {stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11], stage5_11[12], stage5_11[13]},
      {stage5_13[2], stage5_13[3]},
      {stage6_14[1],stage6_13[1],stage6_12[3],stage6_11[5]}
   );
   gpc7_3 gpc4988 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[2],stage6_13[2],stage6_12[4]}
   );
   gpc623_5 gpc4989 (
      {stage5_12[7], stage5_12[8], stage5_12[9]},
      {stage5_13[4], stage5_13[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage6_16[0],stage6_15[0],stage6_14[3],stage6_13[3],stage6_12[5]}
   );
   gpc623_5 gpc4990 (
      {stage5_13[6], stage5_13[7], stage5_13[8]},
      {stage5_14[6], stage5_14[7]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[4],stage6_13[4]}
   );
   gpc623_5 gpc4991 (
      {stage5_13[9], stage5_13[10], stage5_13[11]},
      {stage5_14[8], stage5_14[9]},
      {stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9], stage5_15[10], stage5_15[11]},
      {stage6_17[1],stage6_16[2],stage6_15[2],stage6_14[5],stage6_13[5]}
   );
   gpc207_4 gpc4992 (
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6]},
      {stage5_18[0], stage5_18[1]},
      {stage6_19[0],stage6_18[0],stage6_17[2],stage6_16[3]}
   );
   gpc207_4 gpc4993 (
      {stage5_16[7], stage5_16[8], stage5_16[9], stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13]},
      {stage5_18[2], stage5_18[3]},
      {stage6_19[1],stage6_18[1],stage6_17[3],stage6_16[4]}
   );
   gpc1163_5 gpc4994 (
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[4], stage5_18[5], stage5_18[6], stage5_18[7], stage5_18[8], stage5_18[9]},
      {stage5_19[0]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[2],stage6_18[2],stage6_17[4]}
   );
   gpc1163_5 gpc4995 (
      {stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_18[10], stage5_18[11], stage5_18[12], stage5_18[13], stage5_18[14], stage5_18[15]},
      {stage5_19[1]},
      {stage5_20[1]},
      {stage6_21[1],stage6_20[1],stage6_19[3],stage6_18[3],stage6_17[5]}
   );
   gpc606_5 gpc4996 (
      {stage5_17[6], stage5_17[7], stage5_17[8], stage5_17[9], stage5_17[10], stage5_17[11]},
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6], stage5_19[7]},
      {stage6_21[2],stage6_20[2],stage6_19[4],stage6_18[4],stage6_17[6]}
   );
   gpc207_4 gpc4997 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12], stage5_19[13], stage5_19[14]},
      {stage5_21[0], stage5_21[1]},
      {stage6_22[0],stage6_21[3],stage6_20[3],stage6_19[5]}
   );
   gpc606_5 gpc4998 (
      {stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7]},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[0],stage6_22[1],stage6_21[4],stage6_20[4]}
   );
   gpc606_5 gpc4999 (
      {stage5_20[8], stage5_20[9], stage5_20[10], stage5_20[11], stage5_20[12], stage5_20[13]},
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10], stage5_22[11]},
      {stage6_24[1],stage6_23[1],stage6_22[2],stage6_21[5],stage6_20[5]}
   );
   gpc1415_5 gpc5000 (
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4]},
      {stage5_24[0]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[0],stage6_24[2],stage6_23[2]}
   );
   gpc615_5 gpc5001 (
      {stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8], stage5_23[9]},
      {stage5_24[1]},
      {stage5_25[4], stage5_25[5], stage5_25[6], stage5_25[7], stage5_25[8], stage5_25[9]},
      {stage6_27[1],stage6_26[1],stage6_25[1],stage6_24[3],stage6_23[3]}
   );
   gpc606_5 gpc5002 (
      {stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6], stage5_24[7]},
      {stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5], stage5_26[6]},
      {stage6_28[0],stage6_27[2],stage6_26[2],stage6_25[2],stage6_24[4]}
   );
   gpc606_5 gpc5003 (
      {stage5_24[8], stage5_24[9], stage5_24[10], stage5_24[11], stage5_24[12], stage5_24[13]},
      {stage5_26[7], stage5_26[8], stage5_26[9], stage5_26[10], stage5_26[11], stage5_26[12]},
      {stage6_28[1],stage6_27[3],stage6_26[3],stage6_25[3],stage6_24[5]}
   );
   gpc606_5 gpc5004 (
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4], stage5_27[5]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[0],stage6_28[2],stage6_27[4]}
   );
   gpc606_5 gpc5005 (
      {stage5_27[6], stage5_27[7], stage5_27[8], stage5_27[9], stage5_27[10], stage5_27[11]},
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage6_31[1],stage6_30[1],stage6_29[1],stage6_28[3],stage6_27[5]}
   );
   gpc207_4 gpc5006 (
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], stage5_28[5], stage5_28[6]},
      {stage5_30[0], stage5_30[1]},
      {stage6_31[2],stage6_30[2],stage6_29[2],stage6_28[4]}
   );
   gpc615_5 gpc5007 (
      {stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage5_31[0]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage6_34[0],stage6_33[0],stage6_32[0],stage6_31[3],stage6_30[3]}
   );
   gpc615_5 gpc5008 (
      {stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10], stage5_30[11]},
      {stage5_31[1]},
      {stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9], stage5_32[10], stage5_32[11]},
      {stage6_34[1],stage6_33[1],stage6_32[1],stage6_31[4],stage6_30[4]}
   );
   gpc615_5 gpc5009 (
      {stage5_30[12], stage5_30[13], stage5_30[14], stage5_30[15], stage5_30[16]},
      {stage5_31[2]},
      {stage5_32[12], stage5_32[13], stage5_32[14], stage5_32[15], stage5_32[16], stage5_32[17]},
      {stage6_34[2],stage6_33[2],stage6_32[2],stage6_31[5],stage6_30[5]}
   );
   gpc615_5 gpc5010 (
      {stage5_31[3], stage5_31[4], stage5_31[5], stage5_31[6], stage5_31[7]},
      {stage5_32[18]},
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5]},
      {stage6_35[0],stage6_34[3],stage6_33[3],stage6_32[3],stage6_31[6]}
   );
   gpc615_5 gpc5011 (
      {stage5_31[8], stage5_31[9], stage5_31[10], stage5_31[11], stage5_31[12]},
      {stage5_32[19]},
      {stage5_33[6], stage5_33[7], stage5_33[8], stage5_33[9], stage5_33[10], 1'b0},
      {stage6_35[1],stage6_34[4],stage6_33[4],stage6_32[4],stage6_31[7]}
   );
   gpc606_5 gpc5012 (
      {stage5_32[20], stage5_32[21], stage5_32[22], stage5_32[23], stage5_32[24], stage5_32[25]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[2],stage6_34[5],stage6_33[5],stage6_32[5]}
   );
   gpc606_5 gpc5013 (
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[0],stage6_36[1],stage6_35[3]}
   );
   gpc1325_5 gpc5014 (
      {stage5_36[0], stage5_36[1], stage5_36[2], stage5_36[3], 1'b0},
      {stage5_37[6], 1'b0},
      {stage5_38[0], stage5_38[1], 1'b0},
      {1'b0},
      {stage6_40[0],stage6_39[1],stage6_38[1],stage6_37[1],stage6_36[2]}
   );
   gpc1_1 gpc5015 (
      {stage5_0[6]},
      {stage6_0[2]}
   );
   gpc1_1 gpc5016 (
      {stage5_0[7]},
      {stage6_0[3]}
   );
   gpc1_1 gpc5017 (
      {stage5_0[8]},
      {stage6_0[4]}
   );
   gpc1_1 gpc5018 (
      {stage5_0[9]},
      {stage6_0[5]}
   );
   gpc1_1 gpc5019 (
      {stage5_0[10]},
      {stage6_0[6]}
   );
   gpc1_1 gpc5020 (
      {stage5_1[8]},
      {stage6_1[2]}
   );
   gpc1_1 gpc5021 (
      {stage5_1[9]},
      {stage6_1[3]}
   );
   gpc1_1 gpc5022 (
      {stage5_1[10]},
      {stage6_1[4]}
   );
   gpc1_1 gpc5023 (
      {stage5_2[6]},
      {stage6_2[2]}
   );
   gpc1_1 gpc5024 (
      {stage5_2[7]},
      {stage6_2[3]}
   );
   gpc1_1 gpc5025 (
      {stage5_2[8]},
      {stage6_2[4]}
   );
   gpc1_1 gpc5026 (
      {stage5_2[9]},
      {stage6_2[5]}
   );
   gpc1_1 gpc5027 (
      {stage5_3[2]},
      {stage6_3[2]}
   );
   gpc1_1 gpc5028 (
      {stage5_3[3]},
      {stage6_3[3]}
   );
   gpc1_1 gpc5029 (
      {stage5_3[4]},
      {stage6_3[4]}
   );
   gpc1_1 gpc5030 (
      {stage5_3[5]},
      {stage6_3[5]}
   );
   gpc1_1 gpc5031 (
      {stage5_4[7]},
      {stage6_4[3]}
   );
   gpc1_1 gpc5032 (
      {stage5_4[8]},
      {stage6_4[4]}
   );
   gpc1_1 gpc5033 (
      {stage5_4[9]},
      {stage6_4[5]}
   );
   gpc1_1 gpc5034 (
      {stage5_5[10]},
      {stage6_5[4]}
   );
   gpc1_1 gpc5035 (
      {stage5_11[14]},
      {stage6_11[6]}
   );
   gpc1_1 gpc5036 (
      {stage5_11[15]},
      {stage6_11[7]}
   );
   gpc1_1 gpc5037 (
      {stage5_12[10]},
      {stage6_12[6]}
   );
   gpc1_1 gpc5038 (
      {stage5_13[12]},
      {stage6_13[6]}
   );
   gpc1_1 gpc5039 (
      {stage5_13[13]},
      {stage6_13[7]}
   );
   gpc1_1 gpc5040 (
      {stage5_13[14]},
      {stage6_13[8]}
   );
   gpc1_1 gpc5041 (
      {stage5_15[12]},
      {stage6_15[3]}
   );
   gpc1_1 gpc5042 (
      {stage5_16[14]},
      {stage6_16[5]}
   );
   gpc1_1 gpc5043 (
      {stage5_17[12]},
      {stage6_17[7]}
   );
   gpc1_1 gpc5044 (
      {stage5_17[13]},
      {stage6_17[8]}
   );
   gpc1_1 gpc5045 (
      {stage5_17[14]},
      {stage6_17[9]}
   );
   gpc1_1 gpc5046 (
      {stage5_18[16]},
      {stage6_18[5]}
   );
   gpc1_1 gpc5047 (
      {stage5_19[15]},
      {stage6_19[6]}
   );
   gpc1_1 gpc5048 (
      {stage5_19[16]},
      {stage6_19[7]}
   );
   gpc1_1 gpc5049 (
      {stage5_19[17]},
      {stage6_19[8]}
   );
   gpc1_1 gpc5050 (
      {stage5_19[18]},
      {stage6_19[9]}
   );
   gpc1_1 gpc5051 (
      {stage5_19[19]},
      {stage6_19[10]}
   );
   gpc1_1 gpc5052 (
      {stage5_19[20]},
      {stage6_19[11]}
   );
   gpc1_1 gpc5053 (
      {stage5_19[21]},
      {stage6_19[12]}
   );
   gpc1_1 gpc5054 (
      {stage5_19[22]},
      {stage6_19[13]}
   );
   gpc1_1 gpc5055 (
      {stage5_19[23]},
      {stage6_19[14]}
   );
   gpc1_1 gpc5056 (
      {stage5_21[2]},
      {stage6_21[6]}
   );
   gpc1_1 gpc5057 (
      {stage5_21[3]},
      {stage6_21[7]}
   );
   gpc1_1 gpc5058 (
      {stage5_21[4]},
      {stage6_21[8]}
   );
   gpc1_1 gpc5059 (
      {stage5_21[5]},
      {stage6_21[9]}
   );
   gpc1_1 gpc5060 (
      {stage5_21[6]},
      {stage6_21[10]}
   );
   gpc1_1 gpc5061 (
      {stage5_21[7]},
      {stage6_21[11]}
   );
   gpc1_1 gpc5062 (
      {stage5_21[8]},
      {stage6_21[12]}
   );
   gpc1_1 gpc5063 (
      {stage5_22[12]},
      {stage6_22[3]}
   );
   gpc1_1 gpc5064 (
      {stage5_22[13]},
      {stage6_22[4]}
   );
   gpc1_1 gpc5065 (
      {stage5_22[14]},
      {stage6_22[5]}
   );
   gpc1_1 gpc5066 (
      {stage5_22[15]},
      {stage6_22[6]}
   );
   gpc1_1 gpc5067 (
      {stage5_22[16]},
      {stage6_22[7]}
   );
   gpc1_1 gpc5068 (
      {stage5_25[10]},
      {stage6_25[4]}
   );
   gpc1_1 gpc5069 (
      {stage5_25[11]},
      {stage6_25[5]}
   );
   gpc1_1 gpc5070 (
      {stage5_26[13]},
      {stage6_26[4]}
   );
   gpc1_1 gpc5071 (
      {stage5_27[12]},
      {stage6_27[6]}
   );
   gpc1_1 gpc5072 (
      {stage5_27[13]},
      {stage6_27[7]}
   );
   gpc1_1 gpc5073 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc5074 (
      {stage5_34[6]},
      {stage6_34[6]}
   );
   gpc1_1 gpc5075 (
      {stage5_34[7]},
      {stage6_34[7]}
   );
   gpc1_1 gpc5076 (
      {stage5_34[8]},
      {stage6_34[8]}
   );
   gpc1_1 gpc5077 (
      {stage5_34[9]},
      {stage6_34[9]}
   );
   gpc1_1 gpc5078 (
      {stage5_35[6]},
      {stage6_35[4]}
   );
   gpc1_1 gpc5079 (
      {stage5_35[7]},
      {stage6_35[5]}
   );
   gpc606_5 gpc5080 (
      {stage6_1[0], stage6_1[1], stage6_1[2], stage6_1[3], stage6_1[4], 1'b0},
      {stage6_3[0], stage6_3[1], stage6_3[2], stage6_3[3], stage6_3[4], stage6_3[5]},
      {stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0]}
   );
   gpc15_3 gpc5081 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], stage6_5[4]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[1]}
   );
   gpc606_5 gpc5082 (
      {stage6_7[0], stage6_7[1], stage6_7[2], stage6_7[3], stage6_7[4], stage6_7[5]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc1343_5 gpc5083 (
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3]},
      {stage6_13[0], stage6_13[1], stage6_13[2]},
      {stage6_14[0]},
      {stage7_15[0],stage7_14[0],stage7_13[0],stage7_12[0],stage7_11[1]}
   );
   gpc615_5 gpc5084 (
      {stage6_11[3], stage6_11[4], stage6_11[5], stage6_11[6], stage6_11[7]},
      {stage6_12[4]},
      {stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6], stage6_13[7], stage6_13[8]},
      {stage7_15[1],stage7_14[1],stage7_13[1],stage7_12[1],stage7_11[2]}
   );
   gpc1343_5 gpc5085 (
      {stage6_16[0], stage6_16[1], stage6_16[2]},
      {stage6_17[0], stage6_17[1], stage6_17[2], stage6_17[3]},
      {stage6_18[0], stage6_18[1], stage6_18[2]},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[0]}
   );
   gpc1343_5 gpc5086 (
      {stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage6_17[4], stage6_17[5], stage6_17[6], stage6_17[7]},
      {stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_19[1]},
      {stage7_20[1],stage7_19[1],stage7_18[1],stage7_17[1],stage7_16[1]}
   );
   gpc606_5 gpc5087 (
      {stage6_19[2], stage6_19[3], stage6_19[4], stage6_19[5], stage6_19[6], stage6_19[7]},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[2],stage7_19[2]}
   );
   gpc606_5 gpc5088 (
      {stage6_19[8], stage6_19[9], stage6_19[10], stage6_19[11], stage6_19[12], stage6_19[13]},
      {stage6_21[6], stage6_21[7], stage6_21[8], stage6_21[9], stage6_21[10], stage6_21[11]},
      {stage7_23[1],stage7_22[1],stage7_21[1],stage7_20[3],stage7_19[3]}
   );
   gpc15_3 gpc5089 (
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[12]},
      {stage7_22[2],stage7_21[2],stage7_20[4]}
   );
   gpc606_5 gpc5090 (
      {stage6_22[0], stage6_22[1], stage6_22[2], stage6_22[3], stage6_22[4], stage6_22[5]},
      {stage6_24[0], stage6_24[1], stage6_24[2], stage6_24[3], stage6_24[4], stage6_24[5]},
      {stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[2],stage7_22[3]}
   );
   gpc606_5 gpc5091 (
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], stage6_25[5]},
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], stage6_27[5]},
      {stage7_29[0],stage7_28[0],stage7_27[0],stage7_26[1],stage7_25[1]}
   );
   gpc15_3 gpc5092 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4]},
      {stage6_27[6]},
      {stage7_28[1],stage7_27[1],stage7_26[2]}
   );
   gpc606_5 gpc5093 (
      {stage6_30[0], stage6_30[1], stage6_30[2], stage6_30[3], stage6_30[4], stage6_30[5]},
      {stage6_32[0], stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[0]}
   );
   gpc606_5 gpc5094 (
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage6_35[0], stage6_35[1], stage6_35[2], stage6_35[3], stage6_35[4], stage6_35[5]},
      {stage7_37[0],stage7_36[0],stage7_35[0],stage7_34[1],stage7_33[1]}
   );
   gpc606_5 gpc5095 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4], stage6_34[5]},
      {stage6_36[0], stage6_36[1], stage6_36[2], 1'b0, 1'b0, 1'b0},
      {stage7_38[0],stage7_37[1],stage7_36[1],stage7_35[1],stage7_34[2]}
   );
   gpc1_1 gpc5096 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc5097 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc5098 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc5099 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc5100 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc5101 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc5102 (
      {stage6_0[6]},
      {stage7_0[6]}
   );
   gpc1_1 gpc5103 (
      {stage6_2[0]},
      {stage7_2[1]}
   );
   gpc1_1 gpc5104 (
      {stage6_2[1]},
      {stage7_2[2]}
   );
   gpc1_1 gpc5105 (
      {stage6_2[2]},
      {stage7_2[3]}
   );
   gpc1_1 gpc5106 (
      {stage6_2[3]},
      {stage7_2[4]}
   );
   gpc1_1 gpc5107 (
      {stage6_2[4]},
      {stage7_2[5]}
   );
   gpc1_1 gpc5108 (
      {stage6_2[5]},
      {stage7_2[6]}
   );
   gpc1_1 gpc5109 (
      {stage6_4[0]},
      {stage7_4[1]}
   );
   gpc1_1 gpc5110 (
      {stage6_4[1]},
      {stage7_4[2]}
   );
   gpc1_1 gpc5111 (
      {stage6_4[2]},
      {stage7_4[3]}
   );
   gpc1_1 gpc5112 (
      {stage6_4[3]},
      {stage7_4[4]}
   );
   gpc1_1 gpc5113 (
      {stage6_4[4]},
      {stage7_4[5]}
   );
   gpc1_1 gpc5114 (
      {stage6_4[5]},
      {stage7_4[6]}
   );
   gpc1_1 gpc5115 (
      {stage6_6[1]},
      {stage7_6[1]}
   );
   gpc1_1 gpc5116 (
      {stage6_6[2]},
      {stage7_6[2]}
   );
   gpc1_1 gpc5117 (
      {stage6_6[3]},
      {stage7_6[3]}
   );
   gpc1_1 gpc5118 (
      {stage6_8[0]},
      {stage7_8[1]}
   );
   gpc1_1 gpc5119 (
      {stage6_8[1]},
      {stage7_8[2]}
   );
   gpc1_1 gpc5120 (
      {stage6_8[2]},
      {stage7_8[3]}
   );
   gpc1_1 gpc5121 (
      {stage6_8[3]},
      {stage7_8[4]}
   );
   gpc1_1 gpc5122 (
      {stage6_8[4]},
      {stage7_8[5]}
   );
   gpc1_1 gpc5123 (
      {stage6_8[5]},
      {stage7_8[6]}
   );
   gpc1_1 gpc5124 (
      {stage6_10[0]},
      {stage7_10[1]}
   );
   gpc1_1 gpc5125 (
      {stage6_10[1]},
      {stage7_10[2]}
   );
   gpc1_1 gpc5126 (
      {stage6_10[2]},
      {stage7_10[3]}
   );
   gpc1_1 gpc5127 (
      {stage6_10[3]},
      {stage7_10[4]}
   );
   gpc1_1 gpc5128 (
      {stage6_12[5]},
      {stage7_12[2]}
   );
   gpc1_1 gpc5129 (
      {stage6_12[6]},
      {stage7_12[3]}
   );
   gpc1_1 gpc5130 (
      {stage6_14[1]},
      {stage7_14[2]}
   );
   gpc1_1 gpc5131 (
      {stage6_14[2]},
      {stage7_14[3]}
   );
   gpc1_1 gpc5132 (
      {stage6_14[3]},
      {stage7_14[4]}
   );
   gpc1_1 gpc5133 (
      {stage6_14[4]},
      {stage7_14[5]}
   );
   gpc1_1 gpc5134 (
      {stage6_14[5]},
      {stage7_14[6]}
   );
   gpc1_1 gpc5135 (
      {stage6_15[0]},
      {stage7_15[2]}
   );
   gpc1_1 gpc5136 (
      {stage6_15[1]},
      {stage7_15[3]}
   );
   gpc1_1 gpc5137 (
      {stage6_15[2]},
      {stage7_15[4]}
   );
   gpc1_1 gpc5138 (
      {stage6_15[3]},
      {stage7_15[5]}
   );
   gpc1_1 gpc5139 (
      {stage6_17[8]},
      {stage7_17[2]}
   );
   gpc1_1 gpc5140 (
      {stage6_17[9]},
      {stage7_17[3]}
   );
   gpc1_1 gpc5141 (
      {stage6_19[14]},
      {stage7_19[4]}
   );
   gpc1_1 gpc5142 (
      {stage6_20[5]},
      {stage7_20[5]}
   );
   gpc1_1 gpc5143 (
      {stage6_22[6]},
      {stage7_22[4]}
   );
   gpc1_1 gpc5144 (
      {stage6_22[7]},
      {stage7_22[5]}
   );
   gpc1_1 gpc5145 (
      {stage6_23[0]},
      {stage7_23[3]}
   );
   gpc1_1 gpc5146 (
      {stage6_23[1]},
      {stage7_23[4]}
   );
   gpc1_1 gpc5147 (
      {stage6_23[2]},
      {stage7_23[5]}
   );
   gpc1_1 gpc5148 (
      {stage6_23[3]},
      {stage7_23[6]}
   );
   gpc1_1 gpc5149 (
      {stage6_27[7]},
      {stage7_27[2]}
   );
   gpc1_1 gpc5150 (
      {stage6_28[0]},
      {stage7_28[2]}
   );
   gpc1_1 gpc5151 (
      {stage6_28[1]},
      {stage7_28[3]}
   );
   gpc1_1 gpc5152 (
      {stage6_28[2]},
      {stage7_28[4]}
   );
   gpc1_1 gpc5153 (
      {stage6_28[3]},
      {stage7_28[5]}
   );
   gpc1_1 gpc5154 (
      {stage6_28[4]},
      {stage7_28[6]}
   );
   gpc1_1 gpc5155 (
      {stage6_29[0]},
      {stage7_29[1]}
   );
   gpc1_1 gpc5156 (
      {stage6_29[1]},
      {stage7_29[2]}
   );
   gpc1_1 gpc5157 (
      {stage6_29[2]},
      {stage7_29[3]}
   );
   gpc1_1 gpc5158 (
      {stage6_29[3]},
      {stage7_29[4]}
   );
   gpc1_1 gpc5159 (
      {stage6_31[0]},
      {stage7_31[1]}
   );
   gpc1_1 gpc5160 (
      {stage6_31[1]},
      {stage7_31[2]}
   );
   gpc1_1 gpc5161 (
      {stage6_31[2]},
      {stage7_31[3]}
   );
   gpc1_1 gpc5162 (
      {stage6_31[3]},
      {stage7_31[4]}
   );
   gpc1_1 gpc5163 (
      {stage6_31[4]},
      {stage7_31[5]}
   );
   gpc1_1 gpc5164 (
      {stage6_31[5]},
      {stage7_31[6]}
   );
   gpc1_1 gpc5165 (
      {stage6_31[6]},
      {stage7_31[7]}
   );
   gpc1_1 gpc5166 (
      {stage6_31[7]},
      {stage7_31[8]}
   );
   gpc1_1 gpc5167 (
      {stage6_34[6]},
      {stage7_34[3]}
   );
   gpc1_1 gpc5168 (
      {stage6_34[7]},
      {stage7_34[4]}
   );
   gpc1_1 gpc5169 (
      {stage6_34[8]},
      {stage7_34[5]}
   );
   gpc1_1 gpc5170 (
      {stage6_34[9]},
      {stage7_34[6]}
   );
   gpc1_1 gpc5171 (
      {stage6_37[0]},
      {stage7_37[2]}
   );
   gpc1_1 gpc5172 (
      {stage6_37[1]},
      {stage7_37[3]}
   );
   gpc1_1 gpc5173 (
      {stage6_38[0]},
      {stage7_38[1]}
   );
   gpc1_1 gpc5174 (
      {stage6_38[1]},
      {stage7_38[2]}
   );
   gpc1_1 gpc5175 (
      {stage6_39[0]},
      {stage7_39[0]}
   );
   gpc1_1 gpc5176 (
      {stage6_39[1]},
      {stage7_39[1]}
   );
   gpc1_1 gpc5177 (
      {stage6_40[0]},
      {stage7_40[0]}
   );
   gpc606_5 gpc5178 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4], stage7_0[5]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3], stage7_2[4], stage7_2[5]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc117_4 gpc5179 (
      {stage7_4[0], stage7_4[1], stage7_4[2], stage7_4[3], stage7_4[4], stage7_4[5], stage7_4[6]},
      {stage7_5[0]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1]}
   );
   gpc623_5 gpc5180 (
      {stage7_6[1], stage7_6[2], stage7_6[3]},
      {stage7_7[0], stage7_7[1]},
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4], stage7_8[5]},
      {stage8_10[0],stage8_9[0],stage8_8[0],stage8_7[1],stage8_6[1]}
   );
   gpc1325_5 gpc5181 (
      {stage7_10[0], stage7_10[1], stage7_10[2], stage7_10[3], stage7_10[4]},
      {stage7_11[0], stage7_11[1]},
      {stage7_12[0], stage7_12[1], stage7_12[2]},
      {stage7_13[0]},
      {stage8_14[0],stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[1]}
   );
   gpc117_4 gpc5182 (
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3], stage7_14[4], stage7_14[5], stage7_14[6]},
      {stage7_15[0]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[1]}
   );
   gpc1415_5 gpc5183 (
      {stage7_15[1], stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[1]},
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3]},
      {stage7_18[0]},
      {stage8_19[0],stage8_18[0],stage8_17[1],stage8_16[1],stage8_15[1]}
   );
   gpc135_4 gpc5184 (
      {stage7_19[0], stage7_19[1], stage7_19[2], stage7_19[3], stage7_19[4]},
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0]},
      {stage8_22[0],stage8_21[0],stage8_20[0],stage8_19[1]}
   );
   gpc623_5 gpc5185 (
      {stage7_20[3], stage7_20[4], stage7_20[5]},
      {stage7_21[1], stage7_21[2]},
      {stage7_22[0], stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5]},
      {stage8_24[0],stage8_23[0],stage8_22[1],stage8_21[1],stage8_20[1]}
   );
   gpc117_4 gpc5186 (
      {stage7_23[0], stage7_23[1], stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5], stage7_23[6]},
      {stage7_24[0]},
      {stage7_25[0]},
      {stage8_26[0],stage8_25[0],stage8_24[1],stage8_23[1]}
   );
   gpc2223_5 gpc5187 (
      {stage7_26[0], stage7_26[1], stage7_26[2]},
      {stage7_27[0], stage7_27[1]},
      {stage7_28[0], stage7_28[1]},
      {stage7_29[0], stage7_29[1]},
      {stage8_30[0],stage8_29[0],stage8_28[0],stage8_27[0],stage8_26[1]}
   );
   gpc2135_5 gpc5188 (
      {stage7_28[2], stage7_28[3], stage7_28[4], stage7_28[5], stage7_28[6]},
      {stage7_29[2], stage7_29[3], stage7_29[4]},
      {stage7_30[0]},
      {stage7_31[0], stage7_31[1]},
      {stage8_32[0],stage8_31[0],stage8_30[1],stage8_29[1],stage8_28[1]}
   );
   gpc117_4 gpc5189 (
      {stage7_31[2], stage7_31[3], stage7_31[4], stage7_31[5], stage7_31[6], stage7_31[7], stage7_31[8]},
      {stage7_32[0]},
      {stage7_33[0]},
      {stage8_34[0],stage8_33[0],stage8_32[1],stage8_31[1]}
   );
   gpc117_4 gpc5190 (
      {stage7_34[0], stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], stage7_34[6]},
      {stage7_35[0]},
      {stage7_36[0]},
      {stage8_37[0],stage8_36[0],stage8_35[0],stage8_34[1]}
   );
   gpc615_5 gpc5191 (
      {stage7_35[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_36[1]},
      {stage7_37[0], stage7_37[1], stage7_37[2], stage7_37[3], 1'b0, 1'b0},
      {stage8_39[0],stage8_38[0],stage8_37[1],stage8_36[1],stage8_35[1]}
   );
   gpc1163_5 gpc5192 (
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage7_39[0], stage7_39[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_40[0]},
      {1'b0},
      {stage8_40[0],stage8_39[1],stage8_38[1]}
   );
   gpc1_1 gpc5193 (
      {stage7_0[6]},
      {stage8_0[1]}
   );
   gpc1_1 gpc5194 (
      {stage7_1[0]},
      {stage8_1[1]}
   );
   gpc1_1 gpc5195 (
      {stage7_2[6]},
      {stage8_2[1]}
   );
   gpc1_1 gpc5196 (
      {stage7_3[0]},
      {stage8_3[1]}
   );
   gpc1_1 gpc5197 (
      {stage7_5[1]},
      {stage8_5[1]}
   );
   gpc1_1 gpc5198 (
      {stage7_8[6]},
      {stage8_8[1]}
   );
   gpc1_1 gpc5199 (
      {stage7_9[0]},
      {stage8_9[1]}
   );
   gpc1_1 gpc5200 (
      {stage7_11[2]},
      {stage8_11[1]}
   );
   gpc1_1 gpc5201 (
      {stage7_12[3]},
      {stage8_12[1]}
   );
   gpc1_1 gpc5202 (
      {stage7_13[1]},
      {stage8_13[1]}
   );
   gpc1_1 gpc5203 (
      {stage7_18[1]},
      {stage8_18[1]}
   );
   gpc1_1 gpc5204 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc5205 (
      {stage7_27[2]},
      {stage8_27[1]}
   );
   gpc1_1 gpc5206 (
      {stage7_33[1]},
      {stage8_33[1]}
   );
endmodule

module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    reg [511:0] src16;
    reg [511:0] src17;
    reg [511:0] src18;
    reg [511:0] src19;
    reg [511:0] src20;
    reg [511:0] src21;
    reg [511:0] src22;
    reg [511:0] src23;
    reg [511:0] src24;
    reg [511:0] src25;
    reg [511:0] src26;
    reg [511:0] src27;
    reg [511:0] src28;
    reg [511:0] src29;
    reg [511:0] src30;
    reg [511:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [40:0] srcsum;
    wire [40:0] dstsum;
    wire test;
    compressor_CLA512_32 compressor_CLA512_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485] + src16[486] + src16[487] + src16[488] + src16[489] + src16[490] + src16[491] + src16[492] + src16[493] + src16[494] + src16[495] + src16[496] + src16[497] + src16[498] + src16[499] + src16[500] + src16[501] + src16[502] + src16[503] + src16[504] + src16[505] + src16[506] + src16[507] + src16[508] + src16[509] + src16[510] + src16[511])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485] + src17[486] + src17[487] + src17[488] + src17[489] + src17[490] + src17[491] + src17[492] + src17[493] + src17[494] + src17[495] + src17[496] + src17[497] + src17[498] + src17[499] + src17[500] + src17[501] + src17[502] + src17[503] + src17[504] + src17[505] + src17[506] + src17[507] + src17[508] + src17[509] + src17[510] + src17[511])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485] + src18[486] + src18[487] + src18[488] + src18[489] + src18[490] + src18[491] + src18[492] + src18[493] + src18[494] + src18[495] + src18[496] + src18[497] + src18[498] + src18[499] + src18[500] + src18[501] + src18[502] + src18[503] + src18[504] + src18[505] + src18[506] + src18[507] + src18[508] + src18[509] + src18[510] + src18[511])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485] + src19[486] + src19[487] + src19[488] + src19[489] + src19[490] + src19[491] + src19[492] + src19[493] + src19[494] + src19[495] + src19[496] + src19[497] + src19[498] + src19[499] + src19[500] + src19[501] + src19[502] + src19[503] + src19[504] + src19[505] + src19[506] + src19[507] + src19[508] + src19[509] + src19[510] + src19[511])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485] + src20[486] + src20[487] + src20[488] + src20[489] + src20[490] + src20[491] + src20[492] + src20[493] + src20[494] + src20[495] + src20[496] + src20[497] + src20[498] + src20[499] + src20[500] + src20[501] + src20[502] + src20[503] + src20[504] + src20[505] + src20[506] + src20[507] + src20[508] + src20[509] + src20[510] + src20[511])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485] + src21[486] + src21[487] + src21[488] + src21[489] + src21[490] + src21[491] + src21[492] + src21[493] + src21[494] + src21[495] + src21[496] + src21[497] + src21[498] + src21[499] + src21[500] + src21[501] + src21[502] + src21[503] + src21[504] + src21[505] + src21[506] + src21[507] + src21[508] + src21[509] + src21[510] + src21[511])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485] + src22[486] + src22[487] + src22[488] + src22[489] + src22[490] + src22[491] + src22[492] + src22[493] + src22[494] + src22[495] + src22[496] + src22[497] + src22[498] + src22[499] + src22[500] + src22[501] + src22[502] + src22[503] + src22[504] + src22[505] + src22[506] + src22[507] + src22[508] + src22[509] + src22[510] + src22[511])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485] + src23[486] + src23[487] + src23[488] + src23[489] + src23[490] + src23[491] + src23[492] + src23[493] + src23[494] + src23[495] + src23[496] + src23[497] + src23[498] + src23[499] + src23[500] + src23[501] + src23[502] + src23[503] + src23[504] + src23[505] + src23[506] + src23[507] + src23[508] + src23[509] + src23[510] + src23[511])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485] + src24[486] + src24[487] + src24[488] + src24[489] + src24[490] + src24[491] + src24[492] + src24[493] + src24[494] + src24[495] + src24[496] + src24[497] + src24[498] + src24[499] + src24[500] + src24[501] + src24[502] + src24[503] + src24[504] + src24[505] + src24[506] + src24[507] + src24[508] + src24[509] + src24[510] + src24[511])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485] + src25[486] + src25[487] + src25[488] + src25[489] + src25[490] + src25[491] + src25[492] + src25[493] + src25[494] + src25[495] + src25[496] + src25[497] + src25[498] + src25[499] + src25[500] + src25[501] + src25[502] + src25[503] + src25[504] + src25[505] + src25[506] + src25[507] + src25[508] + src25[509] + src25[510] + src25[511])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485] + src26[486] + src26[487] + src26[488] + src26[489] + src26[490] + src26[491] + src26[492] + src26[493] + src26[494] + src26[495] + src26[496] + src26[497] + src26[498] + src26[499] + src26[500] + src26[501] + src26[502] + src26[503] + src26[504] + src26[505] + src26[506] + src26[507] + src26[508] + src26[509] + src26[510] + src26[511])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485] + src27[486] + src27[487] + src27[488] + src27[489] + src27[490] + src27[491] + src27[492] + src27[493] + src27[494] + src27[495] + src27[496] + src27[497] + src27[498] + src27[499] + src27[500] + src27[501] + src27[502] + src27[503] + src27[504] + src27[505] + src27[506] + src27[507] + src27[508] + src27[509] + src27[510] + src27[511])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485] + src28[486] + src28[487] + src28[488] + src28[489] + src28[490] + src28[491] + src28[492] + src28[493] + src28[494] + src28[495] + src28[496] + src28[497] + src28[498] + src28[499] + src28[500] + src28[501] + src28[502] + src28[503] + src28[504] + src28[505] + src28[506] + src28[507] + src28[508] + src28[509] + src28[510] + src28[511])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485] + src29[486] + src29[487] + src29[488] + src29[489] + src29[490] + src29[491] + src29[492] + src29[493] + src29[494] + src29[495] + src29[496] + src29[497] + src29[498] + src29[499] + src29[500] + src29[501] + src29[502] + src29[503] + src29[504] + src29[505] + src29[506] + src29[507] + src29[508] + src29[509] + src29[510] + src29[511])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485] + src30[486] + src30[487] + src30[488] + src30[489] + src30[490] + src30[491] + src30[492] + src30[493] + src30[494] + src30[495] + src30[496] + src30[497] + src30[498] + src30[499] + src30[500] + src30[501] + src30[502] + src30[503] + src30[504] + src30[505] + src30[506] + src30[507] + src30[508] + src30[509] + src30[510] + src30[511])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485] + src31[486] + src31[487] + src31[488] + src31[489] + src31[490] + src31[491] + src31[492] + src31[493] + src31[494] + src31[495] + src31[496] + src31[497] + src31[498] + src31[499] + src31[500] + src31[501] + src31[502] + src31[503] + src31[504] + src31[505] + src31[506] + src31[507] + src31[508] + src31[509] + src31[510] + src31[511])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb70cc42ba8241309c5a60d345b3b1f61dae9ab1778b736edda211c12f2e8d07398ccc34c047dc2febffc44fe08f3c0dc97a821d196ee044b4ca333ba0120580b29b65ac26266dac2cae6546ad61aad2d32d529b68553ed9e41904d784fee44d2eecf85cf020c359fd811e4c64ff30d52649038365bead8aeb3f9ad47f11069cd3439460c660ee2beef67091def41e5d8dcaa2f119d3ed9e5a0fc4d7f82d3637bacd12d70afe17183ec8780fffc9f887c19943ee3ec83959ceadaa15ccc61f50f16638370fb586c90934ac098924492b095d201acb311634a80e0e2faebee596c8dd58d527e56befba7837514feb741791fb76c1a9aff7e6c46635aa7b76b85a88a71b7daadb3e1a74387140fdfc92db8416874853d8927b4ef5990c62d1ea6044ad30edc697c437e2517d2dfdbc8f740b50fa005155ecafe566dce829c9c97bba54842ae095570adfd4098173c15644a38ba2ab800df38ce2eede4f727e9ecc4a0cf400c95df3d4ed479b7f5fed340a1ce7f46d20f341c49f4c2ee9cfa0cc21bc0bbf0b6a29012c9b06205d75f0cbf96b42b45d292f689ad578194c16299b865985ea8ba890267dae33aa2817806b57a46a091b5dd7224203c094b6de550614d92695243c9a62fad1fa372dd647c05b82d84c5bd45d4d42218bac5ad1cfcdabaeb4192dfbd9d7d514b55a4b91131bd95aabc7f48cd6b6b82fe2e1e557f759069e608d79f9dc43cece13a95b3cec778a0b0112c74760718a1bc579a3bcd1c41def443aae316319a1e4ccae769d2236920d8209eb0327c60e5cd25c7234cca9b5b11cb7a1147814765231da1e621fb48342cb83aab38cd636fb079cc77ffd5788ecd8651b33a6cdc6e61cb5d8c2fdfdb7fdd0620130e36327b5bc215100f0f37e52ed2b9bdf3a42667c6ebe0cf7bd859568afc2baabddd8119ab47c0436e5db5a1c5f81b58e90bc7409a2fc54db7aa6c1861567ae5fe9a55d8b01fcb70016bc4560f0d67e9fe81d1434bc49b3f4e7d6b218b2d0a33294b90a0c6c8fb6f5f89af205e599b51cd280d735d12a8b136097b6afa7a5fb1b1e06d8711da305447dbe0c8bf5b596c69828475142ce596d488c3774dddf0d4a57194331bbf1ff9ffeda5b1f77b5c48d29096ef65de7a7fbddb5867b1c6dc73f818b2ec304314400c00ec081fc266b7e5fe2c5736afcc9ec95e0f22990fc7c574d67266649c943c697b14342f89b37fa0ba180f0941d01b770229d020a922d15170900a219ffeb1575653f954ec6816012551ba0ab4edd381939a6c8b455e23e670c9afc3c8bcf6c451405f79cd23f182fdee37a251958bba0bd3560e7c3e357ef7eb63cbfc9a0431b748c000d09a469d87e8511a2c8b7341a07c2869a729aed305c7e58bc27d0e8fc6feb6fa1f9a8a027c869d91f600f60cca74a678043cd64ed341fa95731f28bf6ca701dd76c697063c71255ba4f626af93f1bb7259e7cdb4769b7e15b56d104005cd0f2b27b5d81dbedcb5aff2bbb6d3b0e216b8a656a07a184ddcf5a63acfc244f835fb6de5cf699446116fe9ec14d18e85a2f07694f851d0c26aa6bbefb3c90ec6d11372460a69e68a07a24e0d9ee341e672787840325e73dd2715a01e01822217690d221f19f3d76751e0e82388cc4aacd001f55b1163c8c5397cd707adfaa46e6ac608fb6c498c85cff4e55a9aebbc134d90875e2f4ba5fbcc95969c7694db7570bb080c592029647cb8b124c3575d476fe32738f044f9103a7d09c580128de0a70e0aed76cb6d0a12c884da403368a58eb299d23f49e40bc38cadef388235a9bcdcdce44fd0548ffa8b9ce3e667823262b2e0e12cdc3f258b5e625cba46f7efe246b5d2f377a3b0ce20df9edcf775754b3e5ab1b443a69e4ac77c1022fa207ad98b4ed758c12d62b5a00b972d5879c2c35ab81b968701c4eaa42854a242c2fa3dc1c853cc728563cc1f4e1a20844fd297115ec598469795644d1676db1d0543432dbfc42640effe940b3b755dd33b7ec8e216a1b9fe6daa995852acf9150395cc29938c893f1de7c214754219d274576ac35f69638ec34cbb9eba070401a76fac080fc8192542d50583f6f5c58104408546fe951c8095d5a8fa454981dba010993fe3ea101420ab23317539999b3b07a281278aa42543863c974ecc229d6f3e2928401f56903b2c404bb0c3696b83f299acc7b464f60900ec6da3059b774bf994c8cac21c4073d9d4ac377f2c6f53f43297fa0c25db8ca64bf9c739c583be46b6d12134c89a9bf607ac3779852ea6b697e5de7a71605f42bd2996c07c6c40ace9b7a5afe123f119180f1aedbf47ac35e19a87b7e9dd4bc369c9e091d47816a4b3b898ab22fc3d8d92b5f879bd70b4ae7310b30926758e128da5fa0a9cf1dcb77ef5ae48e8c9983de479a4e309cb0ea1f15dc3d14ffccf25995a16895938cb1bb37ddd560018db548c20f4fa1b0062791805144816a1c5a2426897aec18b3993d27d101a3336a240b2c80e7cf44005aa1214a1089a9c6946a45e3e17d231448d8cf2de9736461da7c4e69ae4bc4867cae6aafca7d05cf3aa790aed128f0e3e85f4c4b9be5ec705d977c8491bbe619d6f461c88ace1b068e515ea9aa6c3d4350f4dae974caaa2e4a04fd10ba430b73cb228611d2d8628df5668106cc3d4a2fdf256334c3e528bcb0a99ce036136278e3de212ae158c85a936153c37f39b0a19dfec52527b43aa86f950b1497af5efd83739dd2c1d68c8c92841059e6b9da66a9e7e0afde1dcec2b2ddfdca2cde169a33ee1452835e58159ecff0912e6659243186f2dbebf7f9a99241ad8afb99cd8abd37e322e7bf48d505d77b3cb6df843b049576d89cafa635b55c88768fb466c7b9dab9d09165e2d1bb925db970750fe968231;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfa1bc1916c673677a2ccf618530ffedce8a4f084a3fcedd9e1636025be6e67a2ad0efef91831ee73403550a3146b8fc82267ef7832d7a7df2622ba04a71f07cbe4569307ea7a935af2593c5e2a7c32c220b7684a505b409222ad0e10cc6ff01f32f51d257176252c0a2d238b04e56d1b81d7081131dbcbf8b3747e4ac601a4a86965a0ae0983742f568d07450297dba69a36a5483248d7b31260fe33acfee8a7f125cc8a999e1e59092dd13b4a5f78eeb478388d5cb7974ce1d7d7b1c4c89f0705e63e0113f8104008005fbc20f7eea07f82b86a9d65872d9ee80f4f27b5cdd5ef55052489d23c7cdcb7ff59fd87dbb7a4efb5e9bdcc451238bacf6d24c77fbb3ec8c9b655067989e404e907daa8b605ea49f6d800c8cda0075dce6ee426a883de0695c614c755244f8a13dc1c2e94b7aef168b1a108d2ed4bbe15f4fbd33ce6765ad8984609accfea6ade14664fb8033b5700aeb4b64fc123ea5a5ecb5f1b74abe4741b740a03ef77f1edc9207cdcd7b83cfdaf7e47e8af54b2d6957a9e78870fb81dc6a9c971437c56c72498224e24672f07c9aafcbc974d733a89718e6cf38c5d8bae9f9ed9886e28a849c71487eb759c081ecf4d2c205d1e1f6ee3f7c7043a7c1489a4ce7d8b70f7514e2a2ae4e1a70535acdd9e3c8597796c58c14f768134b96317e775fab7b44ca564f8b2ebe323e53f491b64334e647b1d774a9fc6406571bcbb6359a676a292c9ba00b206cdda8720f77bd2634b23a8faea67ba83120a8f3343b20d704c8b202514cac7a8b19258aea1e32acae3ab86ac0b45ca18f3e63f4138c0e5ea4a9114aea943431f9298c5114868d5a4de4b1e1597256301634cd994c114d94ffcd5657720821e499d69630a1bcc71635a38394faea048a1890ab477d96c8c040f15f641dd6dc1edcdac44d1e6052384907d566f6a39d55072883be58cf1c17fb926f421f8894ea3fd5d3ef30624139f27f90d4ba1740d947b005f80f9de47cfee24b6901119c371e52add2df143a920ae1b8c8fc508bd761c85dc76da93b137c05f7d008cfee9e2bd9114eff54e29cefb40f4254bb5e209aaaa7b3f91357325fca57e74c2e411ec7142389e88953e34f5ce8aa72a3645bee6d45d31c95ab93fd8c818f74d0ec7386f3c3c7767b7a0bcf166740e2b18ac8f846fea81917259cbfddbf0211cd8e43fdcf6a116f26859642621000532d6d040e1c04ac2d579792bd2e0f374a830856eba83e1b1d3b64266b886dde191591e5b35e2eec6c910b3430ac10127b1139879ca4112f628d92e7c0807d6686731cca7ec55ad0a4b185b930861f4fe5635c2c3494341a1b2a862cb11becfef4f0c1d1338977abd71cae6f8b28e68d568321d880b3abaca09fc93c95b8a73ceab8a4677d168a364517077f226adeca04f7ff6f5c348d4fa091e974abce5a612bf351ab11d2d247e3e30b19296c02892c621775df5045d5c8a5902e32f2b9c2bcca9a0c67f4499b0a0cc9cae555d9eadc75d348ee3d70e584a22c5f44f1686806b2435bcf7eceb499aa771c0e5e15ee4fe48eb6665c39c934677f0a6bae6b156d74501c8be89d7402925130ed4a40b644b725e386b641fcbe561af82ff2f567a377758d572ebe118a13cc95d3a4dbd35377ef09957fb94036939970c77f6d8c36bce629f92a86fb8620446b8f9552b1194d9be0d4ae587288a09a9b8bd58037bfae6848b66cef170af8dbbf8c5643fd0765eb4b00c9ed9fdabc9b8e6500427431aafd3def961c55fb4d54a3209748db9b3d52fc93f3b162adb0e7a3f2aa10c2b6c232a224a491dbb1495960abcc91e3ddc551d3023beb432815ead930e70c8f6cd98821dcbe219cfb820d53899f4d9004582287d8a1afb65409a7e086ee803c8d895a16b4cf5f9a8c8153710650c684a69afda5dce39446a256b58d913f67ed664f90b03811e85af7bb05fbb576904af2fa3a63409d2f6ccaf3616c345fa2c08509c2cb70993282cb291f1e9cff280ccb155c89ec24e2b2bec2689bf7649ae246d52b386a9487735352401fdd14b49a681adf299ac4d8e7230a2f29892d62e389f71c3787c552ab8f7667009d6879939c1efbe4bdd61eaacfa185122335da3441c26478308c5fb3affc064017be9c745d07c9c07857d5c5f5c23ed7cd758c16ada84782af65dd5a8f80472e67a3e1bbdf1c3cb9cd69a7b04f9c46a3e4b777d4737a20963cd4b637dd871017c7a07b4223a81eb92e47b6a1c40aaeaaa1161342c29425d70194c8471ec598269e6762cb19d3367574f378537609119710d3545127f0dc518d39845d0713ef85bc3f4df8b01ff8f57939d086c9216f033e0da0938d70800a2326cd009c08fc0faa8ba8c6e23170e9d4c4a79e92f2341409cb1cc877402c44d988e0da4d71f6f043a1de5c7a3b11af7477ee79742950bc529e2f34c92b53a83b86f0882326ca6439462a1566d40e2de6de7e30ee8bc4ebf71579eb400d6cf2a82184edce7c2fb980aa9fe46aae8602fb14f3120db613efa2884af7105f0a90c33938e58371af4bbe8a98064d48a8c5cc3b9586d4a35ee48bb09b0adda1fde25315719688368660896943ba192c3d224173936dcf6ce8ce2d4a4b535937ca621d2301d1214cc292c7c33833aa2c1787502b5be2bb773086a58afbff86da78118a62186a828fe0f956a49dfc17eeff7dadd65fbf1322d59dc47de6c09cc8f0bd4d5fefbc2b5ad9e9012c37fbf8000d2f6df3091bb4f2fe9870ba994f8f24effdb8facd33e04529e7825a88652ea2b0894b6f3a640d4f755e7a1f9f3a7ce3eb6bc9bb8303cd303d908bd998d61bf9ddccfc1c7dc47d51a6d20a719bd501cbf93700095f6cfff84da51d812c0276909bf44cd1f32fcda83dda85bae1d9f605132663;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha4482752058159f4c23cbe4902d2a89e3c913deabb5dee1f7e81d0ac919fcc0946a5aa353e238e5bab7c65d278b4365e40e1d08c0e6e714055fd6ed1638d0a231f5fbb1c286aa638c9b3a6867c29509fe97c02544dab495492d3b98c6589e8be3d46ee7beb453fb12f252e7a8209c93f6182a6a52ffd2be8ec3765440a762f35e13a21cb5e6bbf3db48e97da18f014fb3a549073d2afbe0ef704371f75b6c2050f364893fbad918e0dd53eaa3882d3dbce77f07dd77f3fa119f637f99251749512f5ef1f7635ee8ff7799efbcc530fa3404af377fee1bac8ceac634def6a495df17a5da430435d7d0b1c32ab73de1905f07a5946a05fbe1ab048f7958e9faf2a9470be9dd75fe3b258b261b46958199340688c77fa809866beb2ea2f8909068db52c4f1ee296e8c4998e1a3d656613b6c14a3a8f48020c9f3a416e49bb1f79f42f9c174ec06579592e14a890d57eadd7151e2c77825f6cb4b02863186690575c3c4fc25069a6305df27564718d1f60adef3ead02336b8302446b2c5e8bb52d168d4c26995e8b79b387c7e1a974db65b0461a383900ecc3052e57e911444bd12423e45b98fa6874aacde0e1208ddc2cf4a4fd1f8a7ad922380a76e6746cbb2d29b2f05e90455748c475aa4b6943482bdca4da0a874c35b0171254287de63cfeb3ab0711ffbb080dae49e74d064213de5918030d7fb653b6008a7e57e0c26eceae8e35cfa8667ddede6900c93ed08c5668586c7499cc0618f3b851a449d9d2277c30878fb42f1bddccba2d3c59c5a8c4c9701aa0faea56eab73c83aa096e1c7aa0737f01bd2a8e0158becbb23dd51266a441c14b6691e63d838f968484f8a99e1b32527f0a05c146ad2d27f25de330ae6d916404e53276ac17ea9a5d58c04f44021b9ceea0494d6a960fb4f13d875cd1e4ec1dee3c5b381663160da34a86c16220336beb9952178d5619cf3f6b9ac480f4dfb09c417168ed0470a3d18a13a23cd27590642d0b65d5648c80ff92bbe83b6fecfd354602073260b7ecbe4755289534433a2c25eae2d6dfa62a31f402ab3e7ccdc701ae16f13767ed9fbfb2edc8eefaa6df1ef23989d182c52acb3851e389845e90c4ef0b37d26314696e6b4da5efb8e4087206966cccce1a7f99c0af2a962bf4afa2991b36fba3a14237326bc4c012d03fce93da2fb12e4c100e594980491b5a012661c299d647034ed98a85c65c5fee8787665f87eb180c0bb160a1ccfd625cd38c02777261dff3a68b582d8797d45efe3957d0361db8c7c99e03bae0f0391c6ba1b1c67f1fc9e594812a177e5bf32c426c62cdd0a71b263e243eac8274f0da9f314b56865e5478c54e9010857a5fb5b34150f124149aa74da9b6f49f544fe147355457571990e9f403d468e34832abf2383c3e911c2713aee9530cfbfb84e32e61f57b99d613f192c83fb8d960c4258175a7c870778d901ac1f6293f387d7bc40153916523a54a93a2391f22d5b07d1f77d15b8d4c4655930e7ba249b2b64e64aa7d0fcec9d3f23d00226715c1f65d7bea28173477cbf6b9b02d7145f8379b3b89c03176be5af5730f92b137738dda4a0bdedabd125e88d675dcdbd8844d43af87761cf9f16e9a5d3c7be2e4cfa34dfc30b6951a02e3f760ac2d6b50643309a0bf8616c999ad91d14bb2f9269b646ccd0d4008d1398d27bd27a23523e69dcaaca6e2a74b66f862a21717e81ca52071fcf541a2282d87fea179b08554ff9778ceb45ca97ec4ab522537c4323e4e5a6d2aa802e5ab880881ddeac2a211eb6313517abbf76b6519190f9b2214c6859fd7b701e278d66a7b049c60142eb3d01bb51dc0d2b0fc0c7dafb9171a8800cc8096592e2e7dd034a391d4a63bf114a3c66a5e7704925e3f104cb38b03d8cf5beb9ecadd21f1ad848b07e8da6d3ab48200cdc28f4a06f9a6c787098e75508556efc662f2a24e1da5dcdceb6e1d8192691fc29a74d69d867467497ab72275496cd53e0243ec52b4ee905ca1fe15743f79a449e0963136f6afcf12717a87b2ee744ee5332bd3ae6c716353fa24ccf73427f933c17e1903895203304e8948ee3636a17cc6bbcb21bd0cc7c64339d67b78f2eb03b844fe376fdc3fd577ae887669069ae9ac14f5273fcf4b842cd711eee766e70fb19e5834b0f67d580b3188fb555c757d73719b5cb3e4f73120127e96aa278a35a9bbc00d39ec8be11482b62455504bc3cc06bc56f885a310cba37821b16d9431c505e47982a92a88f03205388dc2e4f3991b5fb06595e56eaac84d2dbd9a29b68712d95d4cefb3bbb9eea243a40fabddae4374a21660d5f07beb79a8125310f929e14df017e061a8e440a05cdf5e8e22677a52d8e4dbe3c20cf59d53723736f93b4c711f5482b6ca5a0337aa6608594e89a3f89c95d2c40f878a18a8a1737c0289e316056cbb3a5ab5ce3605be04f0c9d13270c398b0e45e7d5a59e6de6efb143936b69645c4c646863bad7755d9089cdbf0351dc2d90987c1227b4348fe82fca970c54bf0d0ae18922a300eafc3ff196893f8628e4dcd2f8d7fe170388d79d66b3ede6f0fc116ac0adce38f521dbd32799bb94615a729c19c7a1c51bb5aca67927c2c3af10d0b4e35fbe71d8a7ea50378144c6e7f7bf77414f20d5954bdd65477194e7715ce23faf4c978c85c939b9abf60776ec9cb1187738a69d092d61d8f112b9e46394b8fe35f61c2c347570db1f2cf1691db9e672d9b45dce4a625c68363a5207e7da3c2208ff593923d4a25b4f0bb8132a176d8f735b75de4baf5aaad8d5dd29320db8bda0203e6fc4cd78aff6a75bfa07829fab5f2d66ed8c6bf20f4576385fa736ee3eda145b5beba20f3ef32e62a31dc37638c06f6b282ad5df9b2ba610581ae9fb36c9f4714a38af268;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h881e013db755fabbd8d568ee2e779803408f4a1b0547cc2485a8140e5290e644a382591f88463dc720fbd17465d4ad64dbe5fb488cc8713a356491ff4c36700f2b886badd8dbb1fe6663f3447c1132eb1e102051c3f777557b3a3969664d512cd24037d3b82025edd2b4b2532dbf0a5af9c859b03f69c0690b4c6da0c8ad4cfb039cdf66ff60bdcee67858740b2b0d421e2b470090954366e5afe9bc1b90babd667d7a5e8087550560ceff77d5744ac61c60b363a35bc8139cd48532676a97da49937630c4d58ca61b418339db86fa40b9b98a1f514696b77a93915d1b5ba10cd6db5a05a03cc43cf0da222cf5dfbfddedc1b04d4d0bdbba4514525a5b2703fda57413731a853c4a66e2241149cfcccd3d165d76ecd71fddda4cfabd5acf9db1808f934766d0add6fd6452a6daad9e9957085f6d94552a187961e0b764ab0529c34a6ae2844491e24d3661061147331d966bae7be2c6fe6cb8352afcbe6f496d130a9ad474b631f0222eb80ba162aced3c2f78b3bc957be1a44bdf83f2d504665c608a0d31767118b34f841ada1fd7ded9f5679d4704bc2c9a8a590e85ae82faf9317fa2aad978696ddc32b4e88fcd8ae3cbaaa179e275d60b3f4b49a04222ac7728fc15fae9c28ed5ce5dfb8fe71a72372efa7d75e361a4a718d0d56cc75e915462c9edc3ecd497ef8b834dc7174e1e03f3401a69a20fe4179891f67ecb00e5e47d97fd2697591db13073d5ef3debda045d6d3e9c30dd44d1fe3ddd338126330e717c4f9d41a3dfaf24cd8ff5e5ad35d02aead62387b2e3b8afc41bdcccce0c3c21f48ed996bc1adc93c1c8bcf9ef40ab26e56b13e75b542a6464be2c5bf072bf76097afdc296404803cb72c3d4f37c6a6793a6cc007479ae5dd3a64de69eeda04bd08178bc057bab43bc5ca3351d2ebe1da300c4d4a2f023f736def9ed677ee178f4bd19981b76f88278e1cfb274a4f052e8940914564b411de802c9d76eca3ef69b69eb4bf29571bc8a822036dbf8b985db2ba84a7c3eca7a9237b333b4fd034b8e014b7ec0f55b1026c48ac6995756eb936bab680c9c37575266582352efc5aafb97377d8ad6a8750a45194a5a83f11e268bdb65e54e1d541fbd406841cd99db1137ee5f549f07c41c7a911861bda4124426f3a50c20a7ea2639bb6d500ce3f436a964f45c7035fbfcd6314559f9ad1850955afaa0a17fc2538e330625c97e8d7cd5ee997b50a06c71c4a285b1179ddba7f8d6d5baaea2a430edc3bdf666b542aa116da3cd28695e7663e122a40ff34e84377223a70cbc6a540cd40db1b35ca88658c3f68d481ee66054170d8f01096533112420d5141951faf3ea4ef01419c1731f11ba60b7081f1c860e7225ac4fdc132cbb5a1b586007a60e91ed3791436683dd0c64357ff0b81de8aec00dd4ddd6a15db9722c28afcac142c5353e2fb3e5d15ba7de25fa06e1cab0c8fa82224bb01ce0250dbe98df1db43b618dd7eee82bd9f0601020d8460a08ef3899935e48704e29c4028a0b523648f1c8d3ea8cc6c39265585b894f7281e265e1acc709ab76090640ecd0312b136b47c1f80c2edf84e1de466ecd7623e6a635cbdd9e6055703ca70b879f9a1e8dc8695aa8451bd5589fccaa50a0543e79e2ccfae78ac6a705d6fe6a286bc700f7ad54fc102feeed91854f8db381770a6c08a9bf6cb861c321d915f08c822056a02720324582c8c6ff9459e1f89f77142041ef2808871847a8abdd6fc08359e689991edf9708f49e3f87e5d682fd7d81a2520080a7a28e28e5198559a6172274ec4d2df0782480e615beb8aec27e78302ac6a77103d664dcce3fc790df54b0c2895b69d3e21ef6198afaf223a2f774e4f2719d2da7872205e124b0b2cb1f9bbe45ef4d272e5a29ca2057ee52b1dd31eea6fa9df177ca1ac43adb69c594a3d061ccad2b73c460ff3f891c3e5a72e1535f37d0c6e1db8964cfc0f18a67e91b25bc8e230f10d5cb0216454bf5f8f1859347a8a34e33b8d755c71d16898de912b43b560b200ec296ebed72f8e9eb5101fdbe2e677353a93fad907fdc5cb06df33d18cd5f7e7673d99c07a3be7e86707ffa1080d16cab934ac6a40bedcd33bf80e9d06a47a57b300adfcab4f899896bfe6508dc07ad03b2fb45e9efe6773e63472112beb67d2471686cce0fb0e813e30c720eb3e328bce195f49d50fcd924093cb5b7fe209f4c9ccce84190bd5bba1653e8faaf1f6ddc3053082ba1c818e124312ef1c8f502761e6ffa1723d1121647735afb00581e827cd5740cd22137cff531fdd612bce312a731100c9173bbfaf1b962d0bf92988057bdec27c33545b022abf1e080525ac226103e6cf14899a4a6d9b7ef5490277e8b4a092108a9183ff416ba11d0ee2add5a8a96fd1a66798a5f83c17ccfd1d76e47197f3ef5549f94f13113012dc58176e398808cfcabc5949e795a9d22e53e85c999d62c4e2789ae66b4bf7160b71e6e8de96054e3d675b7cc074ec2afcc4bbc6eef17279b1e50f3e159b23b0ad75fb7cf2893e28a6df12b7d60922e79811497e8476c8efde25a3de51ac4cfee4bcc83edb01446ed3060806d0990e445125d1ef4d99d9d42df4be2bca7168ce8935cfa4c1fc19c27a368e280fa3f975c87533446a28929f842edf71ac9383807786f9da3be6d89b5ad76d9cffa1861ed9361b88ff3a38dac243793c489b8da47d4c0167052643e70d8bbdd85a9ac4ac1ace2d336ff0209d194a63856abe0f283f3a1b152b7fb2d013288cadd974385bb7f11aa1751d5aa26dfd52fab20489218aef5d01a17bedeae778fe2f9c718a3a5f9b96ba19f31fed139bdddc36f166e2949c50a36f6840f39cad41400421f1ee0480303df4238bd130a86d651b1bfb394ed3cd4624a8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7198e5d8dbdf45d0e99cfde32cad5ba6e743c127c6599860d2f059e8e5e03cc5b6dd12363029ea16ab395b672df43ef9d5fed4c91fb2c3b70adf7878813f05d298203d3bd938639e5564c681c90874d0a3cb36b67fc6f4f0115f96e546c601b614bb0f34e5e252dac23680ab04b8f43b2c3d028fef548695c95a77619144e1f9bb00b840bb2b5f1582d68598bd56a1a1ef1c5c33bbc7b0b241661f221deb70fa779237979a4c8817ee4023845f5bad5b5dd9aec4c2e9e049e5d17418f4977048ad8f523cb93fba785929ec3fbf9b34f12bee5dcf5b37fabf2d54e7ef09a8588191757455f7cfa94d63786f807297cf63bb64f1267dbafc8d8e01319eee68fb24f4da577ee1a62b276dff04a0e77671ebbc9dff85e1acf5325406cae1bcdc8f95edb23432b2de37110e855574034add2ed91d8d7b1e01e53ad2008ae29f7b13e618725a7e3abf8454e1094361fd4bc2c490266b8563467718f744ef66b90e8f959a9b759b31005c60f7df65db401b271da5ddc6a6ce55608e6a93f15859d96758c4e1259bbb050109a5412944dc7158380d3ee622149db0a6e021a96c8131a405a6681c0e8dd0c6e1a9ffac3cf0b87b9540c3da32dbbf973bd47a1665f39c8551db04fde21c127005e6132d12876cec51486e98451bedb473a30942de5933105edd4f14ad27ecbe1a40ca51f12bc2396059715f0befa30f2bf29298b0a556397688f36b3e95c4a67c7c6c6117f55c0620d3a075d56ef169dccb7578825b7e4729ba0e789c1ad302e5f8db3a9eedef79455d47bf3d16c3ca35e718236a41a96e0941d80d5c0b905a128b28016a1504fe315904d26103e0e9c8bbe397deaf15eeda7f0cbcc394fc7844805abd229e9c6682a01492e6b2eb6af3799934bbe6d8a1e6198128e77477800ea98edae692cf4e9ccdd18c45316d25b315c558e68d3283396a26b82d55ddf4c895297bd3f35fd4f0f68aba6ff60ddd8ca85bf56c8253aa1ca01d432b7db6403eb88fb29f934cdb7c55daf6ff305e48ba6f2597e81f125c91ea993951496a2edc4f148430099307093cb28a48d5266bc261cc0746609782897626937bbbaaa4fcba57b62401ed1226855634cc1a18a014227582dccabdec5d14eecfa9e2fe0f5018c46e6e3ed3f9309f6eaae840d51e2d31edae84fd2652b58099f7631e6237161c5ad883ac85df68ab94b341bad29a43ff85c1f6b54a7f88db7a773d7b80d2c11724a21334c08c6b293ec0310aaad071dca22e047a23bb8bcf71e9fe7fe07fea771409d24dab86911bbb2a9098b460a543ada66fc5e8f0b3b38c06e8f984e164a2bbaf22a1bcbac09bb846fdd0db8fa09559114dfbace5001409b7c1e4028b21f488e69fffb0fabb2a5ec62eeed3fd99b8906e7f4c028caebcc8a647e98cf7cb86316dc8f93bbd368185a9ece5f54efb025426fa390d7300b008316bb11663995f498fd3c87514fa048317bf66edf364c8bc4882b5efa6e2a6afb2c166a517f5a11dd8c5e8c1e7c43f8e442cff3cb14ba31c13de350e724dc7af9192a6d694a345f044800a19da9f7a3bc27b9638b8236265e489eea1ae54b1557b64cec599594d4bad4d1e223011a8bdb3bf79376601df46c67e62efc4af71a9eeaef8f673acf03829913f7198e343dac54ecbc908d9fbd393ad63421d7c49ff7c5452282533ea03dd7ae74d893539285d3e351cc05270b3103b6fde72fcef5ddc79a5378376485fee410408eceb7ff88609fddf8af3b1b5a7579c8895816dfec5023906df862e093ab895a73feadbc7a02aabd112dfbe361e0774a48e9a50a2ca0c9333639e245fa1cce4608349be64ad19967eba4842633096aa2ae6f9ab5417cc93658a095547f6e9ff095bbbffb38667617ffddfa3d4638cfa405aa1be5adfe7166758dac32d8b95f2e9b926e97561018c0082517bd95bc7c77a23d86770b2d7695c45b736870b5ef4e0460c84de24eaf5fbeab4ffa40ddfea879de95036575037d4f7180df97c5fa883bdc2b42aff5b76bc90bc955e59fda6882bdeb73782e79858172570a2091bb269701af5a1a30c4f9e03140e7959b25429b7e6164b7ababfeeae02d219484d5b0a6dcc03f46607f9a65e0810765ccefbcc527e9d350d829a60324a333be3c73e2791bcbeb1143180fda4a61280471f5857dc06cfb740539d531da9e4c1edf0a19364a1df8be6eec65d6bc051ba2c960960b6faae1a703fd45a05aeda4dd799c627987efd4a001c76fa38f90f2a57cadafcb2fdd17da863975f38152a78170842bdef327f0697785ef2bf4e72ce89003f9a1fa50a52d27db7802e0bd2644cda749672e89add621ae803b56871b72c6a96f19f70bc093fcefd476bff8df8fbc688b4eea2eda76af2e096225884141eee384378553cffe4e812ae2597f430d51e4e4f7767bccf6ef3c9ec12037e3ad7833bf840fb49f842b310befd19375e6dfac32b3c0a3ed4954f8801b4ec5f1edb9e0523e3f4b0865439af603e6496b7079c2d2d48130770dfd3dd0b3843dc86a612bd584dee156e1fdb1d3608f0af2d3b1d2459841d06dfab927d2b95d31bcc194d90c02b22bea71958247d66f6b24f95e8faf7db207e5e4533219ed15c107063ca90f371f496d76851908a8cf20e7c1f615e73544af7c2ce7df8699ed74c90827ced79b79d9fb9bb129a0d936d1d002e114001715353b9f799dccc4e72817fde068b768c64a8b619b2d3e4ed81e027e341dd36265dfb37aea3116a248374faf1aca6ed52164599ba4cdcfb9cf4e29ad2c6adc00c7e3cab4e5bc01eb07c6b0910871441c17d1b679dca984d52f281232f77b41471b20b51b93f8614ead7d28d46fc2ce89a1d60de2b487de3aac5a0f4633f9145f1b25194f90f77d35c2e364c3475293f7898;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h17fd8a8d699dafa608592c16900f0538b981a1b7dedfe4732881ac9e3e4bc35301cf01942bc0921638eb8d7205e22ac1b40fcc1d630e91c060e97c8f30adc6c53c0f1e1b951e07874728796479e1dcabfb42b853a23004ae68ebcd823247cfb0a7988abf86bedab22c3ca57d3357b064d78e8ab822e550d8744780add9ea1410fa0956f3dbf643df6250ea0e70d2d13e18b0051840fcdf2f46a66097d571c2792f469c0a6d86d5cc6d3405918ace1c72248c80b7dc97f183f6220bbd4841475a3fce4019dee4ed9f15120348e19c0797b743ef5ba4670b6814a568107637825d328865790a86298f733f763a25cbc242bd63be5d0bded1ffae751d91078dbd05b54aa80acb16b003a8268a728f2813e9116e56540dc094972b30b01c6efe7e788925b91bda16ab6d029aa83ece463f127f2e531cabd0f490d2b08c210cc627eb3247cfd596bc306db0bb3d094e8896157994947948de0441af6475a7945e3840f9db5ea3330335a02b0ebed5b6209612c8741e558d309182faec3052abffda0b2b00fc2803ba0f168a95f7c37c17c3b7a2aa3672c6b7d3667b2be837a87adb89533892037874d7c5ad8248807c7f3ca76cef1b72448ee19974710f92cc5b0cc1b474b4c8ab885df46ba76fb81a6d5f7a04c357ae01fc39dc413eb8b3cd2fff2db0df1cfee3214d9bae4392d207e47b362904cd556b359474ced55dded99a125902009994a435a11e4b7226c5a0daf3da4f736142fac31e2bde3ee82c1610330ff093c1999e1bb7a4ebf3b695538d48393206df5ea3a9ffb63898607b0cdd553729c0e939ae3d49212020d4a8f70b8e6a787666909e09c06a368acd034173e977477fa401cfb746973866929a656c75f6412e1cefa2b2a1d3696cc2f0fedef92b070703b7e96e54f1eaf16f76dd5870f0a15dd5cc55294d6ce127e1f8c4cf3915f6efe2b94e66233c84d2abd36206039ac1c19c4a23664b813e6fa1a7de7cff5f9308a92db1397e4f5865d89afb217329308d2aeb57eedfd33124e65936480f2d76c73f784aae732102cd8a00d5c4385983fe0362f213c036909133315f55b8b551f3438119bf8a59f1b628bc5a60e3a68f56c4df4d131b8d2d93af2ab951e2c3fd0e10bf8f1c057471cad4c52e50f6ee6801c3a73b960b49b3255e4dcab3449418585630cf7c3a6efacf0ab2fccff41ed0537ca39c2677bcc1a2e67f908f6ce7bd75f78b1652bbbe47605ec1b69a77d99f392510389356aca1b346c713b9947a3b2be06d67300ffee059783c7f00882c7267641064da4f42bd0feeb9c23491a8878cffc76b863d2300f15a87eaf37007d8360c47da86240e47356ad73a479c18ed92acef12a277531c6129a79d874b5048918fa9d3cd7deafd7e599995cea5445e21b8ee87df5b89ef4bdd577405abf13e18b0914712086fb6eaf825d6eaa6f4c3960c46ae27e2e9d5f747ca89a7d5334cf9f2fc6140308b01de0ee9a9698c3b1d3cec243ad967e7470f334df16dcd81afa7db1ce74bde3a0238a24223588a05e235bb180b210c07bccf125b9b3d7bf2fdaca653c06cf3c4eaf0857fe8bb34f22fba14ca9d9241989628ac87baa063fe88874a979b56f52cbda2e77e0a035a8e45fadec7915db9e7860da8f5b1fb9592b624f45e76625f78527fc47a4d7af82bf4cb433852cdf05b991d2507145d37e24d7904934eb14d3127bdde2dffbef00ae7380bada55ec83bbf92bf5ebee247d50c66b816daf07ac66767431e63a9d288042d3bacbc6337ed40b01542340fe36558679c4bd198b537652ca1da904b1291018584d6075f366c3111c8258e4cfb0ebbcfbf81bb06c8ef3dc1e842ffc877d5bf491aa5aaba7c605889e373fa4e5c70285ce863ba6c35d567ab7087f98a8e1e73c440390eec89a67c5f053f2763fd8fc2246179e54cefb9408110c188db89659a862844fc5fba5631600c99696ea6954296c927bfb84c1962e22c3859d6b0cd75f74efdcf14ca63bc609e00275f46909851f86e2cefaa5891e5c2338dd7eb9a07ca015128a6a6e7971d2eb4e052f888f7df7503f75f0686b9040f2eebe167da1577f70ab23c7fb93d937ecb9c609b591817b8d1625a20b497b40dfa17b9ded8376e42915e80ad7032a55aea075c5c6e2f362bbafb4750ee7228ee192df366e41754adf1603efcbdd3e647ea9b0ab2b6a767a554d53d35376f8c659bbbd4cf564a04a4df0205bc65a1e4e7e2d504197360c81f198f6aed26c7c408f435804a68b96cd2842f0189f45da5fa3ffaec7991be1231eee82e634a4a8198fa1f4264ac3b69e554234fdee8759ee32ca679ef3dbe818afc344b4a9d904c4c2d59f9d20f59e628b543effad46b823770558dfc61402afaea28a895d2bc2da8ab252a6fb585ba284ce5ebd7271a625e62bfb2839209a47c341df99f2df41782044e9a835d8587b46b5aa58996f82d8c9302303ed3419ab04b4c1f6ff3c53c5c1461be51d5374b91667b9feaa63e6d5faf1439de32ae719dab0546f7746ca27c1ae4898c47fb9054ba30f55821122e8d76da49e854b95d5c5ebe4293483142fd10187d910144ad37cdd5b7b29baae346ae27598fbbc9741c6b6e6de44d156a964692977605bf0a0e869b5973900c6ca9a7b797c64e6da65092b61f42e2f69f7936a9492bda09d324fc1e59287b067aab8d140c8a24f743100a3f2aa57a204cce0d53a59f5faeefd9526cef8161e03afdccbaab91e8a8de6b37406d91afbdc8abed24d9a1f5ac06512014054232da81e6a7ed9031ca6cbc96d59e6a568b4944164475c32a4a40280bb9926bbb9dd80c82a99137b8981b2f0373785eb18df97ef8823b7e77586e7d5075fd9284b35c39711612f34b88462aaacc5d8e28dccc492079041b5687;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf72c73b98ede17a297fdfc0debff9e0184172a8eb4242813222a8088393ece3e31ad643dfdf340e73801c5065354a93dcea1930995f16ccbc99f51854773ac648b0f7e7b478766888d2705e49e8dea86e930a2efeafb4540b46eb2b94ff460acce664fa817ba7f66e64d1f6d2d82b472e1b3d020c93ad7ffc899b4a77f0dd4c00b2fa7e8fa932bab5232f1a5c0b3e132cd18003cb3448190a08dcaf443c734f8dc529e0ccb5c0bd4366bc13cb7b365b000bc9d4d07efaeab7f829b0921cd533f7592647e05879994bad6208e3dc083b1fcd1ecb87d0de1d7cfafe7141552b860b9215105ff5fc61bd7981fd086c401cdc39256a1bfe2c03ec359a8f473d8586bcde2f6b8851870b3d2aa8c49de90a8b61f3d244881678c0c21a8ec09072accce0e7ee900ad12d9c20c0aa359314a1fe8457dcd4819b919cb8cfcbe531c5aa863667107a3ff141505b1bfadf136a8fd510f83d529457723e0f7fb49bc8eba44c0bd00a3a196f89e3db17bfa3cb33e51495bd127ed47bf7e88259fe08aa9761df362fd38fb64fef71860dc312779356d112fd1fc635fbf12c12421d60f8987b8fc80c4623c547ac61a749f31186148f6f6aecf354298154fefe308102ffca08401e22b0a60b9fcb7b2d6168a2553f2e3faa44dc0c40bb7724ec3861c9374b410e12c93fa2a006f6907e67acc55b713042fa2fe54c64a26c2a8681aa6d051c8074872f98977bdba24e4a1712ec2c6326397b3c5e574ea2cae43510ea2cb0000ea16ed8129516ffe6a29105755e697b7713201144b944df683ada77e3e782f1024f97378294363254cf195c0a197238db4067fb1ea84be17a678b332d396703325b9b7667281bfded6e474b8cc78e0fde10b61ea2ec4b7d853b713eb3f26cb6a33a6ec7417f3109dd5a684ee5a4535e8f3ccbaffc7d74fa610b07c5c94797ed0f6a7e32d1a326b930d086e7c5d09bdeeb4f3ab18ff402a4328d6347426a753fe3a81995782c52819ceade976b6a1315f5545f8a8e352255a67d1fa3e12b35e0b85e82b92eb359b285412928ab489b88a89648a7627f36c68f0a7168833df6d22b4b926f6f97a18fb106a4ea8eb68b14bb1d22817b8af497e3261cab9b344aabccb4c24eb0c9d81e80dc92b0763be2abb31a8bbcb0b3b7504d7f2900d23ef187f4f49167f403f0099eb86876b6b010b37891d52893ca92ef3eab570644bbb2dc7f17bf33d05bb5774d43f19632fb9d253e1d4d63252a4e7578fd831f73f0a756de5240d2d2b90a9def7b978d29eae4e65f52c4f14edfb25c0c928006edaeefedf2f9d4328e160b5a62ba457aa818a46ad1083b9007b215e5181ffac1f8dcfea6a161ac578544eae286ee2997885b311b002685e088a7d579fef89cee11e545515b3aa7e8aa1e30a3a01e387ee136ef93cb02603d261f98a0462a86067679af46ffe6aef9244b8394fb4fd91e451d4076ca696c37a5b9867fafd33655385d41c02722a0dc6caadc305ef10975c5f638387e1e9fd90477b77097e0b22bca6ce1a45d5726c6a8b5c8ba68952dc63552b527e09106e65c52270988ea6ea0a7cdfb2c9255b23c8bc35645f77e5120ac96c91b32ef089fb56210c1d8630d2c9d095ce380978eb3fbc447fd75d4ab260c8e0c9722d828eb3f3709df255e1689bd93da755edd3295a8dfa5149861c2d67ab49f245724f0bcc29a3c956c663c46aa7ac825d3519c05161259b393a65ee954609b4b30890e6949cd59c6c8572460fffaa6efcd35e3da5df82e237aa838a0e04806a2055ce9d0f7f4b7843a28cebdc58e870eb44b876e950e04e538a233c9b8617cad95ff9da336fb7103ed9c5bca514ed8b2e6f1cfee463081df771e1c0218f8fca6feb14169e43c14cf533a0f68b849351ee9c0f5b976ff04f7e5a9466432efd029f58915ca2b6e67cc78b4b662ee9146bae8ee073b98bf2e507a93730d3e28b2247b0abf0dbb9b1c91074d4c9b7adaef4f0e0d86fa162543d546b6fac6238b516aabc27188611e6a4782485ac971c03f5926e7eb8612088bddac3317677e20e44df01e536e411b422b302255187e00192bf48355e7fb57e130d292f82e49ed8a147e78a4b2e8b9d967662a2b0b3f930b028b8b08a38045ea70656fa46f528a5c8e99ae47f520db70b44def2a208e41726035ab0bd22dd6483a5fe0f094f88db00e699f877e24c99c6f1ce485284a9f9d71a1a1ab73fed48dd3369f71c2c0f7eb117019d8371855ee4bdec62cc1573ba823fd0cf72d398907cd8ad579e56e91e2eee1be9415cac32bd1d88276370365f2b5e9bdda1a3365037eccda53f9284fe27a3cc4264adb640a43d06a1c1ec5d49a9f0feb259f4acb3e38a017034dadd80e2ff8650b520d0e701f30c063dc26e0f9e9d24996e13e38549e67a9dcb92e9ba8dab9a6ed3d931bd0de52bdc3f25a5f5b0da52c80167f11062d0cef1a2188071c478f9fffacb9bdad6e4b0f91ae38f3c6ab63d9f3ac286b7aaf83c6c6ebd9b32bf367ce9974c3cabf29af23c747007f2b6cd113a351747b0187b8c1a5510b11cca73d7b1d4beaddfa08d6394e2bb6b1ca2b153863294031630cf577712394751394067cabea25d45fed560ae4332a304170795c955aa39afab9e806e97c3654b3eb150fc8a5718a1142b6f275a7105cbc78365da9064dd5d08b7dc7cb69a23380c9f8b8a570aeb187e7cf0d27cb4f6a3a202b0f4e9a83f0d3bb83d5e03c9ff22ebdef99529ed56c49ab29fea2f2fc89df442a741006f5ffffdcf499972e57d02084bfa050731ab4f6739145f39d1a614051d37f0019101314a65444ad0b6a8589f22ca071d6eab658dea1c5b9732b3d36e5a986435b0c8d6f83abf55d25ba143ff877d53387a8db4b765ae9800a2edc62e575cc7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha071ad3cba7c6eb1eaeec2b1e50af486114420f29b30f8bc9a28e2bc0935d364af815fd83c6c0e155cb0cd94b60a341097c15b98fbedd992f7197c4e3a057f19372a0aabd6e50cfe116e8362389f9aa91f073bac9c39f3a20f5c03bc6f1372d2826c0e87701f3bdb1ab6e628e6b81319aacc3d1792e060156920d4a51e8a192879653f590da54252f4198b7a0374bca206c435537750af86fae1cdef5b195670a84d37596fc146440aca85497844df4ad8568a37e297f67539aebff36adeead17b41514c19272101bcf28a9907cef110f05bb275a1daadbabab1262100d21e38c139ce0efa9aa3ae44157ce6c2bc086dc6d4b6a307880feb40abfd62a3f4ab511abcc14c2e3d580cc2dccd22cfb3bc605e65b65baaa1a24b679aacfaf37ebbab0ea0b3c2eca6da13aa0c8a4280421e9d8c00a92bd2371df10511ca8702d0598d00ec083074e055b077508d16e55ce99ad9b87b21ac116b832cd5b2209f5fea72766596f1b36451ba2efb529b60920ddd60e74e1fc19de32f6742cd8eb483d9cc6a5e9357cb19022c276a27483464be438d241731b130b01c832918c4860af3491bdf78781c89c1068c1351d53c02527131f134f8f04a3adbb0d47927d685be349bdcc8267459fb4f6ad4ead185bc30d0844a2427c060e74d333933ab36275a8d7be56b1340834d39fc223759578d28e84de3cf6bd62a38289a4f2c62e8409b8cbb528d8c1324ef2ebc47ad5ffde3fc6acae980415b65b5fe88b4973e9dffa3c7a98e0d4bf8d5af70bf6dab7dd29cf27ef530bf89702ce6dfef91af0c00c95ed10c9691fee158c9e95fb118f516a1aba0c81c616ee967b0a2850bf908129a487a01cff9c2ddfb9db9fd0d87ff5b3730131c530841e65423d8459dd1ea72f1f5b880a22bc8820ea0dcc11d71dd31ee1013577e1198cb0fb9218d53675390f77af217c43b6ef798564572a6899c59874697eb828f42ae21a21d0a266a12b7da5a9df2a078374239b2148c54b782156a9997be48bf20645c39e70d2166ecf9a50f8e681b5ffe67a1338b9b6536c93f4e546e8c085f4aed64ecca70c50233719ba66f447038ed3f99d1869d3296d94d34439b6691d52ede98bc68428fcb16191b311ff3c80eef0ea4f63177d44a713af2be9db54af0884f34788612cab74363a0a1d2db61e27de8e36298b75b4886f13e382ee7826cf8948c2a222a464df42aeaaa21e495f558fdb0517cd832a6afbe783795700aec10717c826a86d0d0d9dd0a13745cf28ce610dae8464942bfad537f560d9cdf7a5c2dcaf8bebad8f91f28d5139902ccea66bdb079ec8b0efaf5162ccebc0afa7dd787bbeb226c049a7750ef5c91c4ae018011f4b6a298cf06334a0e2b51a51e9544bf58d63cbaea6e6823dd186018175ae0d0c6ec75560bce4e2a65c4512e94f057be02ce10e71ec5cd7ecf1f13e08a86782b99ca1ba8fe7230d5fe61d2f45011c4347097183b9e5359a5ae3220a2717d7254eacd2e9aade96197c29ef2bd53ffdb681ee731c12a2116dac6582ae68eaedaa9ae36092dc1d9806612cc6a535e3ce9011f0e0fd2a5cc46ca5c3f0e3310302936eb0e7e7d5bcb00f5ea0048538759e47f3f21edecccb807a3664373582790dfb58720855480082dc705376fcd3d0b3cf123a55f9afe4060655f5be00d3dcb3cc8453856269ee6e3cede66a4a27a52f49fdf0db5c23e4c528e2830647874d55d134a28ff8061f0ce4c83e85fecee5ca7940abb6463a8fe10b85e2d4d9695ddb4489622fc918064a45f52cf7eb30512baee4a871199351223642858dfe18d7f8f6ae3b032b0bb15c080df5201c5179313ce95703aa08dc676799e70c2016b4282f241c8c72b9314618e796805cd156d38fcf182d873a0868b804f539f20ad3072b8418245072aae3669b233062038a535fc231120fe80ccff7f9f96038be3409d55135741421fd1d8b1e31a3e33054c1af89ea7b1302e13665a356997e3c5bc1d7b362fa5cdce6db71b53075812abdfddbfbd51bd1d24ef1bf8441315d6f4b6bc55f8470ab7cdb6a414cd49ec34e8f70f1018b6acb32671ed99ecf0866ae8d721699712eed9943955e0885ae7f8e35002c3a8018bc81005e86dd425e1f19658fea36eb2a1fda35546fb0f77e5e06d738582b2d2642b03020d8d3cfd22b1eefe762defd703f93d8d09966499786c58dcc1c526fe715941cf7d78a447f846cb6a23cb9dcf3ebccff16f36bb4141a3f64817c18fcbf5bc60d4e5b7e3ef23484bdf6139ad980f099e9427a27f5130640a742ef9aa12a74dfc52dd97f18217094710c04910359664993cbd9b7ea36ca362ee1088a55f5d8aefa7edf408955b2040e5e12e43cf162d80dc416af5def36ae4f0a6bf7ed3c71ba2ebf6800fd1eb092b60f9646f6923f97cde4059961135b86198801f7b1b0a055cf90af145490f627f85704a6cb5b381b2792101505808d867b639857426dabf553a0538ba16bf0f8cee0397ba275677bbdb2f22088ad1824868aa4c7122329b929a0f2ccccf897fb411abafb331bcb18f4c253349da85355fb28b1d0c76127dd48f6db7d15ffeddbd0980ab243f86c9d754929e69d5b206baafe5641469d280c070b04196c6f36b67d9c46f307e16d3521c6b8cc8351bcfba6a8307327c25cc9137bd7564fca42b447fc3c0cc12d7067af1dfe0b985fc219300f70f9c383c53fc709d504c5f7d673bb6c38871bee28809e670373450902082e406eafce52f5ea37c6809298d06832b081f656342cb5a4a682a7c39320529102b1021d165af13940a3b1a1c1ecec3dcc7a7f6b8b3e96f3c8cd84e4560d8f0f0f9dd1f47d44cff8c853d89fcca93ee8c7feea5b09e846459efb51c2f05bc85cc4c57f9b7b20d9a6e36e01316de6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4b917c3256beed4075046fa2b8d8329d7c16cc5552d304724fcf2be1797c9734e484d682ed06f48badaadf6ef6c920d196a1f314f5eef57020df2ef53e128598e206ab2958bbeddcf697d2ca752b021fcb247795982d1b48c8678898f8034769f6f718b4dfd7b3f23d2af2461eee3daa78cb29f9b93f9effb46021a6bddada7136e2c4b16999d780f64b1125b8a4e1b9103944e14ce714112ff04fa5ae7268686848581be75b3ea65feb7c9a6d9633dec73b7ef3695202a61b71eca9c519cf779f4d6bfc4271ec427a0f702ff5f4bb1e93201d967fe4976de16c2917b255af6f0040e45a45e0bb0f0361d66ed6cd0a566bb8603850566f1c27a0466d01a399119a34cc5d28788812fac0c8ce0fee846148746a3bdf6a164687c33e8c240aab2ecf68f49f977491f52a076a01e5c1c474be51f6e919267b4f0b3a60d3876f22235874dba1452929bdf280065fa05240f2e2c2bd1ec53204fc45e1e858ca31c8d71f230224bb0a3e495f1d203cb91ba3efde5519a9c8d18e887cc8a0b578c06eadfb487999020f74d0635f86c0d86a27cb55bf11a55d50b8a3a842509f42a995d17438ea2f62941947ed4adc8cbdfe1ac5e493e3da3fdbfc7bfe3319e36357d408da11ccfc1fe7b2740c591b2883e8faebca1834faf0f64d47486ea49d678371e13fa23eae68dffea73c5ae8b70a5279ed380b13a4dfde7fd8a23d305b6794edddc4a305785befc2c1af1421d8d5be270dd4399aac9fe2c1782d558effb98f6f884d6ff471b51d2a42c81dafcb710cdb780fa41a0949d1e3047962337bec9e3b5c5f652f760c69e0f98ecdb0ad9182e5ff98069391e1cfd1921147064a174f23b0a080fed16ebb33d948ad27250e5628e577684c210e181a6349b0a245976c6d16d9bdd1f74b1e71be2befdfac5713b882e05dc1d55f612646b29f1556ff0277849db35809a65a448e7ea0e3f0059419b8ac8a61eca12c11b9d496d9f12b6e478e4e6de93e2c7c249dc11deff90570aca7c7a54c8054b6cb9795fb2ea3315d9014a0f90388167045f949ade3c245a16bcd26a429f58ff917139b12b4d6fe5e7831843d02eda73f925f651918bf41f3ba8c617b3f4bfca549440e2540446544ea8946cdc74b9e13c4fbaf20bd3d56d8c4a0e89e10a27ceed08d61f4090af4237bbec39aa88192aa7a6a017b033d739f6ffe5d09052dbe1824b1034126ab2b9a4bf80887a797f4047760c763c3f5194c71699f91970294035a8fe09730d2871adb885bf84eca77ae67ce3d5987731cea9e3ffb4dd02cf28edb7119bd7ed7d84d0c716ce5ebb38e51265edd687e423b368c80cfbbe21d466f8d89b7378c1acb45fe6a0d6dbe564ce44f5bc6a37a3e5cd109589265994ac6c7fb72fd90433a7a35138e3613df30e23f803f762e5ca80de5a09ce039a4286e341f85a6d7914e02138c6f13958301fa6834c190683ae4222331f14324938de4ff1e567e9601d8ce9a3f7e554693c5494b7f4690227244c6df01cd5e35ef270412381c0f20be9ce2747baa509806ddd9d3f6d47cbb2edd5cddf4962c5541120e8876799d9047b03a7cbdb11a6f4ad884aa0ac3e6e07dfe14350c11095d309d61be872cc378d9e9dbf5de547bf6810321f233dd96becb82b9963b4c6e1218bb3a0b5736e3b0f3b9c765e369a4975b09b97339b505778c11540ce0e71f5592e35a6fe438392a410f0297a166caa21d982469923fb5db5a3215c865ba5eff99b2fd9985822477f81162b71bbc70c69402ae76709fc75d30e5a2d0c7cc8a5307f52301a6486b3c2c93818fe898183e8199b829ae43e8b397ad0ab5f38c50c01695a1a595867ba067a588c3ab4f2b88f7ccdc598c2e7b7fd3717ce9e0b2eebe0bf2635e425c19f72b4aecdecd62af7f36ca51b368aca1cbc437c9bc7a489fceec78fde250a3b2b93175b3ecf14013dba0200cae39067d63f4d8ca1b2fc2191151547c49b35e52ad801f44e3b710019ad02acfc8c9bb614ac8256ff82818e5d7427ff4bb71e1f7e0a8da2490028d78c8493c85b70b0be945349450b9b03e108cc43be5566052290e1956fada86120143931a1f5cf2ebad2eb66ea8caa9f45decbbab6a04af8ddb53ceeba09db4f5322a6002b9f16af36162a5221b7240404e53280c7adbe3993f3bc7aae5a960769e72578b8af91fb54f43d1337822fc3100078604f3f359a64c04330eb9b63d0a64789574430d243b1e7162a792ce97bffec7155e2045060e63c7f2418b71409d192c05b3514e498cdfa547de4b3ee4ca8a1e297d41a6f5509b4502efe32bbb54fb45500bea1de70371f73e24b2dae0dc6f25f8ce128ec65265dadb304a1b665ab0fa38edcb27c2be644544e917f438751bc772f6a17080aa493bf9dc8d3220ce9a47ff540a019a5a439a516f7f2206bc3fd9939d64abc5429b0b065ed9ef4d1d9dc307591f653e995124f69bf4df71ea132bc806aeed3fea27ad77065efd63277aade00ff07735f0e5b2b8f17c33683c88eab63f38b0475d381f0debae4ab12aa69e1775b5a4500702334943b3a0329c6135fbc16d529ffc0d3236b6a83861a58d934e6a84936e9016bbdea997b56dc170af6675414f724a73f39a3593df4324435e5f2e24e4360f05fffb22e698384439815d4cae9ff92e1711ae48885c640b33ae221af12c2a28c35560e115d8af0244018069fc310ca11f444bde51b6a97e6b58a8fc7d4aec44d887c604d4e8411cd4825dda2425af5a3b502f8592767ab72d0ccda4c9ac812c7a6a80da69ba178cbaad77728521ad1c262b46de4848e47f8378727ee29e8fa8b9be1751a9725db2abea57af66c5331570fc1c3c2e6ab11a865929a8317a2e81d69c2b3c47123d14985178714d0caa63d4d277617ee82a74;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4f19257abb79f9f40e19b378a1a97bae132a1692a1687d509c383da4a2776563c8fadbe7650c1f7fa93de5579f5c9a100a654ad85195244190a73c801c059096198eb27be312d298dfaa73ee276286610e2c9bb3c19c32855654015e0c45469fb609038b1599425e856818f1702aa76873ca887ed81ea44e8cd70340dfdcf4a148d867e400a29f1298ced9613e14a0808825ad464896f08761cbf7b5ea78d5531575be0ea3c907d4698bed510665937d63bd082636d07866085773e89041214f7e85f8c0096bfc4c3f78eea339da5e83a0bf3e160374e5b573593c44740372e415cc047af7590552952baf1d48aa82c73ead3fa78384927461ce915f94cb3eae2d4f23d04260eebbc6f8c3ccd8a602ff0a2784896424ade69ace8c226f6fd81e46b186cbf4f3953aee11e23f535bdb0614a6337721602386fc437f4c5d60cf9bd9a95612f532ca2bebadd43799dc2175fd07db48af817b949a385e5d1bb7dbbb0b4aba29f0bb5df8ec399d86899091e7727ca43e2b6abe2866f3f354b36f0b727af8a04dfed2b0dfa79cacceafa1a1e7575455bc8c4d3389038ed3aa4835e3392a366034ba3da47bc69d521c2b8130fd8d37573dfe43ded7b9de28bb48f42bc438c9782a9bf0ae30f2fe592cc710845345d9e94e49ca8f7bf6c550b7492998f2b6480c1de7727fabcbcf0b1061737d0fcef14470db9b63da0263015b67bcd0fc1f09f16e48f0fafad4bb50b5c8912346401d8d606bff588f361189eeb006deacc47f54478e5ad7993dbf55bec05a684f725069edd99283ee2d974b10c58332167f50039bebc0cc3718c7750bae71c2292e27ce14832e93247949a4ccc3658fa2873d522767a4cb22d8d95e903e85968562a750bf3e7ee79f1d3f803d9633add3a651b78e77b2af6ed6d1e70502b4a17f2fe3a7382f8da0253538c177d5c0083cae66d9d1e54c04a6ae0a869f6dc53acfa862b8a63b3f165c1d3b1fdd6e706935e8befdce9da05f55906813e9bd583985f81e63c82466fcfa32ba5d907615fc329a5539f6fda6df3abf1da6ea40ac22d70a458f3f42fd99490db2342766cf59c1de13e25a37faed6fdf80f56c59799b7cca6ec33a901e0958cb652e34927fea772423f67e2603a3d76d6df401a32328b859c4347d9741bbfce0d381aaa973bb208d3b64d406a7892278695860753a21192fc6f8d16ccceb5ad2fea0221fc8a415b5ab521c8f41cf84574f106516c6a0ced7353722738017215ebfadb9ba91819f49afe8d002458c3240576df4cd467a53954d01570fb087673a44139a8549b2959d2dee403239081a864fdd1925149a5f4f4781ad102d8230f2bf5720d6479309c8ad96ba7f59e02c0cb64c2412a709db8ee4bff9fd77f57134feb1521ab1beda208b1b71851a8adc9b3c300146f395e0e5ae866675b84a99b722a1212adf21ddec637345333f584a639faa40b524f38302a67627fe1f5542b2efffc603b1d6e56382df4daac32ef62e0548fccf022d5e7db69bbab3d7acfef2ef07a42fa2c026417d2c353000dc8916f9801ae9f278001de6cc494135b3b5d046fc51deadbef9b7819ae289a25bd272ce8e1882b23454afdcf3186e79573bf319dea7ef54b4bce6fe474d7d688291f42b46efc58b5a8bc1c748f1ffd53995da75a0430fee07a482d29e66c81e5e6242f290a424eb4ef3cab8b100ab8dde4a526ac2385e68915074145780e9147f3763229674d4c418c0bbf493c9225cda73f4d583ffb0af149ef079505b56109b9dcb73b8b560615045f21550bfd753442089ebc8cfbfe1c163d8ec7a8bf2881701c140c8ebb15fe7dffab9ea574daae3b02b5e9fb8ab3993d63199147958c4a0c6306e95743ecacaf65e25f872c59c38ce0f81248d632fbceda02e6b1858d0244252910613eefa0154f2190da4da15720c2644a85474d9dd15cc9356a65c3c90b62b3d5257b3b09d3fdd1ef481a3fdc9d90f2b94fcc0532754b026dc1a496aa7a0d2653703b75f5e5078041c5a51a91b7e26b92e7dc0ab6d061d9cd3215f6d19988fbf24e3547f8ea1d71a27885aac5d69eddb93778618c9e782f6c8cca0777ab2b6912cd62ffdd70dca9ccf9c108b18a3b18c2172d0fb1615b0a97f3975f2b740c18a64edb3e96d6cd85fd6b071ef1297f3bf5641b52f5f7bf74a8426bf6f7c7cc62b3410ba716e6523cdf62ae7f1fef0f8dd57b5e55251adc664f68619ce9bc0b5f07e1dd81c146c388cf688d360da6d21a5b12aedd44f2168bd167b19edb70d365d405f58fa1dcd6b489efb38dbdef304034243aae22921a2aa6ad41ef1ef948abf02c290aa2ba34d18364db1cf1548cb2a06cbb555375df16563144bea77e3eebf5f0579059d7d0371606ce9c8762f46e1ed018a85eceb8dda0e4d0d362caf3ba82470e236ab34ca5ba8407f6f4d11d6ca58c377b126b0e61f8c17536247b6a0e94e023ea0461c7329b9b53f3cbab798813f5adc8287c96e21ae788228694c84c6d0a8ba701c0c09408232466ff67340cc24d061de40860f61429455ea574b9ec4a50f471cc56ef38ffe2a9be86598e635feeff894080abb25a791067139928946d2bb0080c64f1e99212f8b7739bc28d0ad7876ebcf4fe63cb55f0a2b868dba484f2c8e71b51ebc17dea255ca235d0bfe97a0f2a4f512acf28163e9c77b191488dfba9584e16a5bef25bc789eb7a7b87cf3b9d92f1f6491c0a58faf50c331c420826861eee9a57b56ea4b6649e759e8200615b2827dfc84a37b8ea2904cf8dc9afaa97a5bddad24d3f79bb9b27b557c1c77577be99810e9c3bc3503ef176186bba87e7dc40b604a5cfed99505bd2e6a4373e09a00c1481e1f2c6aef63c493be1795b3a74d7a5f4237cc0ddc90fb3a4d9774a8c9a034da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd9005c6d0a7567298f8fa00473d5c19a4a3a3c091389607d00f59dd1e77b71296ed0e2780f29120cce18049f758963abd36c71839a77d2643b5f0ea951a72836eb5921ed193136881bced045beafbfe7e10c0c35e450b518829b151c57b003451cdbd577cdae25dd9a1408b097762a984eaf26f6344012f44a0b501151037d6396fa3f9fc9bbb36c219ca9b2a9ef332c53e28404cf095803289da567d5407b26359964b9b9e5615f9a31971710fe7314304f34d10fe26cf824ba07c9f72f211dba077275ec61720b217da52ac17aee0208372c48f929033aa0f92405d9333d349b3fe26c54d0573e656949a5f41be9dc706c82e5e62ed84b3b2dc3b3240200fb858879da123cf9d53c2b207d3cb99dfd89a09a4fc734301d787d99731d9984e03857a73af9a1e7e5578a328039658cedc609531cc2c46a8b3624752a52b4eb08d673df9ed55807f16cb99818d263278847bb05fe61d85dd032bd70f858b64eda04e66b37675f0252833a9176c84b8a89b43588fff3afc030d52042e561a23ab094400ecad5bff00a0de9b769d90de6ead58c760d0c58daba39603851ac68081689ca98849d0d620150d01b511e4d8e20968ebf1a1d771ea7a078d0640efcb180b02ac9f84d50e444420b39a665f327c0f8f34c701b3853a92d1e3a7f20163f690a10969aa1dfacc40c8113474e95da21e1a4ed7f6bc832628640354215d2cb88f1649f721d3007ce975ddbdb841e5147321ed192ce11da202c98678297bf4a0132dfb8ab00a11dca7d53783bffd486a3589f3a2ebd0411e043fcd46cb09c766390be9214bca59b7fdbaca2f5360241b63dc3519045eed358dc6936b972e551a058e5111bfc9d398cfbfebe9d077d0f51fa802be944654b9e7a1b38d7b6177f4b1371d60d8657565350374dc4937b41c4d6a9e17b11d96602135bc1fe63150dff351ec20cef0a7dbc1adb6c887567f55cdc609dce50fe703fc5960bd5bc2a6015f8563dce12d933f32bdd774efeb80691c7fc7bdb54b7add05884a2f2abdffa7e18734797420031c9d7f0394d552ccfadb2704608046bd3e0759c52fa3cf2f5082b06fffd9fee510df808b393dca3d6a374dbf4c91fbff9e7cd36a58eb0fccdc059de6b95edeadc9f5c92acb6b918bd44cd46f3c723f31ef0906a5ced05271a6d5d008d382568df3af760c62943d0e88c9c373cec270f2f3556396cfa92b5a9e52204d2b26bacdaad02cfcc93265bc9aafbfba69c585ac7fc006fc28e393ae80b05b1cf8b02ae09a7ba281d904b564a9e09212740e268d1388ca15e68702691ce8c4458856e27767949b3a116fde931b579a3e6f244caa2654efd738dd469b473cc0a0192ab06e0590df7d8bc381710569e81172d61dcc9deb50b2da4a6a5ebd2ac58772bcce6b1f097445b094cbb1bda9d3c41ef662004589dba73ec64514028607ccade10270066bc8da90c23235ada87bf7cd67af055c7b4c98b8f0fcab35ae52eeb101d1b0f88661657c43df54b2411be3d7d81108562ed7435d33bd77eadce1c0c5c79a9644fe6a2517edb7cf5126987a29d22336e745eec656f0fd41de1f1b0f03c8c0d1c11f8a6913257859b1e0c3b0ea2ce75df0fa292bfc40fd6aec538b912b16cc1b297d5ec6140e6643ce106ab18ad65e40dbea86ea9969f670d8eed6bf06a531639c7c0ed44c594dfe907ebfe5e69986523436ec508a5bcb4e065883889032ac2080da702ba5709ed5655577c4e88d4e2fc282f95b9b497eda4e4b806e5b6928dbd2df56e06c3ec77c6254d7502e59843e0da5cbd4f5f67f51f22eab25a4fdf5c8535ba29ca4476695a460034859f900f8214750bdc279c730e86f51acf01f9a4ecb9d82e55731ca727984c3f8b37414d2844dad25c2ddadc435566e12f3dd18b54af70892ef4ef05d3f1386e4256119d0997269bf98be86aaee699411736c62e46f8328679489eff08adf5adf4b2757d897d3d23b4cfc1d6eeef1d2e22d685d934d3612fec23d95fb432fc8fc8ed2e0f238735632b2c05c79ba0911bc29235c03ff4eeb7b855418c1640f00935127d5d50184587997a77efde5c7b4f22159890dc71e63515f2ab3a1788d8084f61598dc65a2a24edbd93c5aa82943eb8c96944d47c31c63003ed37a89154fa0d98edae919ff04274742f10173a33137c8cdb0d4739bb049cca2b46f50639456df0a7c3f68c886b2f047dcc60709622ae8bf91ed2f7cd0c5ecc958f9e08d6ad36b52f7bfae1db508e8c1d50395e748c9a16c9237d4f5e25f784af6d3439a4d6f4cd32dba7bf284e2d0924c572ee68579a155c5aeacc35a29398b91491211d2211eee9d08865a5a8fcfe3e3af45fd339c0d9db068442632410e9d0fb82d3bf822af3bca653f3557d8aed15d586d4d1f380cc6aeb9fe3fadb8f3b5a7151d2138da7559932cff5d026c4474cd2fb9f27535bff4ea1048bdc2be9d4066a63f824ce2cdeb7af090b39697e7ae6c152cc36bd7bd4267186d48d3337a0495afb122a898721dc5c52f8f3e36f3622a870f6931913c7b4b491ccd0414b881bfff7a73ad8dc29e1649b434bec9b42360cac10297013425be5bba85914398600f8af41502bb12bb9859a1361fb192daf1b5b10a956952bb12c89531271e9afab729e570f38c7bf729f4ee67d76277351cfc1b33915f2a679c2fe3211e1d1c0cf68a8cee4b7893bc4f33447c3c05aacf8629a3e93574c137ff653d8e76d358637b4fe258209689d03c71bef9d76009170b39d2c8bd76e3ea8e19ed8a8bac1cf5dfea7ecacb69a36f6996be71ba31aafb08a3eb7e8815a4d261d2bd3340c16647e20bc84baaae197860fbde689a5d4fe41f99b8658a019a55c148efd2782603b0d2bce126a1a0da87df9b62a3bac820d3ecb53ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf4efd3984ef32aaa16ab6608d99f4245852bb74d5ca270e4714144faf07411a915c5913008f78c7c44c6ac04bb1f645b727e185e547ef5eb445496d1063fd379ca44a18a8865ad53c277bebcd0a315606547a86396e9e329b3cb640e69a71bf8ca0ca60eca14ec1e160cc9eb093f6013772b41cd8ecf9861eab5b04affd9a4944fb503edb9d18c0865b22f3acd9cd65f6b33eaa27af6884464921d7807674a425e5d12a93c9a986af335d63aa58bb2286d77ebe316d52e46480d1d19a5845f1301dc5d96c8160b150cda6191086ce83060b4ae86546cc8ef4a1d5c48ee8d7cc93ced5c17f305f7a6a9b02a05be4bbf0f33974491fa8ef563f4cf4a7b70a62e747aae8d2f6383c34c4870f8b704dfd5acfeb1bc7b4b6fd6d9f17986aa0b3346aa850d443781f86e3594cfffdbb52974461f33405835555593c03b99a0739bf7ef337d6e95da5aaa6f6ded2d33014b67e8a58ee2f96de2f35848b9e88d0038e946c5dac3df74c4eb1bcf6feeae220d844b04b454b36392d997643a3907f964703f6b5c66b554c87146f20b0a795bdb47af45b300cb95d4918b0fa79c853f2f1e0f8064ec4e9be20dcd3355747808397c11897c3b2289626f1d1eb9f12444d9018f66db86fcbec3ba25fff3669b73daf15c56c1caf3336f9d14ffc12da7a27236754ca8bea2631585bfa804514fa807d7d80eafbd7580956d9ce3512a687e7489ee213b76c2b1b05ce47b59fa9d897d410d9f980fe22027811578639f4a5827b2b278a99d42fc79c9d5ee931a9cf9a98d8e2ae6184632a416cbb7057e126e4225c2569d5592b6bcd641cc421b2329f88f0173dbf0e2687564caa2e3d27f038d9f80cc3126f09605da816ce23884c4064638e7e5a5d59f15ba598f6b7239a2bb2cecd7059bc92add31a850a6b9c705ef25012007bbdab46739188d6c27235a4045d374383862b83d691bd7394775b03985ab952e60bccb9c6bc686a74bedb30b5899a6ff0c7f1200597c78744701955921f04d7c8c1df253184ab0752d0fb4eb38f07302c133d1385b209fee365a255f26175a8cd0f77a4f9b95cb6a040c05b85114308aa24968c6211f00d4781fafb34d3bdb4ab26e4642ec99db6fcd43a71be600807391d8c1afbe2b1e09f481c9c3f974ef474844d801bcaf257a0cced426596e5b39fff5474985c32fdd4576072251d9f1369a2f2cfbd12a8d9278c906c211dd7c8d753fc8ecef7dd052b960d21b9e04f12abe14ecc4b089065c412fe5ba765294fb28ff821f5d555842419fe4a5b73755f058b5d6e58d2bed94a586f732a3101e730747f43e18cabd3e84c1ebcefa2efc75f3eac4a3c39212a355e446f871c5573f70f905f3a9b3047236ebc5189cb4a494295884bd965b70dcc8f7a3da67c2057eefecdc6b742c61a4842ad563be87e02828e6eb59fcf9b41db92aee4bade2854293a9c9680ef9c3e669c2c18893a2871b6ad1df86a323d2a31e3bc0888fc38ab74a869d4e6136a4782b54ae9633c39c71a7d59298d0090fa51336b7f750bb6c87435ce0ca988515c5df8042da3f76a76b5d6463e1523e7ca63f615d8a88244a9aec162b5dba309ae318a12a6f266ae0c3354ac8dd253b92138aa6f025cce23209c749e737fb27a9deff63c6db936a8959bbb5602872c5f9a20011966154d3586ca346929cb2418c78730f380325dd3a107d829791ca40cba6de4875e550f5d18038557cbb7383ec6a05ee9613f0098b9cce0406d300625b517795961b39ddea6b62bf0003539c28cac937f8819728247007406ff555b05afe658cd72b591d5b76deaf15546097058b104b3696507cc84747be2c3ab9807dc0e850891d1258360ad94047818e7581ca4a0420f0f09841057899b039157a269e061b08a1f545a7655ccb38ae2c10d33c3403c9ee9c72ce6031264cef61a62f997683e099ba68e39160875651d547d493e2d5477587bc595a4946ec96cde87bba29cf89921987b402f61e574edfa22eecb1a333861bbda2bce0d33d7f03159f7805c027f99c5a34fa3fcb6c0a0356e04e6975804acfc0c9d0cc0b4627e6a6e9cd0dfa8efdef650b4ea1cbce2cae41206c4ca1a23fb732268b13d25bfb92a415a5eea8d77be6542930d91210b23c37682c095c67cf07589e78a8ca3a06a5999078e6c04c6c98574beb190a97e5f95a88523d455a534b128d356137ba511d1ea23898a694b1971c5d5fe6b9aa38cf88746a146c0c6b2a1c2bd847e8ce48e648e2e69f5c868b5718878677367001999274e06ee31f1e31b7a9456d35c8d835ec4c728aa9a7c6b06e43f2bfd756fbf9ef73efc7dbbb2326f4b6cb377e4ae5aa801e81aba86e975a0e329e63b9e77818c34951414a8c7294b47531c48feef3775081e09ff8380e86b4ba72a54b20097eb86ad4f5fbac1aa2e3ba2c05849c422941b5de4b34c4d1ee24858c195065f4f831c5cf8ef1d3eeb8b14041c7e75874702defd40a1591fc94b3eae23642844389bd3da73c86803606aa92bcdced44a101f6595a34f56fa9f4083f3b186e5f7a4233a1d40bcbe32c0406d81909a51f8c1f27cfd91cce015e343cc7c6a43284b77de145c275546c001fc4499640deff488026c382620d4586bf22771a3c75bbfc1a5611b973cdc8fa1e428e4115dbb6404de91b4abdfbc6b3d3e5b1ab636c10c58fdfc0c13f4f31ddb9b7160e9f9d133b8bae41b2a3f155706d05b05814a11388850e0139951024775b29fdd17e8d042522981cefec917556fdbd514f1afbcde55d9b46fdbf4b22985e177245744456b4288467889a9b925ca6e72201958898b4c668d7bf20d35f3d72802d3d98071fd4752035a7339dca0eeab102956048e5a335f920dc25cfbe681225076e3b34f0002758586e60b253a9bbde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hea5baf3285a5e1abe6977f82fbaabc3415e3028d8a4897712b800a9053ecd7d01ffb31040b04aea34b8442fa2266f26f010fd7a1269f9646fbe9f0e82ab1d88de191fb3b485196950a764c1c64e3056233fefd1901338baa08b05a2e3d9a6095672daae2d860b2e78e808194baf3cbe1b34fa2872826f5e0493f9349f39642e8be348b1404b152e065fb603da9b364f789267376c7feaa1985195499f183cb0b7ffc82718f8f74c7cf4cb7a393f54ab7f3af192cd5b8b1cdbb7f04b90034ddbce697a7b46ce88c2e6807c0c9bd327898f50f27767f12c161731ef605d93d8d4b0d3519aa4d3c0e96573f55268577133f473affae14eccd108cb4bbf18d9ea4a013665eab40c96698ab0eac073cef4b71cca97900ba51595d3ef68496d36527f91dbc2e32894d214097e6b8e015d411d1e76381b1fa74d25356bb22d0b1142faff08a274d72970cd1eb95a1e68f1b3ce1461a529125d84dd9350b504f6c9ba130196b5a642e22a1b4c68e961a9124c6a5f021f957dcf8e463a4369e3617fc13624ab0df428e86b9d26808cc38b27aacd26f7d3a0c86d611d1617bc183ba5f9e9c692769efcc7c16a63b811482a6ad1b0182a4c0624d7528b6b822b15dee54b1e6ffd6ca8885faf50d1787ffbb6f5b6a081bf69243bf8c2cd7af6da711898acba6361ce86c126d3341e429202152ff0f062eb00e2b3ed5601448b59e3acd2f46e14eeffc2f3ed79e3ad839b23974f2ee5019fd122c89d222b5987b37729d9f812cd9d58ff14e1e93a92041ef1b775eb037e5ab77770c7a6d8c4d86f96800030d6450823c2325e6b6a94b32d42934fe91ef1508ae22e0e6a43386c0aecd9bab645a5bdf664121dc944f285c90a876fe6e1e16bee16f17b22eacee1effd0e133a79ad8f961939ddb9a675ab8bfe3ee5d2986b5e39b9c37958a08d0f7f531c03f6e1ac5131342ecf89e61b49162c4aff9db87b2a69bfa47a1c1c03197882f9f19b8cb990a9257b9c33df55b5f3dba172cb56eeb19fdfce451b3e10170f52ee1dcd0c012eb621ca5bc46596f036a409d2a12f0abddd8aca58f04fd7d96651d25729ac4e9c05f6a91bc5b02dd2c24ee32e08da80a7266ae008f5ba448c3a2bbd82cbe03dc10c927f630574a3767cce0019fa1f3b25cf42eb33f089043633d5e4fe4a55cabee938f42b312e8303c2b0e744426e6faba4091ea9bb1aaeb0282271411749b77e62fc858ef6153fb5180a99ea84e40fa569e5c921683d13626b3406eb1d79833bcd6bad6b6d9d02270639f22e8b5df185393871eedb3ceac1c05e69fb3a3ba3145c87ac2d65244ed793e9264a0616d9237bbaa8f655f84655114ee9de42679d6ba5413b3660c3dd4835a5e884b64ad4cb76838c99cd882b29c6025dfb32854f6e3f051adbeb7d6af2d0846e3095de5d59c9846d9494f21a5c162e01f1200506d807f321923182f0b6bf3579158925e6a4373cc08bdfa5e2863c3f3dfa9bfd47f6df3cac0b6b55bb5d9f0a3555042e374c4bd09b4ed023f6900d8924f69bbf2b4b300d3d660ee96e9ed9b20db36ff5995b2d863eb7484c0f7d2fa454d0ebe08d5d4d49b7fe4a7e103861fe92fe926463b3a8507e6eb823055c8cfb569b32ddfec683e8ada91ddccf1d9b6b28611ed4c4dad1f83a77241194e99e8085efd8574578adf14d3350df17e2eb25403ae7db5f19359261be96cea705d3f5ccbe99707f82928cc510f819fb4028a49840954dcca94290460e23c66551e4b1195192f04779373ffd68c1d4c1d57c59ad30d20a3aaca26b6ac0492939f86a3956f951e3389d3b900aca4c0265abd9dd52aa76bc90384a5af5722062bebf49e3672364d525ef837c2964f8752a6715931e77f178263fc6a27e7e737e6267fc9089ac73dd1208aafd5efa72e433068cf3beff54b4b2821e30f0a7a12c15145431e4f0cf39f052e7e1ec348965412b9756777e4979e620a09be000ec76dc99813f43a73cf6a400f39d22eebbc1fbd0e13ae2263bd657dd5c12f9c171289175eacc5fd455c25d4f2d26394f43724eaa677428fb3bc6629b9e3ece6572704102efccc0f2e63c30b126ead1628ec730cdd632e3a83c7527486c5eef09a3d97c99c47a49f231dec64da4fa8e2ee73797360a4e299591ae3fcc10c9e814537b0041dd5852880602906cfa55774ec4fbcc0e7969b2380c5b00fd58cd5c6f10f1beda7a453ba2dcbefb31e41bc75ffa18ce0f83c816821fa4577e5ce0f7827e46e287a35c50520d6433ebb3c04bb6b0945309aefd81e4ade007d6cc781c7c81c526b6e61be374666d6cb5d7ec7ff1809aa2e52fdc3b619bce662b271cc8fb0ec8215a0cb70a8dd1ce5a61c1a6b480068476949e4e5b42abd85c5dea6e4005f261eb57609bcdbac21e8890441aff87af11501605eeb469ee18bab08eedaf572fdddb22d55609e9c33341ce9bfb0c0923f4e49009618e05ad4f64de63f1e646a3581c863eff3469876456cb06e7ccf516ed841a8791db319f36f1c2838056ef8df4f1b2c131489f5090becdf5dd34c6e2b1456f196be7c3be8b628509d982560d65da3a69cc38b5ef5bf43c5845cc8ce512afae62e947dba24613089a4ae25d2c3a2da9250ed9f6cc37967ca92a4d66780a19041477f4b119ae7482e3564d21ecf973121c9e5c9b0d9bbddf9f779fdf47481c8eb47de300d5d8af3665d48ebd38e4e92d787afc3845a6a6e0700fc64cb69ca09c4f40248101a8c5350f0f732a5f176359b1d324fe09771a84bef102d2405b77748aba93a99ac2b676e48f56b0985eb1da1dc05698fa872b437bb5448333a7a8c47c76be3a41bea0733d0a9e42c93412138e8c1a73a3ed9ae27b5311bb95a8e2803f3153692ad0f7828f79485ef6903d9b8abe2249e115;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he6a5cd10d75afd6d9974c0d33da14df5a77366dca90251cf60bdaec050b615b198151ef05a62252039a3fd1ea85315b7c3d0e77b54a705ca4cd09f7b9fd6c14b145c808e91b5515a5a7c778dae177faffe73147cb5fc5dc87ce72faf3f25d2bc6b052f97cb63e4ec1b3ce219a2ed60a899743730ce881bbc49397e3786328966f2d96dc2c55ff5182205a01c17036f365b675bd09b203bfd6ad84eb6d506ca26be28e45f408d4a825f9de62cc43dfe146ac8bc39b4998404bdd344a329c54a8dbfaa1d8c2dd9f4e0e6ac66abf2c411d63ada55aa162e802cdfdac4a0dc9332728717d24a7b40eacd7b637a99e1d9ae0cff9118e03b8188a7a17a1a4dd1d60f17d17b89757dde9f8943cc5ad2e17870591831521c211453264e7741e679184b9a72172c8ab3f38c90fbbbeb093a990d5e91fc8de6fc86492f20bbbdefb293b9e38ca3efcda7e254a69e1f75962bb58156c278db89619888f82a4a8b609a37e37195da9181b3b031f4d0b385061d0ff4435a586ea04a5f201c029fa05c10aff0cb782c542b0aa954067265d72ca6a913c28d3dd0bd4a8160c859f04fffd63ea03924aa81e378d878f25ce11ff21786a4f627ebce98be61fff8c23f9d3409d5b6902e27555c04196cfdebb9ef440160f0dd2ceadce9394bd6a0af1d58edd53599eba9a5c5ffb92fbf45d897091bba22ec290e13b83065255cc47486b1937e86b978eac07c8b014b8808b77533569765b658afbc811ae72568268eef7aebbd29b92fa813f7e86339cab0e6203c21c04c22c1a0af281b6b73ec437b73c8f3a54a274ed4b64eea76a86f18a8d1dc71fa9b56892affef222cbae87032e9dbc8c8b5ac92030aa23642ef459560472ade9ea39e691b224cf143afe8f34e25f1cddae31fa9975779658fe6b061f01aaabaddf6029de98b28598783185d1c06125d6fb2b21543aa31f661688140adf993a82b7985def7527af912546d50a15e4430db3e539eb0e65af6a39b921ad568fd88c6ef17837a963e859f26f0dfc4428dc2cb0affd67eb44d7277a3f58fc5a7bd9e8620f93152aa9d7ff5eec49c8241868907a44b5a74bc530359177819c646c675c2a67e810a6413d7bd2b21b7e7bc60ea76d06288f8275bd2e90e65941a0f4778d09bf922b25ac1c6fab653f2501b1b0412533078a48592b57edce418fdffbd4bde16c9ba87d94771d2795d1afd27d8a0de38034d21305115167fa351456500b94af1d4b9deb26eafa6d0f33ee775f6b1cd486b261007d8fed49dd98388154cb253bfdb0b8e493d5786dec457b5c9b4a579ac0ca940b8e594c0c5f8e93bae00d5fd164c259de818db8632d565aa2d257285ecae3656e71f0913cc2a95261b5a76f8a6f07c67c8f2c89324ddce353fc1351eebe168d5e694dae84120c6ce802f51879ae69ff91ecf36ba9fadce0e69969f2286c42206adf553fa26b286fba027e273ed150c20f60a0f8cda66071c5bcc62f0f2ed7ff8fff226d26750503c6da4dc4678e04b9197cd32d949a43642ae8ad403dc7576089bf137d3a632e22c8fe459865729f0de5ce38abec252b443c70040de72d9ff286dff6cd5e2d186e859fcde2de22c8e9cea25ea527b09867e327d9046c2826bcbf80339609bff2b6119961fdfdaf8d0c2dcd14c9ccb3184952cf73c73e70c790e292e073d6cd0f96270652ddaf40452ff49855c71a04f0139bd6ae1a114a3732e00dfd13c84aa465b9b2ea88c9599f6b60d5c0a5829cc92d2ab237f0b821d7f36a8a1948ac13c12ffa9fdb98d41da50ce4e36aaf80f1147b497923e5a5bbd801b6872c1a0ecb61d6ffc200d270c724179d600b1cda4f04465420a86d59afbd0dbf7bad6b80c1bfe9e0166dc137fb724edb6a74ff158d6fe2a184c47ee34722458eb8b7799f368cb977790d3b8141ec9c0d4d17dca64a1f61f04076507fa5c4f463a78d96efe52795a6ab015d7ae60094331f08398c70f35c541118b14d4bf7a790a6d1f7337d794a404f6da3f375aa1e9fdebdb93bd78fd50860807a5572cccb6c42633c896974764c0302e2268141b835475b667e216ed34ee7048e1a52182362a551f7ed84e30aaea1a59a2937c02b7e09cf745b450618906d49068d4f12f72fe64b0621ae3492ecce3ca9dff20c872062d3a5330fa3ca85d903cada8cb85d17abbfd3a48ab2ab4a97cade7fb42598f7e321d2083d0c7df1ffdd58a9de95d4e69d0032e6265c8c87b6dfea6e34e8c94ccc30983f06e3995bd4005c925cff65264b8f317cbf37b044b9eeba7d5c9d5861a3a717f4549c053fccfcdc7474589e6d095d72a6778275433478e9fffa71436834edb1e6df6415174bcf2272c54d5ed2ca60a9672cd0551d3603ee01082d77f2cb9237fcda6d65dad67fe87253feab819dc84eb55f4cab1492f93cb929abcb33f7a6760582dafd5d7e4476e3a0b6309f582cc5f83b0f91516427dd22e6de6e9af54bc754a55e6b00c3b7ad9a5a4e8298d33285024dc92638e9ea8248052c0133061a93aef09cf683fa9e74d226e9064bc4474f77313e65eefc69cbc72ad026d2daf8973b445fbf04f89cde0792418b66a9e4256f34578d2d60f512787b91bacaf848c64e6adb49a87138fe4a6ee29f8977d45d29ed67ccd13f9dbdb46f499712d29f747926e5f05d680d90724be6609b9ba8e4b25dae79a517b9b385efec7b591d0c21f192dc07e8022de5820efde4d4a85b6893eefaf6eded809407d171a5c4d8ae48b56714f2dc2201d00a6ff479871c62228de2bffde022e7163e29efd2516be83d3d83b005b39c67a4951a9d005d7fd34e8f6cac2a3ffa8ad3b522f278fada8c6def7acdbe4ee8fb41a5006be4c2a1bc5c7382d4095b833e5ac0f2cc8e29463b205e246ccb3f1c5630420b184;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h672b2e014b5b84d11ea3e2e4b40a11cee75b3a1d73bfaf35027d57ff2c50d6be050227a3d306055dd62d8fecebe7f97bf8238f20c548a130c28cf55cd03732f363ffe18ba179a324948e9efdd7a33de0898404313e1c5c20429c4a0a41ae1ccdca555fa716cb084cb45533796d403ae24799cee98524373f01111db55e50cbc9230f87bb6c832b306530d7c573c8fa0a5f0e9ca4839756c4b53dfa5857fbbe9f12e8cecf49636148627d1aa5288a0e5a158bf3c4d53520216c87f46f58edc94c18511ae76a5edca519503fed874bf2ab092654190aa712c556c84963e7f6d5c4e08d242f8ecf58ad797e12b39af270dc64a5db1245649a62d4d35b29a4324d1bef1bb4be2892bcd602e6d39259324bb5eda9023af34fa4e983307c1a27334bf006193a1ab4130b005159c3bb647c59412844fdb98214a9559e04090e28f33a0fbe47d866947a96b47526a783ff9fc3eb668badfff2899f2364c97a9e090a50d0c50f4319505d0e19012ddbe9b39684eec53b8ae934e4a63f432449a1aa9a3d91109a69de5c5f8ffdadc7392af0aab40a00dd9fd661f419dcdced56eaf3d476903d49b800c707f61b3e39426eb74a63e8fe3e3b1a3fe5e606e86011d2cc7faae22dd0abf8f8f77d02569ba7c0fc032c757eb03821a4c57ced0ea1847331df0c6f3ff289f24d047c4159d9dfb4448be276df34e6aaa955d2d3414524465d6bd8ce9c20173357e491eb37c680515586094a056507d03935a016a74dd068f5cb6dd8cb0e53e7eefe5399469c05d0bce8192e9b43dd35bf71210ed15e6736a12cdd93ba880b0ec4e60f5c34dd393cef537bdfa3f2e1e519cfd7dd6d18c3e805631f60991acc933a3e33e4f2a1bd0f60f5da5a8ad05f094ed530f0e9a1e8e03ff9e25e7e18ade7693dede5519a502115d3d7e7346e81983be7e1c69a7a151bd5784d50955e8ba10fc73f775061f4a3d0166d645969e61f3a12045ae03f51edd30d6cf5f1642f5d9d0839e995d3c06491b75adcf9aabf806547614594d0faa01e50b0c896dd7222fe1320739ded4355e3c8cbd43b84dff06ca56c8b78b4ee93f82ded3c9258216e723c90692b09802a2fccf4a37a2865d34d30953db45206768b7f777b582a6e39d4949d98bdb388bff50f607d543da7910c9fd9554beff5a7ae9da985a78327ee60fcfa63708f3cd3ffbc2bb9697c062b920c7028310f27a7b1d013903b1571bd8604f52c4fd64f0c9a3e266b45c85c1dba9e8e1e76a3aa15f4bd74c811f20c599924667f3d6c4cae076d7944f027bc75fb98b4c9eeef38034f58470117811a719443981017acddf1ecd4ecc3e3cff6bce8b01200d7917f6185309732dac1cfc27e126aa1c294d5dd416a93f70cb6cf7be0a28c2b0be8da5fd15c9d8228390560bddae8a85a45eb00e7b4ac77bcf105f94cdf9aad45a1c46547a18473ea7e110096c2b4598ca3d4b31b574b7aeaa908b4d70f42203e6f29f3094f43562619e2706648ac427453925a997f8e5ac4e955fc4ffaa8f795b3174addde9c3f1779495b3590eb769c13d5362e7af74fc62ed2383aca601aa02cd6be1e21e2cf41e462e5194e2a16e007d0ef460b52203707ab2ab126752b9c2879670b99fc7f63fa144588fb06f5992b27ffc1e065ba4e1e36d476fb317b9c609a9f20ccb4c3b42bff65f1f378ba1d5d6b60db71b2e05eb6c76a6676f2dfcc4ebebe68c7e36bfd8d03e6f041d67c60d70d35e05338afed497428e0f479a8fa14b5ee3429bba5fadf676ba125c78b73a7010cc2da0f2e812248d81fc23a7fd77932b7a6c86e28118dddaebfbf542fe40e6d5be5c246c014c73ead479abb77f09f80109710a37615185638bbef28e01f544d3b254215b6b873e36712af11a7feac9376f5b4c908deb41c10f4fb5ab5f7ca3c83b159326c134476d42fd89f669e4eebb48c5a6b49e591f24ac0a629d087382b26ce512cb19635a6252a5e0041c178c62f3bb3005d664e80a5e4935aa39fe28a580c8f3dedd4be5292e694c814882b30928053262c9fc1dbc17edfdf1186326c6530f042ec7147b39e3938d761fb20657e59ba2afab987ea06a2e2aa682e4492f409858c0febe0b755cd10147ad7bb122286ff71ea4a561a00163005f2258a5982f8806c4fecaf1e2131ef9ad927e9bcf036adf435e163e3fed385670273ebf42192b8e630ef7c63bc55e419bf064f258caf48d92518c8813673796015a1822fec4d8eecc45d8bb15c213a6f8e2b221c56b24d0fb2cc1657a062f644374cbe819551e833702d32dd836ad963cce0cc010d411062c22f595dd1bd7509bdd0c825b5bbb1f8cb805897a19e454170b5ab0c54718abfebfb219c94f5d4e445476246523e704cea38465fa59eb22665ec683a702db128dbe1aba2fb476cc23da165b4b10fd2a56d5b2d2130961f0c824f823c460912b07a650d7fb19e54ae158a8eb36ad436804ef0364e5a367733a0fda16dad046ba95e29e0039279c0debfdfb4d59665491a412f0695b74b4875b7f61d7add35d5b5b46d72eb91fa0d1ae66e8cda594ece28b6b79bd40d13352d979a6bf49e7bead0c8cf3445cd502ae25f52137024f1a5dfe32208d71a857eb82edbd761297ba45768d2109b905dff4954b5d04e884192b8f21994caee330b701d035712944975306f83a8675f8c1f7a70704bca077a2ec33f3342d8cb1fc24a69a01fb7ac30d677ff5cc990a8694b9d2efd581d4e6a50a63b21ed98eeae9e207f105200f807a3e60e38382f771aee19949b840662670e9d1d7d549b887e78585ef2366de6aa36d37e1c7fa744965443aeb540cd60e2ba54b7a215a720916cd978584ad41f380304b0b2c4b60ace63b54cfd24faf4800a665ef74e88ebc8b0aa07d2a45423d60791d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9c3697e1af78ed8660d5545108b174820ad06a38389bed967444260714579489c5d994ef3889a1571b95f414aa9280f75a460e2929479109875abe47d4d0b017df0b1edfb1f443c0ce17d56c251c1db396941560f30704c49a979c9643316422b58a81340e777409946c8d12778fccb66210bb34e4e10085c1f90c8d934ff82122f3c1a706fdf2bf6837ced706cb486f7e7d83b00a6f1b89b16ec4259f3b9f76816844f8e90caac54e3d6762ced6f8aef348b2be19bb070a3eaf5c6d595531bb50d72120d692cf531db7e78788096ed0c90dd0a101d3ce358ba07685a51d4591ad2e56b857886d5380c4343e6d836f105f50313d6c8206cf593b596b698299f9f9269f23a1e65100d991dc390927724ab622d8d74d61f208271e96a61bbb73cfe6620d9b8b76c4856f6d470710357b02410af2f8f70e52debf9272e1c1d09c2820e7ec9dccb829277d35f9fe291ca392d59d4289b4210c06be45be7109e57c4c6235fa084c1f515ad837e501918b1d5f671fc0f5cb35b3099efef2a1106e4eea85a546a76ad66480f9dface794b44d648b189a93f4ef6a63683035c84b75e113eecdd7fd7dfdfb352a6301333c8de11b1ca2bf5ebdb375b8f8e1096f39b648cd73bdd8ae07c69257b1ebee1fa7508540fc0c886e2a9332e61b81d20bd561cde5e6d93a6450473f4badff1fcdf63b527a5dfd383f36f801602ff8139590c8cb5fb398cf882864737cfaaac3f737d727452034ee12c8729533d9143a9dbace2e9440995c3b000cfe42dc84ce05c05edbd4ee199cb44d562d1d849cabcb776876a40cafd14024454a3f6dd5e6e779431841bf9c79242a0473bd953c9dc0a262121c9850979a0c4ac775f452cf6d3772efa6cf5e75f0af5fef4f7fa4b38533adbbcbe77281645da260a090e97ada3658ed81e9d3c771cc78fe4421bd096e63a35a1e2002a67311cb1d8927fd60b2d398e856fcc96cc1fd0cdcf841631ffdaf25496dfef008526792ba373db1d38ae411cc28ed2b7cecc5c6036dae1699b2b30f1062af5c04fa35716ad5fa97106f15e36d998cbca019a5cb664de739bce93774c18728d15906e76e14cb63702529eea4efd2470e1b3bd1fd38a49a9a8858ed0258d750d584835c8b767252cfe9192c407724e105fe8cd91ed7b4138c829090e180b533b90df37b15aa53d708df08caa38e0bffa7e3d3cf5fb6b96f5daabb8d0949fbde6dd1efb0aad19b7cdc582759b5b2939c1da6f42359494375ec67210be5f1466e3fc3781c8644a3114299933b99d830bb299b43b6368dcda981c7c13166724182912ee8f19424f700bc08ee64bc885cadcb62b852dee9a420003e20600cfe1fc2967eae150fb9182c646e656130f657ff2bfa11bac399a651ed2e04dacf6b58f5fa4797cf82a77c95ae09e5c82905234cd90636c34c9f0f296387333cbde05d25cb1225519ef4c3fe810e1b6c7177cf11a24162039c46488e5ad0f0f9714876067ab67eb6af36626f237451e20f047e258101b7e54bd7cd92f08372c5b4d9745c00de56a160bc48a1700d04c87bf492566633a72da2607cb1f01a75f627c83ee0407bd1e58f342affe4d4218bd30efa9509aa7042eb3c1f2d5acb99d0c10e57138e587c11929b0fdf55287cbc6f39059594864e7e9117ebc51f144c7b7882697e59e87911497d3eb1d1882a9bd5961ef2eccc4b34e5a0d7bcfd4284b91adfb43adc1ec733a6efc207bdaad96e56d5225dbe4e1dd23feb3826d5e8a2523176f2e1a14f6580ce16b1b8a1afac70002b3de0072332e5c060730d466a7e0ba4ee3c7b6315fa9b2e582819e126e491a2d630bb0660084424dbc4a78c66a86c72eb48b4b8dc117f525dbc0e2ffb338f509ac7489cc86ac406dd545d9b453ebb1e37a57f85434cc780bb92f9da4644e1d423f21a049193b31cdfdee1c2ccba7f3a4b2b09d20376bd8606bb34d7b99b17fa6a4c7a850da1df2ca798963f66b778d120f04dda21a361ee8dfe57c86a4f78163bd9fb122b5d4a2088a41ab38bc8039a4456b4e57498aab692c6dd90949fc37714ebaa21aade326fac6b7be30b71e8a4cbd1c8840eef721a1d28910bb0d28959895f26279efc2e36b47739875433832e1247a6a719d2da7c89929f479fc08c77e4f2cac0fd054d6be23d389b172c9484d291c38ed86aa6e3332bdc48e13a0355849af4a09baece71a46a51a7eba470629b2f06f0aefc0883e870f36178cbae45f3457e662800928cf76a5ade341809a19b1237bdb8dcc9cda1763240595fd0d9773b211b02421f7031969e3ef52d6871d5963fd2490a3d2b338752c6292a0ee613b6917f6346bcb8fd11f0b20680b8b9e82d5468032c031a31320ef11e5461890a8aebf40dac720302557fff730b2fe3edbfcfd46b715dc84978c83576701c19ee8dead7f48193b4d4cf32a4c6097cc5bc92616e5bea352ca55e48b148e4b8536f22e8cdcd8584c6725feb1733dc77d4a9ad69c861811cf69d487b593b4246dc2be83f5fd9a56623d2dd7b438e03d338fe70c01b1c9bd944de3fb13f9a265258e1a17a727e377dc4c0f8dad61b8fee0e56d524e22b9304b5aa77abdf4fff3b9e3f5a351feb21d07c3884b6e27e771a3edf187b64ba8f016c32b0b754aa4d24187d1ee2d208c72608ee151424110a8662ca83e06596958d044c6307b8983ebb44d159a7087ce6a8a030a0eed8a95813fa44aea850a15d9e30cbc57b3be541a6b3f7afb6716c2bae679ea06125ce8ac3f7b87f687be043aeb20437b75cb83f605eebf26f934d5cf5ef42c1b0b4524144971c7b4ca275bb0a160cb6eb0c991b851d0f576d372a585e5b55f47191b0407a6d916aaefb87ddc19e97678ea6524aabb19f2985551efda7412d5b6b4e48a5f690d012;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6c964e13580e20b14930011dc2098883c3ee358584a61620c813d45314fa3b26adc61cbf19928c95124f18f38b5c9f87cbd4aa61c9acd9a1fc838569c226e61f3cf425f20d03fcfca5a8d5c1de08b909543fb564ba13904271dbdc4da26c9335e1e40153117d55fcfca58fbc18c0a8cfa8ee01d0fa656d2878b1172cf44a54372467f690ac2ebe698df6b0254f3c1d65c20183e6f6c7b7c0d8da193d27ed9c6980f76c2637398f127d3af775d4ae3b777994129f3fcdaa4a0a4c8d34a95cf7077867e3af109708f1b1811c8bea9013c46b34a1ec86e3e2f8fac9128101085e8baa5f7709aae99e16d40ccfbf60dd118823d32909fd90f454b83e9eb8bab472cc1a2d0f3b0ebbb88c3d711c7f21bdfe4010df1ba9ca9679ff10a7bc381e98030ac21b1efeba47574708757c8bbe454961f0b96d126aa6f1af58cd031ad499cbb15253cea9fe12089170a2fee93d8cf70619138158a22b792ddda60928b5f53e497893f38ddbdae5b124c059335ca57e8d4370b4481f410045e4ae84631c00296e1c1b6dc45ff201da709eb102c599317bc7d1d75f221f06414bc960569e6f5beab9a3431a25d2fa3a9c125a2be27d5aac340fe11ecbb8c99d245782517de1429dc2902efa27f0e12fd32a9652072993f727f7516d6a21a8997aa5b88e8d302e47d20078dcabc02f617cf916b7b6af0eb6068efd117d3f8c09a575bdd727ae68b4c489c6346ade20d2a60e880ed03c402adb54a2dd14b518d4f626ad869642ec271d92ccaa14b1dc8c30f3ddc399cbd07135042da57febca9fbb7fac5803ad655897c4129b8aa2f53bcff5b027281486ef8d853ecdbcccb813f8cfe55463381879a175f12770375c02b49349d551a3f64775c2b6c508d11ef1b7e868dd128dfe5fcb153aead3828378d61bc46d0e13b2c2da132c494c7ab39e5ae4a3a6b8a8f202f991e2bbbd42695140df242a9533dd77e05d046343a4a467ce38a41ca79d408b127ad1a2fb0c80781f3fffc2363bb7bb32c4911e4fc26fd19b70e3832689962c813e73d9200bcef1cb44c20b921a7ecf6c4376f99f41474f87690badd89fc2291a98384abc14ba829fe5b29ac2bc9f1b5ee709cd9cba6f50eaa52fc63c93f88f32fd870351a2a4dde767960187c3e6856b15cd45e7217c082ade41d8f569076718303258f19904080e43d065295c0dd89ee15981bb98bef990c62147be804d62cbac146fef79ed020f271811e4d24cef23b3c0404896df8fd3fc2f739dc3125007bfefae2b26b5962358f5fec75a90dcc7082dbe08d1594003a3bef80fbb48babb6b734b313d4393693470d0b6a16969ffd20ae51c04785a1c4f17809e33778ccea637e105a108be219e7061ec6901961ee95f4aeb2b1034f93fa561ff604e060c51167a1a33f73ff3c86495663c95c516b849f1dac99fd7837afa5a6415c35d5d5c22236b7297ff1b7fedd0977b97d448f2cfe35794fae4f1d6b6529ef8f2f832ed42d293f3abe68efdadf8372497bc81877d97bfa3835501addf982bb891f3be50237744752be37c2d274244ca0a2e96646dfdfee7ba1f86ac2898a4b4161f08b0dea9a3e0ec0dc69669115ea8c185995cb282770ddc94398ca29ff27d9d776c6e52c910bf66100fc278724aff07af8e315d8b52246cbb482e93396907c2d0bae1560ba9f5a8760a4d3e558d6b16e0e445205808536baaf8a47ff81ed989a0f5dbe9ad6357227f41e533532de82dca349e9772c6a599ff4e5bd6cd8170bc9502bf527da9e06ca927851ac31ed463c816e28c47273c051dda329edbb99805de9bad2d0780487c78dbb571e85232ddf559c5bce7e0f5aa6214abdac4253ca5f1d792efcf8e3a65a16a1ddb870004ab37c550f4e5302bf33209e4ca256e778ec1cbe9399efd4dd63f1a30321eda457171415ae72754b7ca939f044c3085e42a43e7f91909685f504c755670f827956778536018cff1e7529a9a76396264b548185bb2a3b508d8e3537c0ccc688186f5e24dd388d8589769641261f2cfb50dafe82ec47c03cd3f3e576ffacc7f456968e34df752819870db267dc0c0feffdccec1cb24e1508bc1ba4f7ac08da62bb88eb1b8b01868bb01837a66ffc8ba83ee5f179b8086234e962bd0ea2b346af95ce37949c0d2c942e8d8bbae9cd7b0f90408eee34801114c5fd09efc839f2d2810b859d7b15046f858b2b0d7b02ce98d2aaa4e671d209d444f6dbdb7510981f54ab3827b194675e7cf95a7e95d5282ee97430020a899b7a8d82fc7657dac379bac745c75b0cab226a1742c42640187e8ab404e2e076d4d6269a5c36046c901615824a84e684c6acdd6c3ba8dbe75133733958c4db68bd8f7961935c62afb8bd649ca0c8aebd4f8642278e8f167ef34f6559a7b571a0bb114389423994607d6a16c5f794af514cde83de29d183318f80e061b3c7d24214d289aae6722b9fc7cbeff608151b6e391ce192d10dedf3ee9309e55a2880092cef96ce376483d0c45fefa7df6a5b3c1273e61f34bc89001119a5fdaa430bef99bd3bd8d9d5500d86f0dbe03f0de87a917355018e953502a59bc8c7771d3268d5ebf51ecd93a033a950d6d26f60bc86abba871536b3f88bc1b7ec5d71570eef2b10a5d65aa9510312d71f7cb096f98257ef81faf31731d95ab65a08f75af3c57efabd2a15dff995f66eb1d52d59d0e12e6eba766ee85547f729a121c90bedf36672003e5b69967ad536dd75dce3dd3476af1258d4e8d87a61bb23af6a4af13c1439ab014140d1c772378b4ceb572abfeaebdf1800c5c94afa7163df7278e38ef4fd10f9aa900c015a848a8647d3c39963cfdee88616274dce681f38ca3ef78651a6487eeb188e75f2f0cfd05875b2168496a585f47ed484944d77acf85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h15dbe24844abe96f4ea3d7392f7c10d2b498040e1ad6880d1f12d62e641583a27764acafcb0b70858da115bc3208d555a3d9d39311b35901c7f03b1a1cfd7a286315cacfe50cc8fcd425a93659700710a76c16e5c5e0d9103baf55d976744fc94d585cfa103305958fd5f97cc78e38264d765e2b0afde77307f74d7627bcad64767410f07e72ce8f452364673dbcb975594370115123def9f15fec04f33acfa32abcc5f005be35a6a3f52d3b5de1ab1bcae142ea37b8eef70ca1dbf663bfd021b8821b8222942b786c7bfa86a49f0ca445df4d49b426a61cf71d81c21e856dc288b9d532abb2e2911c5e646d74da3e90c1b47abb3dde6dd1e34f63b365a3bf162fae4d136a5093c1ce46dbc59e935d9873d594802f057fbdaa24e1b536150127d2ecb7bb349ce0e8d1878d4386a0726f7248132d6a65cd68703f755934b659d3028730f4b1d2528816e7d767f7b5312c4dd96d1d33fe1646f04faaa164a1ecceca43b380d4f50b6271c5ae9bd4d2d5d6f0c4173f7514a29d8d1aa732ad2854ce589ea2416d614ae453506473f026f35b806969fe23caa6a8ed2ccbc9f47c35cd91fed92b3c301eef635ec6e116ede28660dc07a67841340c429cf30163f86f1947963e5a2edc2f0a8647bdb7a7a7bcc3526d0474915d05a18f4601f9e76724dcb1f969c957e0eaaf80bf981916e50fca42695acd80d1848b713e8cb332b9dad152e1d8fc7421ea24d892435f564ef1cc552e014ca6df76d15ff28f3ae4c023aafc2688c5196b1b1546288ca380b81d9851326c200a3fb038d08e12ea3495df2375444ea6b154bb74cc49c8011c79b020ae65d5daa225ea7b357bef09345d9f89a73577d7aca35b383022f15e00e019f5d3b68ad9112ba5d41434d276888169b5095d85149d7613fb42a3a9ca63945571e052ad7af1ae5737216294f63ca5834ccbe0eb53ce70c583407f58ed6dd7c511759b570e93eef83f69d19e8e88f9d7414f986cf3e946cb576d42c7f5676c4a5e522cb88cbd462bcf35c0bcb52866905eae6e432d61612dfb8361c4fa77cdc48580197b3dae5c082aca7e7082baf0d4f86d96c6807ed8eaabdc3a9ab303a082e6db014a594a217b8210611358e1bfd975b55a5d6be0d13195ac38fc0e2d95139477a0b58fd6ef4df284f5845a6ff7397669eb3a688da3a4b87aa5d0651530a79830c8f23f03573e69a1fb8ed37ed540150ac3a0e7de0fe33fff65549e8f8c7e7f6e15d5f782d8f21f97b812854da3eedc47eedb6270b22b17d3c862ad3b5b7d4a47681e2d593b1d39abd251507a0697ace6e88615a6d0a55f23a6ba4f7fd081186dc13f72c021e0bbbf5365c2bf8710005cee6bd108795a210b83e7d4f3ff0430bc894ebbc81410314413f1730aea2c020c602d6bbebaebd13d9f5ac64a2de1a9aacd0231edd7f59be8d4b720944d08134af82cb374dbad8676e82ac3569d0d0054d03a3ec41ed2549c31be1f94edf617da7b82da82ae172ee0e31d8c82a7aecc664f20c19c3992f58bacca06d414eb6fba1fc0001bcfc6b768fc4dd347376f3c6ad5f9160ea24fe78e5dec91490aee4911c60647be20dae2f22026ab5db6df3edb4b4df2965668092ef32b5a3f4efa4bada199138366f88320bf00dfc4718de4f2128d2e58510c9744c4edd9a5e17c4bbdafab4d120dc8a826e1c60334319963978b666a4c6a333adc799b6083ae63b97fe2d56d30a48bcbdaf40285acf366db456494228d90d7cc9ef6207f7f5bd3cca8b70a4ec5b335e4cabc2bbfadd78c5be764b493b13be333a28e9d5bda766b365e5836b46507c3bc480f6a2e5ea52af1355d39fc5b4d695ef036a3a1c34218c7ab9213f012c5b2265452a540dec740975d8fd228672e20f6fe5c06c41ef9e1c38543b028d1ce1a83647960acb1ccba43a2220bec57324e8ad7c38ab52dfb2d05378fe9599e52c3cb0810efbbc3197b305335ce796ebc49112354d0480753aec497b93371b64bc3a689fdbf6d25bd9ceb2da0544433496b8defe92ecea7a5d524e24f0efa773fc03807aab38f1dc5e1e313be54cfc3d6aba2a775a0729d0a9f9488dc136c039535c3d25d9e2a1fe5cd0524ffb27b297d63bf24ad450df6a682e40aefcc85a9d5f30d63b59db373b2fb6cf539a334dec980d9fff7a53db424b097448ec0c7ba102a84754858905b4af7e1ea9d26cf12e9a36938463633df5e0edde5441a832443a88c200f2f356ae8ab48c8fb4271f9a3ccd15ea563bed47f7e2d91446f0bd0ed3aa23085b97c4441057b706845e8190c5fc68b6138cb94b80121952a3a15e993156225b576fa6d9d7fc86feb1318416f44e033473462bbd30f65c515e4a539d165c47ca1e97a3af0a7f1a4db1ea0439496bcc56ed3c97f246f0c96e173ea40997f0c7a1deb7f7b93f8b42e635c1d581489a51dc6fde1c122593e59806157674ba58a241f1965870d603aef51c5d84a4020aadb46a2b05284fd2712e022f8b9d1ad5b96da86f9ee550fb5d3ce9b90c04e1e8127cf8bf1ac2345fad0222bf3bb9be25cd397af848c2398bf81bb5db28f37a920e0c6e61be893de534b39c249abdb56aaf3923796f3c33fae956ce0adeca8d17e3caed563ecd960a2e6438e64bf2b935ed586a5317e32315933b144403d7911cf13ba35d30278a53bab0722f4b8febfd7142be452c135d0d5b47420f71199069eb7abc90dd73fe384b35d12a5f6826d4b760b029ff8ccdb30d8df66d5f766272c153adc76a742df98e228797fc260a3a9b533443d48a52faf4e6db7a17d6b7a4f2373a7c3cae0b49ac7e4a31540c7418988d56d56373eb8833b24dc1abc3a34c369171079e3baff422108fd2a3072cc06caea742b1d0568b565813cc1987f21585ae59c7412fed8f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2635986651591785f4e0af23bcdc3a0236ca5783174ef7bebbc32a6fce3f6aeac9eff1a2f06867318af4ee3ad49c62a698455e751a0f1a6b8fd1589e448b908d8e5d1d88a2b97d0cc1d99958ff7b0a45f98ea1179e22aa2af6be3c730529d894ae05989adb6e5c31e352f6f9382f7652dfbe10ee56f909bf3491c04d61a2e6207999cd41489d59d838add34b8eef342e2284d840a780c7d8c0cbb1b84976d62acd6e6ae2d875413048685ff8d8f087d824a2856ac40f64ba40bff7c89c454e8903b22f5d63d26ccfbe69470aad8d0173c553a3a95483419296fbe5df90584aa428aa73ff9ea7dfa8396e20b103efcda0279de02b0de20e3ee72499394e8d6d6b4e4b636f389158084caa8d94f9cfbdad9b597be99fc350bb8e71fac6312d40eb86612aa75924377e59cb4de3eea08c8869826d3a2a51b151b4713da50706cf6173a3ea539819ae30cacb7a2c0fec98230493bdd423dd423345b1ef620b0f8937f48d48458abfa13608c42e449570e56b1d4fea3d028cc033defb31fd079cca8cda8e3ee91d14fef0f1ba15d8887f3dc24d910ab245a94e1a8c51fffa3eb3a1fa4518097af0ff3f973a8939cfbc58efb38d22682ba82c2df6382f479aa8e2774e840df117cffbfba6b831c2f1c6869b0eb1cd94d5b9aaff31eb4b1905133ab94f60d968ce3d511908d09b131d843e8db1fd1273bca52af4aca57393fbef1ba3ecb0722f2e51fb84e69e57a11e2050f65517159a053b29a81c1cb4de8328519822e40d5df895fd2e583c2d36bbc56020515fb243ef2ccb31c2818c3817e91c6c88b82fa08d50a030d266846979fa8093ec41dbb433e7df370a27d9cb06593f751e120d03442dfe7931b99c9bf432b35cf85898b7ce1dd53c3a844c05f5acf4bf0b5ef36f53a794f2793b7b26ef25ac7c54b78dfc170c126978437bdc23f09187765fea759a56c8240899931332ea9897597355cc0e1db1b77fc44531735e833378d9cd26288b322b24e41d67e8acb026baca9c99b7ff355b0d7b7c2d7a821f28580801bad77434a496f0a8bd355fe2bfcbb2cc78e0debceef70ab3ca04cb79a6c1792ad284b63d08f51d6aa4e0662b63d46070d46f85cc083037e0f6facae6623e39abc9f32d5b90e10d1cdac69481f0f7848e06af3d8356afbbc62fd28c940461d23139054ed1a89f1fc5326c8df8d38ec23c0cd5aeaf8c58d655c1f4ffc31502f6ccffaa22b84467fe472506391cf3966d2b907812bec5fa1c755f31e487f17e049f5062782819b06615dc6a9a3382ebe323fc99956d64f343be610d941ff5686762c80ff981d90071e95406b9a860ad8dbd491a2f1192c3d1777a7668300e66f2e23b023b5ad06aed4d5fb660bc0bcbcc4f537332427f20c92c9c660782a7ea40ead5b16ab7d7d6f7747fc37805289b7e80b5f5b27d50a95c34f22af07ceb325f3803a925d88a73bfd8ddc91950688857e73c30bbabc944fc931586e18e939fea0e6a27ada69f26a225eb05a03cc0baf5bb79409a4742172c5787d1e834d019c8e1d9195e5e25a6efa3f2595edc3c17c37852f23bc146153de418ca13b5fe864222b3f166855574d8c03343dd980d07e9bb32c740ab74ed15f4f27e5c0508234995302e5afdae08c5b90edb599acc54094e3684c2f81c0f2aefae16af45252f0cf2405a2b05c1771efd3a58e21e5c9e0511afd7b5f1d416d8950c26ea087d3653c5076845a42800485edfe715e0c5d1859e3d3f46608cb95a0e8bca32e4d8a6145a664e7b05f89cb7b5fc2542cdc7de532b21a481021614b80fd3babf8dd6d76acd5c412dc17b99d4a7190ce1605cfba35caef1349473321d29ef6e04c61bb6bb2077e484f7b22915ac6cfcfc7bfc6c13f639a15ddf2c3583cc5cb9d4622437529e4f290bf8593af715064ce9dab5beaf28889e6ac1a7fac5a90798d80941768b3ac12d3214d9fd116af67ee05365cf8aa61ccb2f8cdd6567526d02952733ab8086893c262bac77548b0586485ae306cbadcfc3dc05f667862a4b81d69e14ebb3b85968db5a862e9f78ee878220c00a92a3bba384fc4bc2e0d25a5ceb971c76b196406b8a210420aa352914ce14f8afc09577a3208315b45ba099302a813847fd78578df23fb9a736f4ef37aef31d228f2ea0c3744898efb8f01a50873da0447b655e28b4adf757722cb1b71bc045f0c05a5c009ee6ce7b6aa51bc3a4ae6fb2b064ba4dc9a45f9d2cf35899aef2d70c22e8345139e242c3a3861b57e3c06f6e6e732e015666114c926b4c2dd040876795c48b3c46feac99a443d88c1bb675f6b64d2289dba9f4e01de78f0f0c183072b4a348f5e8578b203fbdcc3090e5f06f936cfb5021e7bb034adcc5e894b658ba78a942a5273e50ef3ddf7c2f503365fce984fd1e20e12db7ad7a36643b951d062463ae71c37e2bb7de7e6bfb939df52043209f86593c5573261f129bcc758e4773ab1929a756a95f19cc6bb71cf4bd0e279aab1b54e62ce0133ea8dc2558f2ea6e3f8808e85976da4e4af2d3afcf0a553a6eeea0f3ee418250520b096959485eabe43aad134bbadcd5e9daa0d695d9189648619712a32cf0fc7841e02d62ad3fa8636d79577c135dd7d7a2b84fbcdd70b941b3934abf26458b9821002bb6e15650500c7a9c449ae1167d3d2d7510eba3ffb5130fe7b7cc03c11d7ea4163987e7bfcdc02bf1f33ff82cb4e37014b430039e0e9c3e943dda55aadb0ba69b31d216d1a62c483321ce483c63d9b2f4b59e8de68f4a0b8d66aac5d188258d0357d58834dec24399d42ba66c61dd2a1164c62dd6fac971de723c1eedf900c9b605a0b003043902bccf251299f310d0af4331b5ab28f6ecafe3ed96700e6f9b9bb3d8ab0a395614b59a91e51b79086ead8f8151;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf209f8b817e93db45321bb73805224a06d4466bd8adff1c206ec47cbc55fb02f9f59d38dd8af22baaa04bad4ec282406578abdc6736dd368c3c9b230ed2cd666ad2eb3b538a7e9909b04519da32ecaa6bb3d3bca19a6d84618fb8b4bdc42a05e88ea938364bdefde80526490e0142c26269c38718a605da55b38a4fed9f2746b93201baeb6c131a93207fe056a421466cf1c2de8840ff59749a2741279bfb04f7feb8bae7cd84774eeb4514e45b3ad79a759b57de5a1c514b5db79099a6adb79a470f1a6c946360ad328386f9e0316d13953965fea24b3da1f4d79029c872fe06252260285977dc60d9fbee3f31fdbc74c6684eb3a9e972fadadc4d15b173c82a290963f2109709f4d0c040208886049f475244c9162e9f233ca3aa6fb697be257a8d90be4b7e5d9f021bdc9913b25a04417396201e53e15d18b1c54e487006d445f84a539bc805cfdc799ef3c2ccd128a7301e30f691fa12fd805ceded72466e185b3bb11e16aebb3fc39bc0c5bb2dbe772074ef3222da62e7392320e9c009bf0331467e0adec15b17eb451394a80050b29f5580426f469b670886b01dfa8802726873c9078eebc80a37920910aeeeb0e18a6519e0c6308630e7168fbf78858f10b386216b5c9feaea3e34f0e7fddbad6ffceef2133c0118b1481a9a2a863904dea819905021d8c19de3f10576d62b9fd48dce2d765173d94a85a0c9f4d090a2debb94dcab106ad6cc0a845a07d4ff5ee3db4dfad41d8f8228f829b8897c3b2c3d5b1835b197246904c776c927b7c4ff2905e14ea45b5d43c7ca36578ee5a918a850f6df923418f9e26eca1e06294d27b6e78cb17991f5d80f70e7a3e6b01366086065d93b3fdf954134e1325e42f172b45196323cfb52ea4febb1990cca2f26373b766ed3b5c2c156b1ce00e82bd87bf500eb2ba19a8be2286eb9c3d2eaeb9ba6135458a5c8d1042cb5f6b5723741629c499095ba9048a39611e9e1bb6bc94f016746b8bb8878490129257390f55bf2ee839a8b4c1ddd19ba53e59ffca5ddcfc96c8c020090e60b4c17c0af969f47ae4165f163979f075f57c41947874ed74155384b9e2d16b7a890888af46c3afecf2c1b6ff42de305c063b8d1a9241af4a56647a0a0bc1a6f9dcbcf8a1257bb77c3c280f41cf1457884ca1e692e1572a8b66fa89c350546e8c8d22d2bc82351d1ac552a3a063050b908590a750d6167289b7d286d839f4672f1f8b768c8294cef7650b9b6b1a14128df7cff592230629aa2904966b1d5d960832e0250a2253baaebbf99131c28788526bc0bc499741975f0d3f3d6b06a09009ac549457da20cecc30701d209eebb5a21f57086c9bbbc4a6b9cdecde025a25b42700ebb4ea5b3190ac131b9a05cce3da19924223b4a1c2f09225aee01aa097aa497d7105748f95269d942b6d68f00b67e7b6c82cb47bc260b01523802751eeb44c5b68f29c74902095ab2464b0b15a3c7a93dfd7c66cf908c0b9f409d7c416a5ccd1d5de46cfb16234871f554ca94caaad56c805fb4a92ff7f37301e31b303da96bdbfdf464cfebce770a3de0abcc92a2a7fd7dc1c26498097fc22e328f83a96227c7e0fd18fbcd59d27d96fcab8e6c3ade256488385ca83bcd349cc5f203ec6c2732415b086a5ab192ca43eecfdd20def67c9b5ec903a0084b145be08ac8dc7ccba7fb541e1d4bc95a021fb3f19fd117108086619228679cbb9f8824a995a8d35d381acd79f17987ee67a8a0c54c0a1f57a0a3bdddbbeeb7fa328692a94a68d153a1f724711099e348979b5199ae9fa8c586089967d2ed56b56583f747938346d700243ae8ecced7b5bbc658fdc27d718f591faff1cefddcbe83bf2ae040292b6ef912f16c1ae50f7a83020870f4ee07c7acc5240bdf3d528a268490365f2895c9d0056eb74096bcacb0091f2650966ab0bb88b94201098867236f5859a06c7b6a625eae57a4801d9b1bd008c206a57c9a8b0231c2ea170f4e40e224dd0729876fbc0030f553a8bb592876a1d340e7b1c6de6339e891578ca82d5ff78383691c1522146516d97d1238964ee5faf062992d514cd0c3686ded2cea2b8d93159788d8b815fc225257cd195b93dbb78f8e4bd84d56931a11cb118c603e2f9e60634bace0c8426a0655b54ca63d6cc8e069b0aff3211ad36fb7b952e0c78c7ce97ff77f3b36ab691b2cf6c66b89607a17f26225cd589c798756cba999557f0dc9f96598c09168fd98d800fa6b4a88fafaba67e5c2618bab8d273f95ad547e29331828ef9299f4366c698f4d8dd7bff22705f2f79a11f39eda9927638a1a11e9155df7f2006e9d23c93d891e10806c9613b86c86303f33c32ccebfd8746bc220d6429810b01a8370af9fe00fabfccbb283fae84b7b9c406ccef842a4c3113161c9f43ebf23aa110b60f5dd74245c9547044bf045773c3b208771226e7045a1873e91c63c561d3d3175958115241286c4fde07a6c1bbb5d2543b2fd3ca1a3983560ccedd4296b80af6dd141858c9f941347ec759b3facde65c13c9f6f19737fb5a20e9e3d63b10c4ea9249e4ea63268b0c2349adedd5691f1002529ed81f067cdd2ab4cb8ac19bec87305eef2118aa2e8dec4fe98372a2296f4fa071708a955e65a74aae856f34279c2ac5425b034b24673808f9207e0bebbfae7e7acfb4e8e5340a73827cf7747f9abacbc231be04d5616942367cfedae3c8c5a618483d74e139c4efa7b0329c2701868308cdb96075321e509754674f6fa24fb5228b99ab06236edc5b71572ed71d41b2ed9be2b3a74950e8caca6db4f1d553717170295edaff761ceeb6bc824fa4194250682b628cd3bc3e552a08b2d178fc6d917044650835c474768f25a456f95241d81f227e28ecd2f65da82a931f1cc97d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9fac780e58ded6544406238c9b1085a3b8066b2bbd021e3177b4759baaae152510325b4c3fa8684722d229461b37e22ee0b28a509371051323f5ad38a0c07651d453fb95269b4915eb441ad7cff1cbb982a04d7a4808db5aafd3e2e8a691a90416c29ebda9b4c057a888e0b923e877280bff3a2d716c3dacc90bd099f9aa9123126bf5939402487c7d646c9ce4bc49e79adca7ba0627694bf47f6297a85d3647649e9bf264f16269d9d17cb294997bd5f57401c7c0fff0b531a329606094929cdefd4f8d28db70918f017f5e97e8a49f65c0230145a39b077d7958cf658c2784cfbb1d25294f9f00d09a554007902d7446562f117787ff7b71df6651a504011c700b6ece20705709b6031f6606a8bea2cc3c2a7c0f92866fdde6be481202ee0a821a0fd951e81fb604023dbd2dd58385cf5cc11cd9c4b94144b609f3729f37d9ae0e45dc4b03a37d45cdbddc5ddf889979302070d6daba610c0eb91cfa0f7a208bf7c2e8a8b5c957d2f48952add5fa1b5f0bb8c42c96a2db7fbbbd7c7f9109d5d6071581a84c04976fdce66e515c13f8cb56c8e7e807b6e2db4440aa6a57a93ac7ae6409677807d3cfc1f511aea3ad0cdca2c581e35fa9cbf5c03093856b66d0f41b4afab25462832371beb8a263836fc267742621454e8849cac957fdb1587f957439c8f9250c8836009ce38010573e8c990b65709327efcdf6eab55f1498bc6f8e0435fdd04f0e338f2d9560c5526f48a55e2fe880ba4a820b87e27670ad02b7ad8132ec2476af8a4c08349e6d5d6c2d271f93ff2474f7dba00c163c30142d1e3b100cd55b15a0729babdfe605b082a7ec125d1a3520ddf184868cad5cd74086094e3f0ccf266dc4227e9db18ef908ee77d44b6dbcfc037c7df3f0f0388b14cdb64b3486c4d1477c1a794d123a239cd9147793a252c87ee495239dd2767cddffe73a6f21a42e4cd4053b15704b4b5391c28a4db4de9bfe2a48bcb0833011bc2daa243b513d8b025393f0973ab9dbe015a4f3b3f961e22dabe6f007e0ddde8e2dc1086c8850ea87d546211b574e4e08e531a1c5ff528dafaeda8960e2279181f1f563f0064fedf310b1646953e0fc81f9e24f375fd29ad4cfb87a3fe94ac20a79acc8b023c69a22984c05b0569e064b6d93da4e63d286480dfc49382a411edfa1cbc21e390a77b95d249a639719d6b353fa8e873c00bd61e7ccfdf58f006c30c6446574cadaf8279cd20cf75bde7ea2724ebe5bcecc23d16a8c02462e12100176c3829737525ee160c2c4677d46e9e8d63bf2b67c0ba79fce2442079e134a54020922e83e75ce43e090d6c433915b122235d3743470a816c305eb4464111b4261080ff5635da0ca8c4bd5011bc36b2b2c1bc899a544fd8c5e2680c546f55895ec5e393a0a748d6089313338babca9f7c6226eb90a90804dfed3076fef9c574a27ef902482f80a74ca2cfe69df338c78fc95588c8d15b76681496bf058e26fe88c53f87afec38279c9607adc4ea1e2d785e82130d882bb9168efcd02eab2ce7d7ad301c0c77df18e12fc05a825f4e495552ae984e8f908b495ad4f3f351402200f19ff7aea0fe1687fa4ee1298cac16e7e9373c7e18581a9e8f500ae9b8debcb416ce2e7e18682b206d0b8d9e6caf29d6a1524ec6b44c0c96214adb87a5ebd443eb25ad9aa416b61e6e5e64a19fe8978194be0409fd039fbf1912f254cffd0a0e44a5b32d3e6eea75ad63f5741c2508a5719a58fde72d7cc17d6427c1728a289a5146cbcd782ae51611f8118997d2500f554ba0bc7b0ff0ab5050e6b561ebcc661c1661fd06073267685ddbfe5845a75d012a66f851ca9a0644027b351d53ef4afe5a958b7782fdf485e8919c1432ba838ea72b12a83d0d7940fc38e24be1ab10efc2443fc620ee68a616f167dc961b73f90fcce0c0626b952b00234ccf6da92d1177248f47d681d70a36ecb17079301075b3ed9048bd31a37407a7a28d92d54f427bea998546f0afd52a868c18be428e3b5a9b345ef0d5263b7ddeb0f1823fa2a664ef03368c33cd21128479d324d3f547adb544864c5ca75556fa3d752116a83d88e8aaaffc30c75147a094e782cbc2d9181ada02d8cb9690aedb84cf539206a320a02d8904dce6910595b7d3b39c3ffaf7a3c4a8043af13fe40771b5f22f4f1c0ca7d29bb72bb374e75098636a935594d4cba0bf072d7bf14e28ce4f37c9b96800e54404747280bacbb60fcad7195d092e04c9169b9892f076cd4dbd08781cec66ca306b7945583d297bb10cd59fa7812b9b118566d1a87fd74ff0da2aaff14f8fd0edad25579b8dd7097205c3e7418198707e3e56f336e0b7eaf7905710c83ab41f3366ea9c4bff66a5ecf706f4334f5584cd7c97cc8e2ee5c17530242aa085ff681590f01cb1e6df319b588994b69a409345d35ef6eb269b42b9d1e333a768bcefa5dc5e2bdca0b3403a805712b89768e83366f9944aaf2d6952b822c9f19be96296a3ad658277199755be00d776720bfd44f2c7c8ce28a20bedd31bb87dc215fd32f226548915fe0839bd0543c8fd728f45884164f4757df0debf6df7466ccd575f191fc3bffdb4050e0ab366d32ce66ec5a318b980df40f1b31b4e3756108f027fb61aca29c4e743ab4739e86952127e18e65a8c7ce0a17af23f168fd93a1391ab69b3b2456b7c0d730c763c12cd3fc6d2502cb12a0586b88e8d8fc47007623b18b9b78724324514c4216d82fff27032a33bbabc9742b896d0f724d6213224751fc32334bfebdf4ab73346feefb3f1f2a1478cefa9f5e2e8707523d4574336f4dd02be1414ad645f1b55d83f4821b854cf6b544e3a22d422c9b9bfdaadfc3b20f71c8b368b0a7adabb948f9e1703c10686d79be54373326493e421109;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha6ab2ed36ff1d51e0589828a141eeaf00292531e009a2b534017923e0ff8b82677b56fef9a782d1b1f5fea432d72e76166e24ba5d36442209c6f3b1b92f40858b446af1a01cc0d6a65af56f33c2de36834fe10459c1c2da9d0112a7c02a47bc0c5c30249980f51b72a50f27bfecba3ef3c019053eaaf3592c7bc479c7ee5e6469d0ff97be6b3407624352403cf7186ba8630b1e310e05d9c1e9a3a75588e03ab678c7b6aa2dea0487fec7e37847b4738e11ec56dc524eaa5a8fbe454b37a5e593b196e553a334cb44ea97ae93d874d896b84b7ebfc3ee1f3ce0a0d871ad804f12798481ce3b1919e0c8b90640b09c00829b60764863acb60ea0c13099fcb97bc0b81d6fce6383f2728b9a8ecd513ca78a365d5ca1a86a3bda8bf902a2ef8cfe9819d31f143c3cd7938cc6264178ede62a7f57dc70b065575187d21f12c3b02a4d472ff405f6120511e9f420e6421bacd46c847be9217687dc8813720485efb9ea3b19277296e5a6d24437ee9968bf5ec7d232abd8a3f34ed19083ca817cc8e4528e628b789a3450767ccd9c95b8197e7f8fb94d17fa38780b5c62c0150edc53bf2251922732a77672b8b2a2752bb5b9a12857d44d5ab6190e41adaebb580a70d0e6a5eceb26625a90b49464bbb7974468c5d21514888d734acc54ff08bf99297dd59596463e9a32edace21b877432fd5a59a67c0a78007875b402be8705c8f5aaadfd603cb006a86a506389d4fa499a561745c772f163b4a83fd9c4009d2a8a1a95cc1491571472b827b3d0731f6f77069eb0bd491fedb3377089e8c89f23da22f3784fd08cf33f120fe9966e3887ba34e5ac107488139af9466d0750c4bfe00500d9206ef09753a6b063cdf87d246e2eae00d8cf257c1927870c6573e08764853be50fc9ae49101fe5d81132176fefbadcd685b775c69510b1ca26b591d175d4383e792d64d338a5c8771a52414217658993b4168935e6cd5671b53b46f557037293c079416085aae4b568b0f72acf38dff73bef7dbe17106fd3b801a910e1e19fb11cf547992be26f7ac54948588c9ac05601938fc775a75b78412243ca1510b87dfdd1af96f048fcd119a2808434b1f32cdd9ea714a11831b09afd16a5e8fe98e0645bf91040a5206725ef7260902548f3498d3d8f077fde52004214369ce78bb721149d8f37e0b7da07db3ba17b7c525d74f72e83da69fe5799340cf7d460931f8d22f8b4eacd5e266c3ab74888e82ee1adfd2ea4033c19dbe0fa95d9d4b9825a17140d78566351df1a2772144805ea41a0e64be89708b6befa67d9c5ba6f06c9f558f4edb3e3ff1d6418a648100e473309911cae2ec42c875af2f05bce46c301ae89d719fbde6c00d39d3a07f4e03703639689f2fd4fb0e23548efcf3fe6321a2c91e8f6b113d8c2cbf6466a190ea6a30e19a17c90faab2f9a231448f91f5ee92f9734401068ab76604e2a8c66d9db93b64654f0a55e3212055a05ecacdc390cd01dd80aba91698970670daefc04480175d28484409884e5653da277c605d940bb553988daeb5957554507c9b3bed4b6667fdf45e5229a80d79b8d6559319e78f8cb37a92f958315cbe46ecf11d8610bcd6108d702eee5d1646fb2c6481969f14a9c0c5b6ac3bbb20cdfa526c5005a443781bfac7d4d0b675f7a4dfcf94feab2191dcb6178ce7f0fb98b53eb96f572ee21767b6647d40f0ab34290191965b57384c82781e3d046e6d4c07caaf45b94f5817515ebf78a3bc651a24060b26c556e098d7b97989d015d31c97c43a8b9b7d1ec5d6c93de6743345a2e6f28011a1569b88dc39a5f19a2d1a2a5ec4f49547d2cd7c339220e85965222acf9c4254be95e67e3e1aaac3f4425829fc25ac685d8427342f07cd7f264027acfd0603858254a04c9bada462b33163599b98bbc9ec53abefbb4c195006551fd78f44af35922843c93464c64415ecb9556abdf8938b465bed1e82991e123ca3e512d80560aeba06fb5bdb4f3b69934e6557d990897149d4b7e1e76fbedfaa91a169b5818ed401e7a2b02d34bbbdf22fceeceeca83d5119ba7a0c51dfe99cbc7c18376e4c9e08cd0c3a39fe87153ba520410b003b148a5c9b4d8ce3e45da118569630694a1dc8fac7604140ffd352ec7c19f54b9c8cc41e04941dc825e1a39ef3ca5ecce445cfdba0e9f533a739d50814f0765c2162f21d258f8bb52108bec0035d5e6131a6c3bb435e142d71b6419a1d927dd8be6a2d4505e930c9119c45e7918c51f381d3bdcb95879ecbe80b7b7f9620b3daa8b5275421f16f82cf915e036b74033b0729eca222b76ed80f0ea0d5b357c53ea32b60d7a43f9bc1935c70eb5dae529c16b78679476cf79886147104214a7c8d867f6cc254f8fe7fdc9c80c03e5ee3c48a2577479ad9738318a4670ca28a84aa0f968eac7fcecb8234d15f6e5674bff8a2b233b382003bddcf48dd81c1b4879a7344465d4f1c549c04e4440911fac12288dbf3f7a59848bdbf46095fdaaf67bd0914b43c29ebf8f600162d89ba5d72203aba26a78a6c11a80ab27f36e1b18bb73509ae20aedd056a60e2eed378c51680bf30b613ca56dd3e71df9b4d139769744ee92e6e143396c80e9eb95a6341cd2af007b46d66687296fd9fcfc6d064af8400f83c28669d5d47d65c652ee3470e3f90a11aacb3ce6b9b9160106a31d230b11c05206652de63f00273a0e7d30669758360140e623ce75973656bd7c0f18292d735510374c597c18c8c909749cd72a4b663d394b5957740d2dd58bfc286c4e34c2da7acf504ee77d973cf0b9bf7dda880d8d7cff429e6ca4f036b9db4982c33e2487e70260865c23e0f989cd251b958674af7122af1a3cb4a8346e66683f4f90c2cd6db326264e2bdb404b3768c013641a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfc04183399e79fe4b7b8eb603ec45c6fa6f52a2d0f5ed6d7eeea44083d09af395d98a62dc04041a7eb4200ca3f0618409c4b5f27bcae1df47f62c1dc89a712700ae270fe02f89088b3103244d1ac71ca08f29b2cdbf21a35f39dbb935bb075fa2f7d88158afb9b1b242b1428d60cc326502217892dd0d9c9b282c34363cfcf67a85d75aa7faa92c9667b7535609bc184301ba27b74d408e1135385accb3eedc2b396e92743a74d679d4324815c8a0a6b0bfee133219a8261361e2d6acfbf418d1de62c066e6414e6c24cde3e516a0ee0f42407ee6ab79b286def7930941e1cfc6eaeddfbb50811ee1d67e10a598992e2f7c94f3fc8ae49b42cdf0ed726732f5cb7ce08f73a77369d986f440ea033b2a01bfcb2d5cf84a805295e46bc5882387bcf414b93a5a595a6687d4271b6db0ac4d63a2047c15b623f8e182f70ad4b8f2dc2c31b7e88cc200c1929e3374080ca3a8cbc16f72db6135c917d7dd7c73be8ea4c25ebe6541e96cde2995e368395d880b04b4796f7d6bb9a0a2547d13fa05c70f9228a96bbb675ce9fdfeefc0ef51e0d1d361ea4f3f6551a5839c32fd91551aa860e8531cc9f50f9d0ecdc7d03c2bfaaae8c06be49773bbebfad9f894be1a0e8d841a3a7c5897bda47666b1d9a762f2df96cc89f4228ccb3e6312688c2b3e23425e44b14ef80d7a9af8292a56a02b5d7aba0334fee4356f6d14757f5db39f489c435401696e9fd7853918c59fed56856ede009b41e43f50dc29a570ca9e35f19a426d9eab00557215841fbb26ee6cfa307a07312d7dd5943e5e2920026c58701e75252f73a4fe6a3cceed14611f4f4c9c65cc93ef9adb1de83bcbd3b349477180e04ac95f74b23b93b01342541d261b986c84c5345c35bf98d527e196900f82c73c54285f8f5a5835850827f1a94ea266795ceeb45ac6216a5c8b4dd964f2811634c5bb37863e0df827a4dc80a30013c24205d8cd800313e9a541ce2941522a540fab47b1311d01854dd645f94cfa57cdd35595d3fc4b12949100cb25facda5652bc1105188d6f55fe4a637bd5673b4c7ba2afeb6e7f5c3db2452b91ddfceba44af7d8b67f9bb7ab39a3f37b7946faf54f28c57628fca8d8e3091d2ab9e7ebd097c58dc16b7ec8df85da668305a58f8ad9e0389f711e465194291b6b62567cca52ee22274b9d4ceaf5eea4656bbd95787dfd3318d6337aa8392ce8dd8b1d4d94627317489f2296397f9f42e3ad38ff06c01a36e6e55f23af056fdd5adbc7f21a1b53d8d5a8ba1173ab432160eb9035600d14c6ae9b1a9be213711f9a0cf273e93e538691891a181e2d308c3c205dce35168c94600ab0832fd7725ffe41fc030f1d968df8ec44ebc6593408a71d44278b82e78869406f088815e0a833985b17a14b94bf43fbe04650d2da4e27e3cc68a68d9ddae899fa0b5354f97f60b7b1e4e1e0172337a58e27d78a8bdb90f8b871b4293b284b6bd1288ec10c0180dad0a425058f901e9c751e24a982f423e7830add6a74fd1a0ceb37e025288f7f70b8e96db63904cb47fcb2c162e820d2d52b9799d10a775884c01c1d720431e7fd862e8de7c5eaa7e18e66f536d92f8e89ae4824f9c2c6d18e5262fe26b32a60eeb40e6bdefa64d865c8f3e10fa2970c84b793ac591d7ffbb2d2870749e7ebba1cc8bc9d085172ee4c8e32a172bcdd772ff7162878930a36feb3751378f7929fdd5e7d63780be29f559b2d55eda10facd3e7ae48e122ae91d1c2a7da490dc54d5d4283fc03b04c39494b0b9053a5a1826d3a0f55691cb9a7e20a9cc8aa263e9bdbb57bc65aa59a63de8eaee6bec3cb61425883ff94f2ab503d4d5d87bfb6d790d1d8d44e8cbd232463d23f5623f3efd480a6332ef0e841571c3b37876fd657888916bf0ccbb97ee42851be4405bb5c338f32bc06159d0418a358cdae87e196215f66d3663935fb99859fa43940866a1f0ee6fa6a1a7ed8f6df425bfbbe36e5ecc64789a8bfea825982dd86910e19970e485434c0d6cd8aea652f2d4df567ae8a2f37f64c54f8abf0bd949fb4e840894811d96ad77e5b3cd6a6e3395aeb47741217ccc6ae2e643b29349e4aebc204297441fa535a0bfddb2f225408e0c4399a9145b743d0f7350992f3b5faf58d6d442cd52cc61837a8566c454dd94d4f8fe943a503f0b84d6b5da81898b05c07fd351788ed832620cbfbf1aeac85a825ed2c152f515c821db97a81c87db92302f45468295bfb36a6745640a606dd6df6e99d900956df08a63f77624aa5e7be3acd471c53f272114d4a2f62b75b85b9083f91070d32d28d984c80a9a651e763893612ac2e948f2ba9ad6dc505c9fe4664940f20fcf423457748186045c8cdd5028186b354adc2a4924c34b5dfa659f67710eef133470ccf24d6f149c0a06aab162c293c96bb236d84330e966377b3c7b7323cdcb551613605ba084502d9a65a5035e1786c14a84e946f6e803f574f2c98e47d11d0565b2b28ffa8c032d8712d60c0b52c999d8f4a1590c08c751425256e1b396593bf7cd34ce26d79102f2029721ec3fa947ce100408a041ddaf2bc69704ed293492ce06370a5865a540b0fb0c2a3ce3523331e68fa34aeeee8fb2b666fdf18724719d79265db64eb394615ed186a77b570e09d908d5d86eb6bfe67ff8c12fe785a39e157d4f692d1f45f6d6eadce35ae5d260c430def3bab46057f88ebe4caf41398d1b013013d3113a4744f3f25d8aaecb9494c1d1fbbb0fec78af396257a917799f15f14a471ddbade62b3ec78b0345d8e06a899cb9432ad724df538bf066ef7299f8828e981e76e240050026e948c5063a5043f6fb2ba0c3f54f6ff615a1840d624e201b4582e8492848ae193475ee04acba398ad534c6a3283e96772a1bfa31ecc80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'haf95ff682545e775785b4c095e488b0af09d7a9ed5465c2f1c3390bf488b955ef007100c7d11508f3c5d02d7455b210552208008f87e10d2770abd6f01f2084b498fa716ba2f325aa4f5b83d03ed85a19ebd4e93f23e2d379361cef3c7d1a964a6c9d9441f40c65ce70f88e23cb435cedfbbf6eeac33f5a000eeef44c14065269dfa81ff3bc5995c5d70ff169313dd1e6ab051cbb1246a87a78e375a0c4270cf107d17c2271f4e558fee36b750149098fb365f4c0a3b14d2befa285ab18711520ac8b47e01ebb77ef9c565fc8b5076139bbf58f2c5824c3bae07df3aa6dfcfb758b878750ec6d17c1c469615b5e38e471410498de4804ae383f9638c49833c90881448b5815a8c6a0b123ea25ca1be5c07687d2e5b6354a1991c6f27ba529759092ef8d4d80716e253922d6f8444703bccb427b53e6799119d669dcc93f518e57cf842adfb96f1bc8bb9fb7332fbbec8dbd807d5383b89edbbf31b886e5ee4d20a4e175b0d985d8a25be95425a2206317338ab133b69240192fa5d1e42db2f5c7daf47b98115f46102111debf89294adf3370139cb2503ce0d4c1ebf45c6d090a9c459f94d99e36c8a53ca833bacee915fb8f3232a0d17bbf597bdb16ec69f4ad3ea34e760eb4773aed94f8b47634df0997e764809a610f1cff5fc5c195447ba05a6070c57ddc733c9c91322c1a76cb0f1a512349d776e5be98c4ec466b656082e64187b0768699ea439bac6f61252fb8928d7f0668283d441a9ad95b80999b437e538c0cd0f25c9051c0227e750ae26c41f9d741c11a655e23bb5f1867cab297db9636a26e393cecf655f1ce88afe65a42690fbba303594ac4b99291b98efa5fdccd63f5b80c6ec7d6a7450504399324303fa5f6bd9460ac1f50b26a0c40f9b696344493c586ad40e19c94c369813fb05429106652df644818a20d770f08f5f2fa6566ef7c00f799dcf1cd0efe9b2bc23dc3fe8c8aefdb0c3f4dbf7a52e28621801c5234aa8b93c7ccb046d1c19cb90926dfefd558b1dddf7c373edc07acc059ce05ffe1f7734ec05c2014987947be10bd017ddadd49a179ced7051278849ca14a6ade9e1cdc046f697a54fcd41bd9b09ca5544e8413a7d1f6aca997ec909e95a5f25f815e7cec413ce09974bdf7edb7e043be491f9d65b22f8d60378940516ccd4845cce9ba84a8552afc2e4b6fda130d78581a2d1b33ed73c8554a523674e304136e3ceb59e0ade46e19798af6cd40dc9154d0ad43f22e6fbb8378ff3813c50af1de8c27c3ec88f4099ff372b19f6660effe6c8a132653aaa1b6ebf12b056025cd478318cd1b27db9da4ede8b0064a7537e1aa4a63c9f62b16e9ba25291f6ae802706ad261bbe5108f3465a8d7b04374d14a8003498096b4496235fe56a924abb256e26a8cbe7abf29b2bd0f34ad66f3918b234ccdca3e63b23b4b246a689e12b5d227ac5217aca1629e01ba5a9d492268d35bf844fb3c08a31e04a6a158362db0b225bba7c43f804120dafbc03d8a25a7f5a985cf4984ffcf5de090232baa7fc834c8cac4a7f43d488c21c7d3b7ca65af6a40e30ea3baeea0a6b2ae706513e05d1122bb454518e9354132c1f624b1d8ce6a67e6722641e014a1c74f2329eeb3bf19c2d5f962e00c660de2df6947f86ffb31afdde607322bbabfdb18165690bf5b163930f0be21e31006436d9c5d2ae51f5a0b02baa9d80ca4d6a6d2339e438d4efbe30d05ba9112af303ee4570cb0a36b77915bfcc7e8b8575f1fee794d3db11ea75e3fd9e9c45f673c2b46d076edd641668b27268a9d0ba98de71f700531d66277ab1694b49d21cf6afb4a9d288f6fbee7525d32a550c5f27d8fa270a72b4234b4dd97e5109a7dbd3cc4680e1aa38593d756a42d52406b9e56cee73e59ae1a95f7677bd73022f48eb1c6b6001cc6d4f6be69e4559a535a939ac13f6687bc955460f6327ed5dc5e5b24d775dc791fb861446ddcc66a8b933aef04b192323b6be5a715b8a7a64d3ae7b4f0a072cf2e405d1b447e21777a7f2ee617cc8dd7d2a5cb40ef8dbb6e81ed0388b77f0dbe95358020e9e8d1b90fc1569eab6ccb8c822fab485f339d9ff8c8503089392f84f4d180cf6a33750582cfae5232602d522620240d54cd8c40603a3b95fec229a65087b4a53ed8f30dedff09f4b4c20a67649126f2fb301f0d1a145a116875dc4d50ef3b956361e22afd194e36ee634adef9b7c0c7918db638ef4140cf94a70d5614f2d85fd79cf4cb259c195fd5d2368029fb2ec90668786bb7340b0850476f791301c19bb03f0bed973aba1f573b260b1c850e3ab74628adbb4ddc8354ec1c757fb5019f216868165e0b4c721641dcd8bd2885e6aa468f0f926b93450d490a67c89f5f252be9a990b2e5a3584d7bc1cf2833ce1ba367f9ff0f3f80bf04aa08bc0badf865c23bee3e87c175a01cd3960175a271f28ddf9157aca796b081c0bbee2d40360b9b15254272342f1be43bdaa3a38c5a44f43e6fe5460a0ca44b835558017f2010e20d7abbf03b631430d1f7ba5d7c1b56d061312b21c4e3dd7d454f2e1ad451be24659d87509b00d319e541a1e31e2335024ae34d9771579a2da3fb885b47d4a18beb9b02d74a1bdc12658bb8e9703185f5ab3e2a6bdae5d95ef396a186f2c0e29e73fc0da3c156d789bce00859dac6c0cc983c037e0b3dec4275b76762136a1c97f4215a9df35050fd0aaefb3a11a46c615090b91adc711984c7ac1d75d0e3c6616102ab951d43ce7739431aa457fccd685ed6d18425d2af4021756573bdcc044fd5469ff805aef2d83a1b95f3f310563354ba730eedbeac3ceb14c4f70abe5828018f68191555f8ba79454a3b27b70e7b4c8708b73c367d9a225e8646ed66e6b1cab42e3bb0ecf113b540573;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he2c9cafde6f310dca1caff97683b78537ffe90d035546d5827b61af098e06319ef232af1bbee0dafc9f497fc4c9e34f9459ed0e4af13f2c2981a97c768850c5585fb99be107545f92184e622ceec5e7b685b97b1669448d7c1a9ee1dc4bc1acf23b9c88ea21e4e1281819968bf42db00a00c7ba3fcc38bbd8eba1eb61e589d4f723363c91221a41f2d57fffe97f0e33e8487befef859fd603ebe5396546cc9862a2b7f9da9a5f03dd6a218d051600f511b2c7f288876d4bbae99fc9534ae1263480fe90d6f4f2cf648af9057e97c55e4826683a9ddfe451a806f6ae7d7598d68c401e0280e85fffee01c1fa44339ce95da8061fc43b2821f532fcc7046724c9635fc0f4040ab8c2714ce84117ea0b179a168e9ac64346c492f40c45ebd7f175f91e993d8accf635267d8ef9144dedec08517b7e3fe4dbc17bb85d760e8c6831185e1228db2960de55a7cf7c320043d337d15782ac1064d4c64dae149f4a68dec333de1bc1afcd9636d536fa8fe33fd26e595e539ba9e9a79369002e0494390bc3a256f12155e66b5678fed38841660b239062be132f1aac85b31f3a13f96ded7858115a72e4e0f8ba377bd98ea43f8ff2f15b24e434f82b6588460c8e0c80d638a2cce065d65fba999dadfe4fc17f72c75f4d21f68917ed0499a706767b566df595aa9477ff2297d780184c2f5246a5bdf376b298369eba24676eacb95a8e5cafc40c47e5d7a8bb9dd07a97dfa29669647829a4b18a84ccc389ea1cb428fc00377b73d77e4078e95ea173aade21ad5f8699de1694fc0e4791a3e9482ad9501ce980ab3d5623fe9c36a69a306565ab3a9671f49075950d527363f438fec8b06d26b60de934bb07c38a373b15c6deec16fe4492cacc3ccca531c16a33822bbd14a2ebcac49bb6e577964c3b33073cd4f4c80c60e2aabf2ac75d2714d95e44c76b94919fc033e35e4f9d006770c06914c8868b241dab30ea9316ff2df6c9c8b118933c782be019dfc508da29169f72f00740f9ec815b150fdcccbcafd60ccbe4a44a76aedd0e58c2952267ee3f8675abe6434ea0fd0fedc5de25e07f4e6332056fc3b4e0be179905e566c1e66bd6dc9ff1cbf7aef713033f865f9a2c5936deb43ca9121dbf4045c94cfd93598f2b928cbad3acb3c92c2b1900dbf206d2ffbf8069ce4eaaac4db542d286534764adabb8cfa380c5d65df23b47926e3a103bf4632585b1cdbfd6c3269ad8e5953f658498585d035a0b4a51fffcbd34ac2c8cf7cddab5f15525485ba606ec10c2bb83d00dd2ca7cb8b665da2e5c38e5b4b66e79f2996d67ff3866cc405e7f61880a2becb911bf7a2b2c2ba2164327a79e122ebe9ea987ce9a959a3d73b5a46ede2ccfe44b4c2bb0ad4fd9fceb8c18a4b6a70f9c8df7869520159d2ee29d8c6cd9f208dbdb5793cd00ab3a06767cd33aa86b6cb8a38f2a13fabbbaa4bfd7388f3c94469d1de4ea9df3772b00fb2e35b6600a03706353cac626ec49a735adc17e545a1a5faa9b45703cbf54f771b032b9978e98b4b2e3493bd5c58fb50cc2127fa5081e73cfee5d1557825c30fecbe45383c944f28651f08ad4a2060b4da339ea409509669f9a84a8ddf8d6bab87034d66014f3e858dec4b2d151bb89c88d3fd649417fd7c08650c33229c9039f93462ab86301b4dea032b7fbc506805213c3fca6b241618e523788bd9c704542fd834f937111262be62550b6f8d8f75b88871db702edb50135d74421444c4bdb413665228b51f84947b2fe4a1517e7554b01b9f0f5469fd34247ecc7f82f2ada820c1575a61d4f9b6d096e22e70301cfd788b9e7059fb463d540b4a0069b1d5fb5a1dc8f23306ef93993ebc3fd4995abfa83633a4b23453655e139b7334b8313af0c9cdba46b9582817fa70c10f4f3dc3f90dcd6d296446a0511e0c0a13f1f0c486bfe1007390b84ad27289ff48d1a3c952706b07078229313095a538a159e92a46bd6b97a951d3e200264afdc06a363bbc8e995114e9ca828e79b986b85d34a6a2bf5f72705137ad642702697c64f193e47e215763b4dca21d1420a1a0c56d0fda14f86d6f223e2be3cdc4964442a75e1a84f7075e554ed4506cb2ab6c2f6458f108526b0eee871f93fdb546c086bb56706015015c0f4262b3df113edc70ab6960321f3fcc6bdfcd06de45f4ea7092e2ff445b753c046afdac928cacb5fd7bccc73b13e9980dc499f8cd01c67124aa533a3494aedd80575fb11a6386d135cd70bed46c7a694106bdac2c05be1c8625c4bbc01fc512dee07a39ae817d8f7f5ec9b666a943a0a39b1fead549ebcbb1a3f6a112c21359685cae3d8946f6a40fd155dc864f79f1ba5502c2a883b547ca1033f9fff8a3415fbd7071ea2717a4b6bbb558fe0b602b38d01036e84f3f5771bb1526939afc9ee5f7294908cd1ade49348ba3ddae397dfa5ae560f00fe191e886041ee24c0fabdb29cf4c366c91f1f45f6ac12a43678dc13a0a3c2e351f6d9ad9e261173fe196214d9387c7cdc5effa5619de6bbc3a1a8b2e47ef1d27a940fd362826714d2db4a0967a1cb17083df8ccdce463d72a64fe72edab85d1dad661bd60e5662aabac12245b022c343ec8ce871fcdc5c4ae338daeae0438df4956423ce3e9545e4687f8b72aca8f47aef03c5c05921986aba8af67e89721e13334f8ec9470361472e95b3a1c42223e3457cdce5c2a60790b3543778af4f1db20ef21132b17c88929aed974c1490cd59d2cabbe76215d4feba945b1a66dec78b1cde8cd4569450b540938c27e1d208b838bffb6b67e8dd3d455413829e87e048cc739fb815ce70b40d1cf10a1d6efe25ca4373b103e6ab922786831b0c9c154ebe66fc0422674332ecc42c909d235ac6861e61f6df1ee5a83b84382d7392;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdd0958234c8ec63be66f86dc2c383631c9bdb900b294eac4fba662c78d06ffdbf90e0c72370337d8e47dff22c68fe38885ce606ac838702991214f2922ef1b2eb1c5808444e9d3f4a166c93743f65f1f46c2840d4ca59e5ffee1e68d337d106a20968333fd026c660809cbd2ffdbfbc4a5e94ccb4a4f308c12bed9c33c83849af0b97330ef2f842b7ac91d28645c8b714b113a2a83198ced50b2d24d8f597475085b7e2f53763caab50ea8a3a7203481b11ab03f8a8c17124f3c47d90b3d63dff699dcb732c29a1fe8ebc0b197e5330caef39971f6f7d7a56b30357f009ca0333ce68367e134409c3b1d6ee6f6c7b16d9f2ac89769f40e75a118e93d554d901d883242a48f2ad68d76deb8f0b60ac7989c24aab484e6c19caf8fa55272cc13a5947012ec1ecb0cdcd966ee7bdbc2192a2b68327fa7a1d655b148d774076735b56b60ea8f689497e8b3b6ab779823ebefc444e6fd76e94e8dec684ebf7313c3d58b1902eda50697a87460b1598f01261a016f22f8fc4089b2af52b2a7c5f847b4b7b2e357437726b7c2cddfe534871257711e9f5f15cf419f01117424eb3f521c2069cb47becac01795e33adb0dc6b1d02ffa20183968014aead4adecbac3e46e0227c860b2b74020379edd4d721c81d7e35fd0d52415a3965d2f7005ba41d3890a4940bcfa88a4e87665cc8a71b51c8ea8639644186c60be11f29b4a1f72d332dfe67fd9acd09653303a131873c6dee3987ba5ee401ff3a24ef3a91f1b5e5f0f1e841376b53be28212482c655e718940abbc839f52051c6599e329e0ccec94c233d30b11ef68a69c9dcde7d58eb76b620c1cf05f6b1549f9748c954dfd9515331873a256466c991cd8ec62fb067ed6c0ed7031e73e5c6b6c877317b6a79736a8a25fc5a935126edc6f239f9caebedf07d7bb59cb26f4e270a5635ea62cfdcdcf603a61a26893387abe06cb646e0b029d731bcdf244a4042352c1430340c7f3a4e2086b25559bac5deb906de8252cefee2c61efe42c93effe541b737d55a68b9f3e5e657bf6e51ef96a3ba08fb3df50547c83699a7687645578dd7bf230d8a3e3051094b2fe27b8b0d596292e9fc3954c612a1c55b3e86462ca3264c58cd5fbb9b28fa90ecb2435cd7389114f867a5da571a6328ffa17036d5f7d2661c54091e601b512028e7c00c9e9c551a28aa57d829f428e5867b335ec71b0cbbc924ead25ff6b0033889a5784cf28b23f13d5a86772e4286a0f14130bfa3e518c5890271e676bdd58115fe3163e054afacb9219df6f3c42e3efaabea32841d538389c6a998cc3be454097ae0ea0aefdf2adef1d537d8588f51455830822b5c0d42d642fa69cffb7c8e7e7f9c33c1a9ce647fcea76a1d888cb1745ab224e3e6a97b0affcfa99862587c56d08331d9e49b8498b681f1dbb9f45a059c8309750b371f6f27fe1b0ad4697e3657d7b1a92bb7d22e06f33b7d3d21590f3b916fd8d836c598683c4a9d64d357e0427461daedd96841e966847ef22f82568a247607d5d8d3e778a736dc9d3be4e53134dfe1741011165db471af0996149b22d126e2956954ac51e8e66596f8b54ad6f29fc924da4c102b24e1b95b54e3feb1f2bdd55f6876758f4042fdc2491c26118193e89fcf670615ee9e64584973c130d5bf7d6467130ba6974348059d65066edbcfc70409eea5995231c331765658403336a3a7699e0da6730769010bc43a3588ce9143eadd999a2a41a53035fa2365332034fcb684c403f7f422671d005ea11a84389c8cb4fd62cb3a7e8a2d2e3ac9d7b60a2ac9cde2f0f7f3aeb3a4099986912cf5518288736fcd71b065439a32b2445212c2fe9bb9a2d024c009de4fd2183b98dfaa2567988677c32f2a0d7ddedc8822ea12472fcc31f0010be3cd002dfe854d3d7b6ae96fed8e9faa365163b7f0b0b36742fd5998afe7bd672a095e30f664f7da245d82d4b8cc923989320baf693a33360a8f2d6cc47c1765b55d8a75d32df7ef73349e0ebb806fbcb4a162aa7adc3a282648d6366fa18fbd69de4ffafb7c809b87320a7612edfd32040f9954e6cadea690b477f7042db3f507dd56ef96d83e569dfdfae7259858f3d9498493a5241b9046bd77983a9ae1d51eceeff330c9e1127e538235a6b4fa7415a7ca82ebbef44e0a363387f6391efecfd2b994cab269998fe86ca24c8b3f929e5ad7718026131f96d3339794c33219b0beb220e01fe25d04bb19c10f4ddf19202f1951af999fa74428f1d63fb1f1af880425653fee78abd5ee90870786e665e270609de361579a08c1ca94ad47aa0267390d5b99a5a285bcd70b0f1ec43019f477c95bdd5c18f0475ce27edbe8f5780ec611f69e1c84eea9cbbd0dfa058f18eecc6625f406c141937c2347234a005efb1080bad6256236afda5f1684bacd50f20708145681f03f3a0661feb2630d4ba8a76aafabb3f87de448467779702859c30c1e0313a2b5bcc61699598e3a544de58eadfba36484f659a49e5a8ffd20a78d8e3ac99b7a5e10a7a255952996a4c56adb06ad9923e07ac1164436e4cbd3d1dd226f5406e08b6bb24c17a9125fb300c026f9e3176673bf9039c959273454d274514d2875da00b598f0b28b2cdbe8575a5b8ededb5888fbad05187b37c9a2b25140553327c9a43bb117c27ddda977dc19815ce5847c111d0bc7187227391a883d8a11abf3543c54552a1990d45e01194502078e779adde631a67f776025ea63add66c61388f2b8163abed3ca4003f24a847b0216c88393362173883ca118b7d187021b67b99049c8f3ce2704860eae1868d8180719fa55260e0ed8ec09d312819944e092f80616729120274604adb105918dee7861ff8e1342e9e409222a288bea0a65631ccfdd013f4b40515cfa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8125f108907a9509144796b38d327a45a33fcc989384a95edf2ba87a60c0b1c377aebc8895fbde355c4f04449502c20f17d055021de22de1ba5d36f70910b2c0ee4b895feeeaf2687ab699a64552c6efdaf6a2d8f2a811bde8209fb815d72dc8e8cb0bd5847d602c17ac9e5dca7a415e8f8cd02ea2b54d031251f8f2f7ab750f8c363365192d72a8c4514912956ddf66cc16bc056788336c60a195e35b31f293973ac8b036e7b76e695e83490705f5624b4142c01996aca330d00819e440eeaa9af808df5acefdb998498662b983192148867ba3a238ec97b6192468962d7b8eedfe0410f2efc87c3e474892b57c09d22ed11b7806d96d37d2cdb6bc8fce9ce7e34790d071555b52dd1daa7782b4b9c95c6a907c4907fa54dba55ca865e6f701f00a6b42236e7e3bc7e926af4bb4b8f506463a81492f9a3ad0886aa7a16b95d440328951add2026207a90c9a7ef88f2ff0c2e14eacd76b903a1d9ca401af542641aa41460d18c15a5d9c513081e61ef555ae05f3018830a1a271746c31cc1c8c0fb887531e64f25ac131d0fe8b977ba4593ca28bd69c285fba18a1e3aa0e841dc57472572160d5dd99651ae8912fc77552ca846f831330758d2ae440e33730bc78cb92667b836cc9ce8d66c5b74db49d91c6ff71818cc46815cad11e1242c71f3f864c48291adf9ab2d21950a10af418e02827212d9d7bd38b48614b3717684df02adf6aa9c74a2949703bca9749959044100a31e834eeabfcf5fc49645550fba0d675a64fcfbcf66e404ae3e40df4e050424b84d472ff0071f2cc5f0fd236e9c00922a4174aaf2671330402e7c944b59c271277ac18279666b448b64653f116a09ad189b5e90d8d51e8255bc46c1af8be3ec63f474d14653ef62ae40b5b10661def83aa30bbbf5a889cf8660228354069db0300b482ffd28295d31438e21d4eb8922242ea61cfe8e8737e51034958e7d20a86443c243be14342562b7abbeb6f37bb855df0f76fac5f2cb6e686ded1f4049ec582f71dcecb1d734fada7a3eeac0845819075d9e77bb202608fa2991f252639d1d2827a9fe382601eb10e2f1c74f327658ffc1da6a29d917e343864d3353e9abf88e1cc51c626519342bfed905aa7270d673d2ded04b50fdee88d124dfc1a2661c922dbe4210d07fb2d8d769134dce9c1d4f0ab3f6c380bfb92f01acd3f65fa40a6cacb76bd4b022e7aa67db16a2807bee494dec885b84d6dfa6a0dbb346510b6b37962993ce8286694539c117ad1de245ceccb4d67c8524273c873dcb1ad439fe1a45193cb2345339740a761e27e3b5dd0a47e422e921b89b5afe868be5a6aa254e6a557209abb490dc98eeedc7a58acbe7ec3ccfee688667d155db581bc92b50157dfbeecdcde12b6dfbb3cc93220915f0a891aea1c49973d8670c5ea08ebceac8583a57d7e6cfabdc1c7ca07bf0565485f36365ac492c4b318ee20d623c8a6e40d8e749e1fb2e2f217b1433f13bf4e8f509bb4415ca617e89e88422230fde30a8e10ad766670a8bcbe1765f5704ca8ba06060c31578d39adb616551822961d49a29133cbf2398b4a35b2b3c481706358c447a7adb44c57b008a2fb383b95255a20f11ae986f0819e764b666cd703b00e1ff520680fdcf6e642c48ae0903402c98a68dfb9408f391a9ebbca4e528086a7989883198afcdf6377541021d36230c3f3faf2943f59b1277ee9d9eaca320c6c1fb21bfd788f6257f1f293ca94b10e90c5e3de3a1fc0edf4d5d3d6ef28a3bed371c27cd532e28df041a48f6822eed2a8305ac1d7417d6c5162d612f270eceb6c48516017b97dd8540c7b72fcb491a53cb725a8c5477bd9fd5ba84307e68ce30e23b46605aac2c767ef37b26630072d964472ea19011564634f539eb33e3038bd4ba30e024453f5cbfb16e5d03c8f29172bf09d5b98423cbe081fd233889bbf70afd84f4574b8390c8b9cc6dac1a62f23f19b6f31c8b319a39ee3063f9f7d11367e00279a2f088804385e350b458fabcdf45d14731ed98e201a1af90a36d8e494dd837c436bb998b902c0f0e6dc0c642ee3e5c4b0b5b924396de5a30be438736cf9dd0a8129181381b137a9b0a7b69777e242b880e11b8f509f77cd463a87a47dc8c7c49a3ec06927932f22a328a3294dde04b049139af7ef43e95c3d1d2cf5c320d1d42c1f47f0e69cb565b5015108579ee4fdd7d43a41a118738128dd474fac27eae0e5446395187fc1d0d9a0cba3d4145adf15cbda020bd87c48d05d44633ef2c0eb5e917d98ff2255144f4c829791f881d13e2acc6ef06def73742986911cd032e3fe48e0b4da379207ee1c589b365cb89993b6312f9d5dfc452b585933f1bf7e74cbca3ce190dff57d706da3ecce7a48d00738b1bb7b2ebf54bcefcf7dee3c0f92b9ff9e2510955ea8e4b3c134015c0f750d05135315edc0986473f3be48aed9de4e7b2b4f228cb277d10b03a0fce0826b4d795e409d677f88b9c6318ac7f6b2c1231f94cdde3f761520cf3d73c6c5560cce3d04b9872cd2791e45663a7b9d34c06f8874843cf0f8cf78f4b9022a2b75ae4cd9ce346f9e5c66cbcdd1a280fcfbc42770a59a084b9e84d43e152cf80a9285539bc4ebf3e7158c532b5b361bf2246f49ad1aecf6861f1c736a663927137eeea7b3f951ac3dc9eb648a9091e8f7929b176c009b1275e28ff9d03d982e1a1ea360fd5537f2f9669be8626a7ec4b7670bee4e1865c61383568e3d5ab4cb153ae999a29f9814f5f2b421533b7e7f45c68f4d9e7ab5c392cffcd12114d70c90d768e081dd88de7355aa511896281248f973c82b06a40a0340d9945f45186f397f75797e1889a8215849caa26297239f69f16407ca2c007e8d9d4151f21ab6d3288eeff23abc604bd3dc20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4e94c940b2684e1bf05852b7fe3433efc858f1b3693811b072926fa475a66c5f3114ef7e7bb6a04d1b469b32e7b040502b81e2fbd4faa5851fd9f2323948fc1bf6f767f92aa5ccd4fe7aaef48cb38f4c506de7fcdb89878d915fb8559fb4f608727c575f5662b0b341defc1b0ee81c91861488800759bf9bd20233831322c19b7ff8b6004e02149d06c2dc6483202e55c7de04d0a2c02d9a08225eabd10df725a127425bc3084c5fcb6dcff08c8b52626d0fdf0323fd7398cbf0f7c15fb64e655fad289c2da2d055650692ba2908fcf7f483cee0eb6ca5eac1ffd89b6f81f8e24ff9f612f4776449eba09960ab97e16f5c92adddb0a43beff334f6c9fd692fc7116f71673ed519bc308fd7a4763bca34d06b448848e64b6ed57ff98c6b1bc24872af4c3a3315cdf67331284d3f1df21525ec58397001300bad9a39d9e3394566ec3d9c8f81a35ba856c9b163bed60993e1073699ec1ffd05ff47d6cf363701942d8ce1323a1aa0822c37276f28989fd89da45218eaec11c05bbc4eb171c09ca1ec4fa71e1e00ee82afe83a6c0d82e22309a67680cdbaa14907083cbeac8755932dfc39aab545b19bf5d639c35fcfa38f8b02bf3a614e9a9265f51592e878c17621a1fcafb4f0180c0a888118f4d687fb7626ebfc061069d6ca6ab5a1344b608b4f74fffa559b415533a2b5c324e1141fae2ac8ef33ff1225de10af05899b486b3b9240000eb405ab0ec58a6e47cb57834acba20830b01cbbb840c29888a975981d7a475f2ee2fde7fd45d0f493cf0a934c41d0e286b21bbdba75635f45560dcac66121bc2b15537db598b9d1e5f625d4f2597763235e4566f3bcb44f2b6810adc0e875e837559ae29d83ab577633ba6f7f4349191326bfe6b1e2c0e8c7fec4193102191a79c46f898c2c376a428b066601167b3d49238029a7c329bfd02e43bc2e70a259d5ed3a15a188b96042e1981e597025b693a630f0ad8eb858597fba897985b842346ce2cd47d6cf7e1b8d35d6887d557c4dec04879421fca733a49a17e9c05209c80fb32f96aa33f6e2b425470342fae32eb0511356be4ed0b9525317ae7bf73acc1702f75c2b85ea0f17fe26e3f3335df153cc47b0a24d86ced0481b1e926cf81008d476614d7b1b1b40c3fddb53721c0e2980cbc2b433951107aec27769998bf0962b6481582bf2d92ad3de52cc4276e8c335b5aafb9a218ece7fdd29b15157fbe894a718194a50329df9e64636f3ae4e38c60b950dea09225c2ce296a60d49866f2fce1fd64b977bf1e71c8b6df8221192b9ef24e24147144735870bfd9426d8c368b05597e3df0ad747f17dd1549a6235ecfae62f8a9056519e7d2416365acd97a1f45c3ca555fcf0d5bd6711d83476dfa56da45bf41365354ea8fada92311440f9c8507853615fa435da65bcb47a254b8f37a92b56ea1f70faa06392cdd1b11bb4c63bacabb687e9c8d5747e65cc0e20abc6f18d8fcd4b136f0d8ef83cbea4f4b2a1523ff5a1dcaec43dfce193640f641eacea8d13117febab6a25a13f3ebe69f27fdb65800af642640b28b37449d8eabea055f86771e8ef949b25972978ccdd0ae8459372d6e1af681f6854c23382b549df060cb9f8e52210d70e984073b47f5ab1cddcd4d757a58a21a718956f860be7d54163ff232d5397594a61032e16a9a26b68ac7a23a5a8c1c35875658ce8845a697745e90c6c2e4d8e1d2df0411a263851282c80140f80467d41cc6cc52b1e867cc84c44ee284e292ad116d5d12bebb273f8ee4bb88d6ce4a80fee3a6f9bc2640c5ef897ee6df3df18e0cb0815a33f13313d7a7c0441e0bc0a8c03ab7692ddf7d65b1e27a781b81f06b68c7e1171c4aca8ca23cffdd28b34aaaa7c676f3054cb91d1f14f10118bb5656f0d041998adf5b694ff11ac17d2fafc691368faf4b79e42403e24ab16c6f237f8baa86a6cd09f5ee62c9cbd2c9d2b23973099da916229dc26c798074cd14a08f08d8712b6f4dedb096c0a1b25a26dd4153bb59e565e181529c4216e6d6f0487fd4bc22ea3baa034242f3abde62afe42a0e43235e3851926a4164e0895140760bb68ae39d1506f143ab52035aeb1d5d24d09aa41d1b7d097318045c238cd7acd1517978b7f3fc5e4cd1a4f8fb4cc5fee72f13c227251f8daa410b25d88b064c588dd1e913d2cac48dda0b9774085c0a2c4ce2cba809db31bb53e5153570c3c552108766474aebbdbad35a88d5deac114d7a64dd3bbbe0a26a25f466f19240032d4d6cced77b483803fb5ea581e0a2c794139eaaeef19836345c52187e4bf50844a2fa95633952261e3656d3f6211882126d00668430cbb153f12f8384ba4367d03b2f4e0e8d34786485510e3f0d123a801c813e1e8808fb0c550e6ffb5bc50bd9eea38bb02cd99c3cddbeff85849094c3ba2bed866d8bc43838f0995011d81628cc98fb36bba855672b8808d5e8c2c75a3b1de079a43235fb74a5187861aac861816c9f10c02a6da3175d3b5b5716fff3d05d6aad6d3c8bd6065e22c6480d828b4fea1e6b6e337f99559c8a8cd7da02c64aa7d459045cae2c2d27fa1c40ed91c98b6936cb120fa2d5f61f014b9b0492b8d7198c644aaa9f2fdd091e08fcd728c03497eb213a93d9daec6a97a823b1e9fd498a3fdeb3ddee8f1211b0df45319ce117fe40b99470f83af18b1912e7ed31a35ceef6da26653f782afcfc9a28aa4159ac118378fbbcad19737c39c90190058d1876c58ea757738fe7a714a630ee87aee360c7d7b88d6819601c9081090852ff49957379ce326785a82c36ac3637f46ce7bb5df66d20dbdd26666a4ab53d00f40e67a7f67642307661caa1008fdea016e0bc31dbe9d2c20aaeef0ac847b32948ede41bb7c8fddafa02abc78a05ae779;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3d64ab0cb04e1948ecfded1ffe86883728df32b56e0be3109d3c03ee79a9de3f52dbd47bd2dd8f9091895771d86c38bb978bced5b3688d6e509e33ee7f7d018cb827eab8a0b6e61ddb0725b2bbe98dd22f60b8f0926e3ffadf87b494369c203bc9a699687c684462183daa7a49125605a110365a748ddc61f8ec7efc7931dea2c100bcd527be52676c1e67b9c6f3bc94219b5eae5196bcf75f150fb695c70b66c30ff618dcbec7b47b20b2c3b3719dedb528664c8bfdd0b9f9e824d4486f11286461fdca006975d05c369f0bcfa1f2239914d50e0ab1e209e8dd1f4143366143fda8a0438ae7b6392553637297b3c4ea09b36ac850fa1c30cdadb4c89afac3bbd375b941d2a2ce90fff7fc27c26cc1f21d9fd619649d00ac61fc8bee494dd15145df47d0ae12ae859238cae0b59159117bace6d374c129987c13d5f7a1bd5558f801d800b9f495acc35dccae8503c3f02abb603d717f7517a003b0d23229c3cf3336ae26c1a859f04208ba19fcbcb7f3cdd5da76f5dcf7076809fa605d0b90cca2dd43dd18d23c8eebbc678a1ce320360257c3fd575ff45c9c736afe5c490f2acc98b3a39c63972f8b7fc6d245befa43bd32d91ef37ded9eac1471ac647f93711e7392e8c1b0a9c46daa6161f3c56080ad3aa71265b47cdf4cd7784c41729e40eeab67e12e53febd9a0aab5044425221548e69d26d8a410d678c1218ce35f69dc311e0ecb161f9d3524c1d3a74e8df0e49079045b24d5ab963db0a78145f59926dd258d4aac2b256563b52a76409806132324d0445e227411c228c36a918406f0e12ca897468c59b868d78865fde91babe679ca8213aab11b94ae7191a7851b0364a1f06251abcb190111e59c2f7c07f8788741e8254c224c814076ef7111cfee67b79a41dd7c01fbf65366da97b8b9aef7e4053f6424d201114cfd492733024aadc70b28a8899d6e97c487593c9fc55421b38a93b3b6ef746d605d654bb4b55454d54554e432da6f0c984501fb9755a709841676578c1c74df32ede1a7bee602d87b6b7f415c7a7db2445f403391aa4717f3fa66ecb2a3c6b7ee05f0a9f3e3269ab2df5bfc22c5a5d7b0de52a3d93b68f41c6328db3d80c23420bb333d3c9cce02de51731bcf028834edc948e8ba662f7d2e3a2b7415d097e7248056aec254be00ae4e67a851acbeca72d0e198ea6d98c9ddebd45aae323f1cfd40e996ff3c49edc225e721faa41c0035cf9bda951c474519657fef1cf3a987d943ce95144b3673995207bfd47bf78418bbb44f52adfe640297ffe74021ee4650d5e6050d882ed247a754b1da5555360216dc412de94b04665ba82c7d9385cfa4a0ea2a0f7ca2adc99190db5f91f17eb750dfeb26254fef065cac96d3f5a3df2aed7434532d67f0f9bdaf3364b65fea11fbff31b14ca66c750d9d00898371f8e0d4da1a988e6ade86508e680e41e77fee4591ec7880cc4f2613be1b01089705751e16f120a9762c7b637190ee68a32de48382acba0396aca0f9be738c3ac1ba611833e1eaf5a422469fee36e4c18a80f1d679d8144b3145f73ae297bdc75856fa46cea8d2ed1c9dabdf8a557b8d6118851d53390222a4b05f05a53607b5cc40e0e3239176ee0c84e02878065c6cfe92224489fd15a7c845ded8df6d2d0f6528a32e9a9ae9490bed917aec28a6042038eb51f150b23bbd30a12755c41244bf537c0ae3f74e9cb38e94ce788c36c530a0d8a622e99bdd97c083ffb397ce03dea63e91864a957802cb9111ef25069d686643215ba1900739abb3b2341490f2e288df7c565f4c4935f5dd6719c0055064eb8f08927832f16360c37f1cc349800f5a7b4ce595f6ca42dd0287c96bb87278d83fddaa8b7a26ed4d7b2b5ede91e2a96e27bb352f6840d618496892a78dcafe77a98325518e25e438ba630344b5b6952fa2fec2c03b9ed53d120ff9477bf588de666294a82825d2d8d43812f6f8c6cc516287d8a165ce0fbef427f599014a1d6d5e217646da1373043442fa1984ba0c3a73fd5617dd7f6952f266142c04b8f927945bf60cb0119b161460c6495098f00b0066a354b12a519fbd8d742cba8466304889a552d4a1699e7dd467b7e956996c14fbdfd1b7ed0f43ad64f518bf580a394ef254e42641a18b68837e2674d44cf0d3e865666f972d3f6ea47a043de55b023ab81694ba231ecb6020fa9f0bd634d5405237d177e29fd9527d8d0c679d2844f802f0d61419a0cf292510bb510c052c0053836a12d971679d09df2874d515f2874c1c3351536b8aa945a9bb8ea26bb6f8e38ab7e6c4e31b06b11faea8045bb04c59d974fc631ce98f30b9861b07e7a6587535f3104318e92bb7784e7f3786ec507003c8302d848643bb1af9d8a59b6909ff11a2083a5294696bfe15cfda60b05582d2aa924c19b07a75a3ad73271d7fc6c3b48c2632eb034b6a46dade071fea01c26a9c577f47c5a3507821b8772b9e66ebc8f6b6624f43c85ff00b6e4a27b295aa5d0d3716d2e562faec4becdc67fd8f83d62e71000d434458f49fa2fec84725d39afd243aca15e1d1d30b962e8eebeacc319445d7e1f2705ce21967db4c66d8c33e81d9d207fbfb23ee79c5670938d448f2c3d5dbf1b886e692492dad6b13d41a6da62006d89c2399c0393c1cb7e26b70ba0446647e886fd375b648e53740f8c0c6e253a9690a17c2764bb9a87fe186767b3b24496f60a571a98f72095e10259eff9fdf7829d8417c45c95637b1975f4408296c3eede0028933fa9fe5fb99a2481596df48c150d6275981b4f2706be6ef1f26ad2de95fc267a69a3b8cd38d89805781a5e9d2c0e44f4188553df56f892657cf00b4a4e612d3286aaea190ee69355b64d4c5af2a6dc61e4c88f5fe0ccacccda18b0b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdace698158dc1e15c6b67dd3cdcd7ec0fe858d51902c5edc346d2ad9e608e667d5616cb53a397ff7443f15ff1054f930a00d3a35f3ba01492751d51dcac4a4ba269b2b8621897d094fd8d4db1f9f76d50a92f1bf2efc18159effd6cb5c591e9bb1d253aacba9f440c0609c350ce42040d560af6da9549ffabc22b8f6373841dec0a2017a433d76d51b4665d944eb0e6d9489b2902aa75f438962bc12044592fca2eb00a6bf335382c4460627260800f33cbd57939fafad7fc5021d903ccd2a4a3b7953d13a49fc86a552bb609b233f798b27883fdd5a5886f6095d13c09b0854968855199bc887af6a23d3f4017bdc58d0079e9a663c9eef73e9c0168265b93cefe730e196118f196b8e89653ccd37ae2461d9d837deff98734e8c6d2d25a3f231bcc4eef82937f630a6447e13dad4513cda018259b3d2ad4476fbd6d2275cdef5eb0df5e9832cd942fda916ecbf9a69bf7dbfbc2ef8d650cbc0573abf6dd6fe4341f5bc4501e3ed1be4b4082f1f3787ac804e9323d747afb91cb67ddff1205f74d4834a853841d02e07f17f07a0cfb1647d9a13d20b751f584e3cf4e6db069daee40a845ec38c2d30e3e7cdd59cd12d9784e8e598cecbf774a9aef92223e8fe0388eaf7e28bc5ed7821437d0906654d58c1f13c3d4f21d7a73d00e4b980f43ec0635e3f85a4004984de16350371b695352ca770cde2f70f3c3a15d0ffada44f23c8a07bac9a700e232f0fed9fcef8597069820e35ad64fa11009c97c28fd7f5bc754b3ccc215e7e016e1dffb6de557524ab128787ee279f7abc2d0e9026cb7408c06f2ff0ac0603fd637290569003bb2c96c782a1eb8f7f44ca3ed2dda95894780e6ab45fc7f23d7aa4e01e8d9b00bded881f173fdc2ec560849e130554f44cb6e26367905181ed8fdbc29d83ef07178f04b694d8f6c4e7679589cb62cfd5ad660de592332883d2fe3cc5f6e1a59f46fd5b6163edc8067f615e80508bdca231bda302bbb5f0c6d5c6a2a2ac7948c2dca8782bc2311e7a17fee99988bf456f6f85292e16f6f115aadb921d675f9930ec3e184589f05920af97e9c5217c28db561d7f3e070050090cebc52addfd946d8b699f22a9aa9ef02399ab5b75a9d86d8639ba17e6e52c3e792bbfeb729c936629710325558c7512ae1fef60e6a08bf1fee76526d414c6109e6c8c0d87bcef4e881f93af7b0ccbe4bf8fabc5b8e8e968961725bd46b0762bb5ba4ff73414c4a8ab1df94457bc592adb51761bd46caab9ef1f3c4ea1e90455341312b1e9516a571efb9fd00c01248e0d22a2453d46f1c126d1fefcd3852c1c9f04bbd29fbf22409fc078dc797670dbc782fb8568d4df9481007458c439172051db1380147cb823f85c45a9e1b9830955063150b4f9f889bfa7f776eab17605d6d2b46dc9d8bacb826bfb46094cf4832c7be5b31f399f2e4840e252f388020d5d86d2678a85171defce8dd4bb7143cdb4b22074f3e96adbc95e93339d11ae65bfcc05bb4047acaae70a552acaf25692065aa573847e40745f5f9dc7d048111f861ab05d96c09ed59dca72c8e844779f7fc14b2e60bba59e313d37781bc8443350988efab895ede58ced4a000b8fd63b2cbaeef58ec2173d18764085717fc49c3f58dab157d2f7f5d750bf1d878c470f5f4ca9ed6f3b7d89bc55471b92993f862582522a7624066f13d7d12e6449b828dbb70fe8c2be466df3f608cae43c67c26a019a93d1c5d0db1d90ed80c440e6292839e79b8b51c48894af3a1219f989b09a8f9252d16c03734a6ae2f259730ee59a07915a3247158d5199d13f521e2b497b907fd14013cdfa004c622b117a63d9a2c6daca5f4af3ac5ffabf00d341fe52c7a09421de7e8a2dea2b5148c4c4811d00581f4a47baca08033a83ef622f9c93f68e285142814fed62588824304d0a0e9dcebfe6e8d7e96d2ab43512a3e2358b3a9905990def95f09543672250b83df1fe286bf76c0a56847786f1497feca618efea201d978291b3633db8ee6c18faf215dbccd15a2bf4e1bfcc375d6caf1858454e14c197ef4365d26b205a7d6eabf366f19716ece6a6a08dee2244d5221451e4c9579e500d2e1192e16509a4b6072225530075ca05262408586fea6dabf8a2d0d10d7129170fc891dbb7d3a5a2e343d04152b0ae15b53ca50728bcc4a7145bce1dd68a0e043d069c13acd255997ab1e7dba2c2c4092c903e5d65e0122fbd98b3b12981f99bd60e24cd22e73345aeee90bdbe4955cd064248edf6de24cc669722a2af95f5cdbd1cad6ae8c03163ef6d8db8ef087cbf79e7a3c75e0e9f95488f3fd0e0ebb2a7c474bae9929413d658b1a03bff4fc50450d35b9cd82aca63c698bd1845c15c3981282b61b9d05a2ce1c6b2355b01f3f08efec08efbed33355789bc53ca35fb0c0c6b8c7c488d5e7002f7ff631e3125647903126d5ce63468424e5c8d5a29c7616b7252614d00a4610751af29d5f5b8d588fbf76b4dfffcfccd7a9f72f76b9bd157fc7e04135e71902b419d3b90d0908cb9fd7148f552199037058c20be95c5bf182a6fc644b07fefd5fc2452ab26c5df8156aa001eb5986f7f5cbcbdb93fa5be4bd65cf190304174cf56ca4dc315626d04b031b140a591a585f328aea9ead3eb86b246a71ca0a7ca24882f24ef6d180b795dbe578d4782e6f1a5b2484b91ab51ca74e9b1438c94280797f21121ef0b641c0629269b436c6aca2423c03807b06e87e8002d905912122a0c344f422491dce96d443eacba41e19314f4d865257ed06a40d6e34b4215ecf31d57134aada60270f966b03e45e9eb472f30bf4d5363013133ca64542a6b528b9a590d26da2cf4652b713dcd8cd48b37506b0ac5743a1ea3bac53699f5a7d076c3f2eb1c9b5f15e0c5c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h20f83af98f0cd8a7930629d92801ae9a7426afb0bf541c00be86675a24cdf83db1938898b4cfc6dfa762cdccf29505147c1a7e080fe5f1d6a89b16d91a9dfc9b1e3f4fc5709edb9c8bc82eaa818523bea7ca833425c56dc017031c3516d3453d54822d6925b00ff1ce2556acf9d0e5ca62e6a0c46d7c287304b70668434efa888c758f18cd40d92e4b17d2377b884b9b3b1408c3c72f529a4d0322d5a9658a5bcd03841e5e840f80bd9598ad27b637be867b609fce0ce6172b9f5bcdfdb57c6c63b5c6803762a951ac8e8ad887904b9517c33310577cba891502c3f21434c4d1488968ae138a2ba97a26dd939a092cc14b72adf62689155faee4bc945eb2093f3428b18ab2f524faa10407a554a51cd5557c5ed65de92be74659956a793b6cf408358c454c3b98149cff3dfff79ae4b688e34dc98ee00ec49b990bf42854d5a55d16b164dddd23cbc66f8616da8035a14870d3e5175ae3579c47d03e114a3423b1fa4de34497a9e7a8bdea354ce2e01c583e38eddb642d2fb7ca47692d1b4e9c08f26f7730a30a84805c3d710a372d747bbb48ccb8a39ee89cd59dc1e2119ca002c1a65bc86ab9c6c35d04fcfc74db3c755dbd5bc691e3e7ece431b31949d61025f0f1a8fd582990266dd303df7e34e9f70e18e0868b388b9d69218598eb10c57032f6dec669b91e50f74da9e0957785f101caf9c96ab1774f3e6d1921979be81f9e8f87201b6c562db603205c1c513c86ea66b4023af9e32fdf1ad13c486e0c4ca4fcf31b236a3f100292911c8282c8960fd4b1b9d1056a2b678b7a919c4da9f50d819fc6b79befe2a094f1694aa96b66c0391491ac4baf964e1ee07b311db18ff6ce125a819fa93a2f795b476fb3a48aa91da164672392e6a35663eb6ca72d9d5b6fadaa0a235326910b1705665753564634acbac71ba22fbfc9e2ae6d64749b480d15e275dca7a68f8008dcdc718271f8a98b20109c06a817bc732f7d3f536d97e97f89bbe48526525f5156f2c9c1ea8929302510741116323b94549740a12c9cae9c23bab0de1dbab4ab952c571a060da94d1d5d1619a21af456a776107711ac33f0ef6002ae010885698e2ddc1f5b0d51273ff0822dc752612aa10d9a88eddf62b9df46fbca702f29cd9e25e7b8fe8b518bb74c35e3427d1623f92b080011879b570e3aee09b31d0a947ea95fc0b48fd16d5cba6a05bb2a1c9827762e1b6f157fa044ac7ff789842b81d4165097796c5d6f0febb41e65ec04c4889b1b6288b7fdd87631da867f3c7bf72ce8b4d40ae014678fe57eab69af319637316c8f4746508245483e664e4681944b5f4a7e8ae764b3b207830f9b4747f0f92ad10c596d0f10bd736a7ef48198e75ad56610795b7d3f50264c559fcd94f1d7945530277fbf727818cdf99aac43e37fdaab5d7102bcf65b1fe9b21408e0ce3e7d0579986ecc9fdade202de3af1dcb0a0bff1734f4edbd9fa7611db243b9b48390254f93a5bc3e230c838c4329020a704311f71237d6d30c6f834878dca3828fe9c529792d0ef2a5d1826de380f2b19693b45099ec9c3ead08b8169423148c75c6a3e4763a582e05222d59e883b6117f22a4d3031a8c8217061c935d2ccbcda54ad70482bd534cef51fbeaeeda8faaaae32eb2b84257b476a4252d744f297bd48c76288f9985f5bf58dec43228511893b2a07443f4163848fb0f1993a56c32265fe62ece6ccde296d60c60905679b93929998fbafc4d2d3f5670f4e8ae79a6d704a0675b6635e6f9736494c08e4c1007e0bb2aea57ddaf40dabce8dd388b73a57cb2335a3b19f7e6d4aae4fed27b3e6b80a1650e699cd8ba6208715a22af2fe053992da3b7b17db74493e3a572eab7d1e0753a6f3710472d1337a1c6f7be489ea922b5dd32020bc718f298d2d3e2196ce9a46add8c6187ea37486b9bfb6f3229a1c9d43e30b34edbeb0ad96ac5af25f84b6203305d485ed714f44e903c004557c846d3e13cf909d0f6d05115c3c1107e3e308465a9c06170b22c4d348f0c5bc5684c752b11d8423974294a768b572ff8a8356c7d48ad4cd9a1bffba9dbfb9b39d95fbf3f0f330b436d22c3e2da3d30d43bf3e86836dcd1a5b661d8cfd4e2229eebfcc88ad5fba4cd3cbfb07b198c4948a0ef3a2c7763546265045c948a17fea091e34f9405d6450a4919ff5c81d95fb0976a41e15955a0e2ad2a8a901c944c17d7909c4ad3ecb3c931907b92b4b4f3ae2b83d4912cf95409c945f2c5e6072c80fe2a0e0b24be3996b30f7f253825ee2ad02d3d2580d94cd47837eb4549fd48b65415f798043628cbdfe03bc777e3fe1be36d21477c129e7ffb3b9a1953bcb0f2497ce4148223e7d25bd4c7e41ac5ff431470d74104c5cf887d8507026fb03f2b0d493ca5a53c8537fe47f787773e979af0c90bfba7a5c02acaa3167cf72470b958c0eceb08531e649e73abf30202663f204895f9af38a60ebee0ef44953f3e1a5575b441028ed2b916f51a41244ddb3ae24f69e41f906a4fc34d67224d605daedfe5f7752ea38b48cf7fcd9b4654cc46b5a5311f670a82b82a1f1abd18f8e0724bd660537b161d0fa7359d51ccfb56a36727a04f0571d429276e1b4100dcf21fd11a11876ce2a44ac33fdcb7b5a45aacaf915b37883331268308c6e7e0fc771d89c70d6f27dbb6fb69bdd994011700cc1e6b77cd98c5b8ae35c1b5802eeda1877cece0ab647a2d61a5d0bf8ba3ed68c7989b2fb7b1ebade43156c2e30b91a77673df17079c5a3fde43b243ae20c0f10775e90fba981240ebe1cb8331dc4c0786e109d30581e653a5bf367ef8023567dc584b52dc3170f1f2e03ca7e5ce640b546640681a7a52c3e32f9ad9a26844da025a3620321681a720510f4046d136015a57d581;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h888ed8960f1d15b1ff211749c6493ef71e26ae33cd040a23f34479c635d1df3a59272bae6b9934f54687423c07047dece621930e39537ff8c3dabd65f0f58d46ccf0bb1db70eea6cad8b266c2e71367fee585ed34b18b4e94c620366bb0a1eff4959f30682aa37c6c9ddc77b906b491f5955ca12ecde716a0d8f4d7543eb48ce75a8d09aa3b93220125d17bb1782147bea148a08a67392edf636434cf86c83437e35e11472d96e185eb102a53d822f37babd413ad515fa008d68b3beb758ffc89e7f03452f750c0316b5eb4cd7bac71c81b9b8c66899937c8aef78a095d74148599297a9982db05278e5f86f9cd03568e9d24b8ca3acf0cae219b2feb5c2b730c692802aaaafe746482d98457b672086194ecba796f1b512005a0516ad10f4bd8f8bc7eef9bdddcacdd036f96475a5e6db29a7a89f68c2985c3699c77112b84f96cfdf025fd118685ebf3ca2ac218c74385eb553e99a34dbf81b163c866cadf1895d2180b8083fc742f2c8d2c2ceaee6b85812d998c9c67ea4326db5a5176eb519c0df39142489eae3d44c02f924f97b882e692ab28d9013f2bfe9c2e3b34471b439ed5c9d215e483af3b267537065297f8c6d11ab2c589e3b712a5e18aafd582df2f9034b7dd0c845bf9d474813eca980996df936ccea8d30ffc12abd142eae9f30a0fc01f949e004676556af938cfd4128d6e632d7cd9ccd5a9bd45877f7ac2c2820f1a2a2036cfe26706e78f671cdbfbafee42e0d835607851dfb52119fa4493dd23ab76ebce3cbf30f6217590c6ed6206fc5ad0815465a0563041bc750883a55ef5091c63d24f6301c9ba70661b8cabb969ba886290adfe6a051083f3e327709138f225c21e5e97266c4bc3851d1e50cd7bbbef30498b46c87f1a04bc0c9d88b7eb02638fde9a594267f93a5183908a9fd51976703fd9f912c168b4c811b70d5377448ae648b31bb756e69890ba61815f97844d8f9301fc6f76fbc33577261ef2d8830176ce0fade078f28e0322502f7324f5a27e533c2ce1ce9b2e804bac9d91390bb20d5a75784cfdd8a47812a8b22884af1cd056103ea7f8e98c938e325c40ce89a759b1b6602e47dd37b6eb7da0e00efc1915d02e8cd9a6157b6a3c0b9a6fad7d1285d6fc06e8f95dfefaef6fd2632c15ce5c19e55512f0f8cf8427d73924c57461989ce631644896695e680b48fd4ffc95f8b70276a6b21fe139b0dc3d05b2b98e38fc1ad509d38208d6bb9228d6c5043ee576a32309dab8781bc5af6538833d2afede32229681c41191a7fb55e16c982419432f09409a36489ac9debe99acadb8cdcec1006329ba0615619589e6bc2b9583c22d9b47a4b006ab61feb3384b0704e669ce5f9a0d3ad88a9a8d14c7b7a5071906b2ae89171b1107c6709cd7ec8925183a40cbc36e413e8f1f08b4495fb48c9e45326921a5305d892396398bd063b74f4d2e54cb168b94cbefb0c145cac7bc4e6b3ceac32d8997af4bf6f6a9577cf67744a9699de1cbb53647ddcc36c292a993098b0f0a8affa914b90605f3bada06647b84a895d39f74b2b644c0bf2eec6ee67e7058e7670029d15969265530f595931933168962e66738d5e726874f4562ab7ff5b092f4a39c836d660683b68007f589463a2c8295d7c706a71206ae3e2124f47726ad970ea49180d09b014f53df5327d8e97b7b6b68307e9cac8cf9c65d202e48691180ea175b19d7c6d2278486379357d62b73d484cb2ca9b0f8843a80d5e03ecdedd7067355d950483955782230709b69ab36435111b6cbccef753b369fc9ad01c3dd68b29202fbc68d64747fdca126ebf5c47becb58a529790d18f76f1e7e2b752fa56a63231954811125839ccf64f72c1703ab60e723eb6b21b920efeadb70096f99457c1f5d1054f5401e459ac07dce46f33a63bff89424fff555ecfea046734c34a5135a87f8742a1d0675076e92b0df6e26d7937214be599948082224f238c10db5ba838044c2740db266f2d73ca758df0a0bf1a9d753ed7a5555739eba007e28f1bb6e47a0c9c4bcdea0e2469d024007052c8d76df9983f46c5a21d7c2080d05ed6603b0a7b29034c0ceed2402e7d43aadcf1c1938147eea5a13b6980c95649152ec6a1e3c8362c8dc94f0cdb4de5a39e41e619114f4665a027850e4c6cd7b0ba23faa5e6d39ef5965824f253b8012d2cce268308f07e546cd26b84f41ec482ea64787829c2c619cfdcb8dab37edb299feea3870beca03185499f3bf248e2aaf29e21f5d13b7d5a6ef77492861e1ed660b3278fce14d321d18f0de35e0a238e390a09c9d2001ac765dd3bbb5978930a05be160635db1780fe6a3c114c1007abbf558dd9dd517bf5215a6bd76f5f011b759f7760072cc1aa9fe8554693abf156c9d1983b5a504de8508d7f72e1e083336eb488eeab564b2661508c693c36be1fac1af2f3a20dc623072114c8b96d5f250553936a3af8ca71da4958e95eccbf9ff5e0eec9a3d0b7fae1d34fa979e155d71e99591e0517e017a88153ca121493851717394d3bdd9cd8f74596974fe3cf04ef9af1176c631dac250feca831fe839ec3339000f471b2ecc6bece8462aeceabee6289915d4ce86ab1c445f6aacd936afc0e9f215786c536e0f92dda6cfb8a5ee656da582b9a215372e16a30bbddd13c26f827bb0c4b4c21f2c561c9bf74e98c9b9068e4664313c22e1ea103b30078f40c82df46e61496f593dcc9542e4d9ff39f27bfd81e437eeef6b713c83fc61e7f55f882b08238fff1b8aada0ff358923d08b4a441dade4ddd3c94a94697815da5ab00ebf9d4920c73699d6f3cb0180ea76c338ea53ca44c045f7badad732eb3bb37e2c2498053ced21f8d257154a4c73bb2484c31baa0abfb3e575a8a37409a05273572914;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3a50f1cdf411852d28786033789501c480d7259fd7be716d92047c3dadfd42135537892c63bc3a4b3d36a3390b170fd32a6874dc711218732c7cb607207e99e75b9411d2c6b5c5a529c89328876909632ff63c7d1297747644614630e5bd497a5bbd676ddbd8af3b95f0f052f9426c25c6abf2716fc86f52001c1f5964c80377744558a6d9c01e14a3d053a42fbd8da16c6147e418c763bec3f2fa47bc3dd8293273549dbb5d857e5b33501f6fddd515d90ef24abb58a72eef06b871f6e218127ed61d08130c39d6b44e4b1b6bdf38672a50f27bf2d303920775d0a05db951d1f209326902957b7707f42e0f74e6ca09f795f5561b2aa76f1d0ce90a7e958eb004bb14f0e60762267acd3bdced703b2edfbdd06dddce984c684b47954f0436e8e2918d8566285a38fa7b0c527c995c01c8b2918aec9a9288a151d59a848c7ca42c5eb64d71b2919f992508cfc312695ab3c3088f8f579e8c672db8413f4d36455fccd203bddc246db57d64a8376d6aefb25ae8fe8f143dbf16ea890d4b125419f6cca6e8dee66ee218e4574ee31db4ccb797dfb502b3a61814ebb54fbdcd74c3c4170cd962ccda299291d75ee9aef5df825a16659cfc711bb9fab7b25c02051ced8c31db10ea1e95ade0fbd11a149fcb78a45fe5cecc6632eb36c6fed572bc39c974e521f34f70f6cad4f42b74ccc5b6ff3cdd129dc22dbbae196ff58fdea1c33043cc8cbf2a1b88d10936e092599472e79a2a122c12393f36130fcab2427710d28ca683d7bdadf9076fb3c7000d6b74b0179895cb88920aacdc452c43feb38ef071d28b728bce38e5f7cfe1c45ffd76c1a23ad6be6f6297e2d732c84c1c11dce22fa5dd4d3248557ae2e0b0fda287b4887f407c343fd64a591934f7745f24df6800322f10ca8307e474059aae9fd80f186a83cba146c9957b234acb0583220b41c461bd96159f4b155e9cba96ce33b6520133d29fe30ed015e0c98bff52c1f88df0e56c929df85255611b067b3e16feda2f5229c1cc9305b25155ecd259f555c1e9d111daf786462a10467ab523dde29b564796ee6601cdcddc3d667c9457f93f6d12b7dd216de63908a47603bf1d2a0e5a9b3f640fdea9cefdc9b4fb78abdef0556c96367ec8380f68798af3dcdba44f0ac1415f98303a228e13413b761325a2a78c68648c7e069c6bce30d1bb0d209bff03b330569e673676a9a27ac0f85be6be875141a7425326c8e9cf9e8da690ef292a09f6e6d21d0042fced78133c8628e6076607cb8acc86c883ad6f90567cb32d6092396c20895846cd3b1d3519ba85b346b100a07ef2a279aaa45770df3e075e7b46568ab64e451b0856a892d78533f06a4ef3761eda1bbd1fc30c7ca5a0ad8db6baf32d39e5278345bbc081acdaa0ddc6556e4464bc542b617ce7ae17adaf6deacfd0dce92a68c699917132f19138cd470635070e7985d0f07ab27e92aa1aa7b9b1317403e6e15e12bac7bbcd1012ca7941128de40bf4317636fd18449376d50542aaa4da1c8cb5a5f643860bed19ac70751a8ece6f1218fdbedb258cc893f7f94519ede0ba503da025254b67f9af37be83f74f6fd3f714342144bfe6bda123727eb113331fe5862848a845cb6b6948975c2629653d9782c176979d6df6145e2a469141124fb6ca84f29b5491cbef3678f56ecce3cdf64458ac1630b200e05e6fa53aeed504116a430a0ed815477be2ff02f912b64bc22cb5054c3ccceff6f02b679774989edeec042f1cc2d5b812f7f9d94ca3b0949649267ec451e5046429b50f95f4fe1ca6fa135881290f2cefc75d0459cbfc018ea652ae32adeb54feda268c63d16d1ab6a4a8cf231810f9c9da0210292b33d1590e2de97ec9da9a8045308fc50ea2960559465e7f4cbe5f5e4941b2afc01c8572d6bc686e72e53e6174a0af409f86d4b06edcb89b42279ee856c6c820f9590b980a5db634d07442f84ee529db93f92b42619cda555c1d0ebc676fdbda7ac016b5e86e3db45d175123ae46eb18a013fdb78da180776d8bb99f11b15341288899820784fa6bb295e925e244f69aff263e8f9602434229ee3f55935ac06f89b3a5e5ba596f1dddbddb8916c8b85eb41e8828114feb1ae5b193e0d1156cff78877eb384429b90b2104a2188f7020ddcb3699772af402f7df8e17b2c689a2d61356c93cb58ec4caba8c5939f54487aa7df73841ead3fa3cf9b669a1e6198c230383096feedb3c658ca5a08d08b6be5017ee662d4195bd39a438e2202db49688ffb67a8656d06584e2cc7bbdd1219a986bc4faaf38e08a56635dbc477ccb143b15a0101a8aa884114eb5b5829e737bfec6c0915db2b5ca776731eb5bdb25f02cb39b41554f1088457c82c191e35400bfb9bf2f39a28bcddcf17e1faba68611de80a313666229945d303141bf87575394356b24e6d27488d958e07841885cef6535246546525880c1822263931f15bdee70234c95ebfaffe97145441f65c44a61c8ad25249ffa2799fbb6c1f3c8975f606abf70b8e6198438d24449b08f35bf4b2e1e9b9e4c58b7b9eeeb5f33fb0706fcfb406e21b1abfc3ffe52fea6a41b1d95bbd02069d3e7de8b74e6db0d1bbcff7dc6084e7b9b9fcad4c5ca38f225c878fab392142dffc859d21aab2797852ae945163e61ebcdfb7e6a4a74237574ce7667e455a84c4cb27866a1ae53f8e24d3e49b4fdedf20dfb0ebba6cd09175921e096e5f72c6b5d1501a3dc5f0c61e368be697c047ca6152af729b9c76efcc2234392d0511611f31b7833256aca5c0ffca8cdaa6f883c595997efca8069e44deef2186c6c97571e7a417732fd7161d18638476d2a7c9fa475437e607919906ad0452674230d9a48988fb5167b9840d5583b87701720741ee278cbffe28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1c8ed19ed8f006261b682552e4958767abf102936f9c00465828171bd431cf2d1a72e1344098ed5a4079316dbf55a5dd9406f1af4d5f6720af215fde7443ba8eff9ce3cbcf20fa23bddf48ae762cb418d4348b2a113682c7c70594833606d7537effd5d48a1270b48676894f9d4a28948b6d5bbade4e33c33ed26bf5fbb063bcf3d8f0dbbde19bed60283802494f106745131709146190d47eb8a8ac11a2f44e5d12acfb3b4099ca67646d883b70b493155ef5795212eaa1027a0438df961a5e30a980c11dd052a125f2d246f50b90d6b523a7b4910ebc6f8180ed120bcc89938fade3164ba9f0c48e3a02dd96e2d01b39ff3d96762564a06bb72332219822c7e3a5a3b88c5594bd954bf6bc997d5f91ad55e97e643d076d97676e131b919faa2e7bac55ab1776ee97b4cad458abac30000464b7d7852c3abbe66b1dfb4a7918a1fa2943f62fccc56596a05968db05d8bea8fd76020c8c671cdf4c1511d0c5eeacd4a5947e3c6bc550c15db511870c99c4cb2f9f20ca8faab158e2d959b6c427cacc4f227d280adc28e10649ce54a56461178fae3ea2bd64f19b83cdbaee0c5bbb37f97c7cac917969b6a9ee85d8aff5240c977f65b7304394b1b2073b57c55829004da229ff73bc59ebe6976ca4ec79b076748cc3255441984820797761ca1147309e0cb2d13054169dc3d1e2efa9dc807b61a580d990554f5912debba1d560ec22b5b0b63a7cbfd07567ef1ef9c4d1a5e799815852cb345e9f044bf83442128b6068ef978462843f7ed0d58242c43de73fd76202358102e09fc5eb6f7ba1276c3112e3aed6d3f9a8f08a98c7f75cddb14a3de5ca74bb5860e20d5da2de1d0c5da993c81d86a4f689c83f169ef1974ca15b444f005d0c04bad6a11e90f770579b2ba7b7161bb4995282e1462f5abc30c79f7063baf5c369f7dc38443dfedc90b525b76eb8152eb5ec8f1c311734079f61682cd58772b98a226436f101f075858e215d302ef89b078eec5ccfb5f6e5bdc72986cef219d94cdee0b918611e4a550067a8d15d0b4d4b632c67bcf1800eff16f0e5f4e93026f7a91cdf657660f62f984607c5d182e8a2708e1201e197ea941642104955541c14273590a753a1da560215d69929e9f7b2ac6b695c2303c5f03e55741cfc62cbbd6b264eaabfa042b19c26465939874a6d79d8cc99df4d050e172ac5e5f73bec43397b0b2512af5a8be30bab07c93c7b8daf5e6271d8fb1a4b2adce8bb0dbc36cd8e79841afcdb7fa27cd0d67c7f216809ff659ff2710163a53a95cc43a20799b95ca51980071436fbf01c6337c100ef0b23f04dc12d7b6c2cb236af368c5259a3211796a6765a367cb70f46571d3aa1b99f0b343ab71cbb639022d34e91d03a24b99eb457760d37eb0237b7ae119de26ffa67d3a4d73c353b8fe4817915f1c29790d6ad66e80855aa367c55c548db77093e6803cf78a1a5640592593da32e4e49365f33032c6542c4a1bef51f6c947cf5267bf8ae5397ca7b6bb0715dd5d8177a6e8c1e3426b45a20571e47ef9e2f9019a4eaa1755bebd9aaa0b046ca8a8402b4aff98c240692c541135f835f2083d8db5e5231872491bb5a8fac47f92ee7bfd5a4978ed68451e2762b5d930293eb0bd437f24eddc6f39b8bd9a2963b51a514e02a49d2ebb8f7e3439d0f802213b05d92f8f125253a2e44379f59be03914034682e6ac7b7a05284b14f55ec741fa1ad2aaf7c3be1d8b875803f7f05935c486a0f10b7b39e4fbc7a6307b83528d79ac1f0ca81bfca8e2f64d8ff14d598ce657c3db7d812f3c16b1af1550f10de3745e2bdb94544e6be85ec005e68d2c20e524d42055ab957b17de506ed2062f885bafc8f1f6b96f98d8388ccca5e505053137c9e2ca0d57ea2cc5250488f54e0de5ad7e56c4303083cba6f4fc2cd546ef8025a5604d557307bd8544bb6b83e2c8a9d8bbbb22c700a89d73e6ddc14517f369350f9260950f0085828ddba7b72ebe8be4b8e65e39a2a6a1ff2d3e0f62833df2429de57bcd0183afaa720ab15556188205b78416e1c0100721d774f31e8ee3241808b9493a574641f8eaf809fa4f072bea47f5e04753774b3e154153bd134cc50a3ad6aa3426e928e279eaafb9e5d9e66e0b37c9a39d89f8f81f08c9fdc0b499f74ce1cefb0c5a443ddf130ffc991db483a8bcf28b55bf2d7d29453c21ab2ddd181feb592398a9dc78de9bbb0cacf94769e95f8ededf0ec80becaa950c8fde47f4821f1b1b8cc068135b2d1c75adefb4b3ffe5999e35f1585deefd83f19ef120a7392bd0639a2a1c580f2ae9a21b5c7136cddc01a19f3e139a760c59ba2ffea07f0a8da29dadad4f15f58fa9d44b8f6e66de6d885ce495868a957c22344b2bb0f670fc38bac9f2f110fbc1152affdfe89bb6b5148242c2dbe467e2ae918de0cc1e477f72a2ea42e7a04e09f9b5985759bd8eaa4bbb32092df6dda09a2078aa0f593c3ece8ffb52149e9d568853bbb7d9ea761e6ecddc014b1e74c8f59612726e0186458df22c27ea5b52b4f97fbe30f666400051f490081da50c70eacfd746d33c97905cd46d79099b531cae66d2e310aa044698de89f77ea6794b45d87a1e467d35ef3178b5baa3704a17a84c818128cd1d29af9a8c7ea7cc717476209ed4cf889b50381d50163da620224a0e5181d0d5e35b14b1c9019705d3e785673b1b9b0119c0deb37a3188d0111fe70477804d86aceb7e2ba48f8d83e69b465830c0d261a25b4aac9a613d5dee390f431947f5aff5143861c252ce91d38fe573279594684774f989e7b5a3a1413a736834e852ca73b4e00abbb217ec0fd091d8dcb20d1f6f77e6b176c24b877bfe960c3f484af1198181ec73585a21f3e43477a09b3bd5c66a3fe53c1a8056b5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h777b5475588d1701de4ce7eb58ff35691f508d2ad618644ee2caffdfd11e32414978595158cb1e64405cdf4aac1b7ab567918a31ae2b51cfad57743635b66b3aded2e23e86ee7a58d0bef45c168b32289e0d5725118a5126c04a5fcaa4465841d0aabb9abf5382b3574d457f7117f7ab289acf033c0f059dfa7ae3eb341938c63690a5d95bce3e50c3467528c5d11e8b5f9fda90b0b6947bcd81b5c481fba387e72116a62dddffaa210c0018111d439c91b0ec17d50a456edbc0e0103ef32b49dd933e39b7ba61e8fe9d0c2b05990dca5ebaecab515c52b3b5b99847bfe7923a1d7b93bc4ed39f46a98ade795a0815736306df84cbe93bc26cdbf533c6b7fefe191f060d7e0ceef27086f91b6a3083811068e4543bfcbd146848de192246aada48a5168ba147ed3da315ed2890d2f8d02c504dd09ecf6b84ef988b2aaa54dba90d7eaa2b028dac87ff087b55e7391bd9ba2c73855053ba809fdc3de8c161f504ba65b991d4334b644cd6e2a3585bc4ed799b4d7aaad4255b80ad85a4c12b17ad21760ca6fb47d2f1b656b1a411feb3fe2fd84c242bc291084ff951657ffb6752f9c8b6e016323d8e4af24e955d52a7af3a4ebeb233dafb8cb7cbd0e8b3b521c333bb94e5f30ce1183f505141ac93bf9f34c806da5ad1cece6ad89aad13d4c98b5c3bb6b0cc244dfeaa31924b13a1ad4eb0efc5e7a47cab8754ad2aa78bddb75b581ec92c9bfafb3d5a1a948ff8922347018f3178886cc889fc9e7a2da013f8cbb93587b52728bcb288d476d64f1b6b64f7cae1d3506c1e714d33b2fb211364df80dbd54739943d4b6089d4fadde64184d30f26551f6691bc865dd988b2ee6343942e695a252d0108f3eb57890b3ac7417fe3fe6569b10a1510953a0bdba3e4843533a7b32d86ac91f913a42882fe3bc8098fc33ea7a84573b1164274e2e8865a8cac39f16292d8a4a9e99dd13e07e8fb49e4e47730ee48761c7832ea9a09752dc81c532b104413bb4b7a965be843ff940f6f839f370e00bb5f1f61cbc6c014dbeef30a99193de1050816d3d59218e169636986f63cf8ef76730ffb09e8618141f1c6c55b40055b43e77db132117871c4f15958a7b30591fd790743677387508446be96bbbdd85b2dbd0e029eb6e290aafd135521a3c9b7dfb098414e5805683099522e37673d7cc55748d86e33aa290d56862cb13f56a930571f953acf92c7adad1249f1d240ebb3e2fb414681a7f8575cf147ad177762b675a664d51307ad4ce9edae7fa3d33612cd90982526c43606b0bd898bde3369ccb8f2e14bdea38929557e6b3f2e4fe4f6423b51859c0457fbe2f45e065ad6ee0842de223db7a2408624a5c21fa0014e3763a29e4ef4e9fd7d353ccb68f63196a3838d86f88953878b779fd0d4502d9fafa9d57db5ffc395ff9a069029a92da7757f4b7b87d6d7df95d82892cb7ae9e8904542a597e7541e4e28fde3a0b1a261ef5509579bc5fe855a7dd759b30f5615238cc2b56b6bc1466c6ec96c3b251f3e84601b4bd6ae5fb45e1c6e934f397c9fba501c4772273a0f864d86389ba22a73b11ff66357ada5065624206d9fcb409372aa0dc1e3ff66306bd4625c9473630c10eda141883c8d1f6f4b370e5cab910a2f18e190c05d271037775f5f533db0790a42d718edf301be3407123306a7fd77768695d4c2da58882d0614e9609c2bd3ca2add5b17ad812fdf3f625f609b4f2372f63d1b67a688b2c740ea840590960558c0324cfa3c3688dbef0c606f83ceb10929466ea4ba0af8f67dacabdc99e139e0063a88d89be8100cb47c5d2020b55026991ca7fb77b2deafd6999b6a0bd9fa6f99a432ee32f2ee90f8defca86f1ac5c3e5f7e857daa140473368468183f6e47653aef071679531de36af84e212035cd5f08c9615de9e1d6e9dc47fe06d027171b13b5355d10ac77fbdf5c4fc8644ac30687343fe1fd4fc1665eb31929cb6293b8d4b95910412a7066e82a3487d7a2dcf920b81b5eac0e7637aba7b51a932788f24ca5aea892133e6fa646310027e6fb635f5c69adfcb0a5b63bbf5ebdaa0045399e5addf1dc995c4da50d4cd83d9f0012e24096eccd12365a1ba4494b4e9d94f5646bc33ebbbce5b3b82c16a1c12e777d606bcf13b292d988c20dae5611594c764c34e1ebafdaef305b5dbdb76e48f46d0d92315b718c03258e5d94fc0048b79ccaa425dfb965f1627e3d6c9a22d484912205a6bfa0c83346f4aa0e042d604dae1922ba3b819efc1e1c3b88246fa12c3234c4d03eb93d4f1c28b4b7030db1119d9752dce7216d511771f3d2d0badc547fa3a9be1cd6e074bacb9775b99b689041f08665b919086cda240c08617a47b890952685858cf75069fa733b9fccd004e8ff2b3874c35a72a84af0109fd3bf64ec93bf0ac35211d45b12d0dd6d03ce77887d2e36d48a63330a38db5ee9c3d0a097783784a813a83a68f6adb458d6a29688b3ba99fd65bb41dc30c3fb6eb8059f829c3399b8c9ae89a59478cd7b74514f1127f3f5821bcf8af6f2dc07679ef922d92cff8da185d3df160c72366a62f316b0f05708f1212292cea71b9e5f73e80df307f95355415e127019cc71c5388e9e14ef22781014f9da10fbb715fbc803217946c939b7460f35ea24f4b01cd8ff3f66f0eab1447b697aaad16b4095ba86c3f269686b1f314cecd5f1078661074850f3652126ae77f9dda2b5124d61b3e02c22316d56158c566d8c4e9b18dd8c0555cc89d7dd4f4051d0c67da63044260a4fc5a4533e1876dfafe1a1ba9e7e1e0b9db7c95bde579ee92445db3022f637028d3c6281557b2cc1e98c15296c8b8aaf608a817cb687e1e7375ef746affabdd59fc4815c4ff19878448f4a2b88f13226030e050df2b2ed30e54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2a2380ff682cb5f9c3072b9d8fb5ec8bd5b0ed805af3b21f03a3a4a186a1861a0412ed2d8755188599853b1740ca471f32d98b8364930e0f68a3d8d6865d95b3f45a229a776ffa80190ea817f459a9cbf41666ebcec0ae09acb457287672571df75720a30884c665278df2020fe4bcefaea5fe78ac3416243e808c630b04d2aa9bcd3f30fb8dbce87eae7794baef245264ac6215ca1ef8d5a27be1cb6e57f5119a8b038b6687b9f98df81e4f3d0d083da0d992726b6dd2ef665a47c1f9a504ff4b9d300bf0576364dce6e5e2e4fae3d63730a1a74248e561e3cbeb3033a90db200af9d5e7461d44848e14e985cc92f80601c6c8e3f9b28807ebe22147193790524f943f2a435589f6367b503a389c9d191498851c820b79e511e4055fce75ea5c275af411b14cded39f252b82f67ee0cbe979213925bab5ee2d4903d6781ada09105d55036e12ac376bd8430b03a1dfe74005ae6b898543ab4e49b3ceb3721ae7d7856538ff86d4111f54b380f8370fe65956613cb3bdd7b9c8b252ab2223da63cbd0ece55330faca38dbe1f338da807df9a1435601bea865a3d89d9bc9c02ddeedce329dea86a1b440d0132bba9cc25af5ea6f4baf2e5c56a03f2445bd75352e030fc9dc374c606346d9fa901ddca0d04841c43615c567032631f26e1162895ef4e3218894a420b1de01d8a9031b5c982e8da86fe9b3c762f4f1f3ae9fd1e372b7ce3aa7cf31a0905b7b8d7d6bcafd61b8a991eb3427575f507d9957a8c2fdffd96acb539103b2d80c72250d5916f936c86bda529c4c85ea43b5e463ba89a339ee2f849cb0dd21ebdb8dd6f2850a312ff2262b5db206b6af9f63986e2b20d4ac6e21d019f5aeafaf92bdad5819fbd974cf55da87cc3e92fb4a20af2b6218e532115a2db036ddacad7c8f6e81bdc3cd04c961b4c4ad201063386df9e77e859de5f6f23319c9723d4df3c317774d3b67dde0d499407c7ff2bf947d095ec235f37e3f903ea373cdd36bafacd45962c1e78f67cccaa571ce3e60d309b29cd5c2d686c201268254be91a325b89ebd45a803de31b25a1dc12616b8cd939a5647181613c48970f8c6600f03ccae944d26a47fb90f899a81677d300f871a340324631ee7b901fc905f766f0cec4ae5cf6295fac5b36ce296d0562c265943a637f0f9c310c5bcb0ea7befd481f814dc35a838f6730a69bd22f641f64a55911bef439550cd8d3e898ea9173917b30730ea2497581bfdb5984219066ede857ce154e89ea67c6add54ac3c04cff220a239bdb3806b42c2abea69e20d01127fa29fc1b2ff42d5b7e74e18b622e2c61b74f62a00aa0e667c01b9f76d268d4de309753ca1dad581610affcffcca9aad07fe577a33fc985949061a946ebb8bb447ebbe3243ce6ec9b53cd1cbc307a0d949deb26fbc84181175438360e09509f795ca7fd89281063845388ec3c501fce3a78c3408591a5bc1f6de2145a6ff85c4a6c4865dcee9e6988cf1b16a69e9970385d92e16c5d32b83ac9205f9f69088321c1bbef4075b6694929f9795ca129b838f6559ef4035c32443fbe482c27c4243d3a2f17b98d83770177509c613e8b2ad6d4d3a804aa8707bc98544f11c9613f793846fc213f3a9a9464ad42aaaab8dfa76d5fdc0af02f8ace40a215bf78fb924fdb91904cea29720c800574739f4c9ef279d2f7f56318820b24a394b61a809091816290e9874e763606b97e05436fce84522039f0d59b08cc7868c0e7ac946116fd14274eb5897d4b483683a0ebe54ee30d65774bbf69b8acb0fae117074c0e9223597b342ae49b69a4efd5b181a21aeb6258696a74a081e337b175ca694dde7a4b4873f8a6c36d0d27bafaa36f3a4c5a29a40b5fde1257d45ef78b5a313aa70d74338a541a8d905341eb7feed0aa31f2acb279f144a91ecdeb856eaf2da732e7589016077e395d98593a2aadbb564beb0a407ba047eee8c70e5bd335cd30b11d2acd346aaaf59a0c6ad17efcdec10a5b09439402ebd00aeb668592190dc2ab6466c8f2861501e30357889300677b572fef86d00eb3b2f860e37f370dee8b430d9cf542834c5db77441feb1cf3fe29ab6cee73ce1ca60e9ead4277807acb1cae0c3b7eae1ddfbe03879d1f814d7b3c1e10fbfefa15ab1c36614a7fb1a2970f6cdc99879136035a0639bb0fe0469080d914e4ca90123a277fdc07ac5bccd664a56f4eb616302911a92cf2425e0bb822c563310f5ce7c1da0a312d76ac35901e5bb23bdd0c5ae3785261d494d554a7b199a2afad190039a64a5736083f15080ee5684aef771101a0dd54a1d4ca53e3168c3d50c7952c58dfdfe49f6e9d9b54fb8d29e2e88efa770b4b9782bac375faf3f947ba24ada0e6e4ecfc39f8634dfef1d80f24c844149d3f92e08e9ed09f9f8fda007adc99c6625cf5aa692069a69ffa19b1a709d20b72aba6cb51494460f651e6d5ea62058361a772e37f9d1cdfa6c82599b036434aa6246d6c2e5255c0ec98d6fc38bfe8760f4f786cec5d9a91df64384673248974726ffc9b9fe50c33a006a253d47469921412d3d54cb8716e79a444bbebbff2494315b585a31e27d261743f020d7b6792da73864d5d456435ff2588122a63c508c1774896a720bd2e0ed5afc1e771aaae29e28b125e991b3a499f5edb1126749f73ce24ed5809d5eded274ba55f8d73292ba80f74e5ccc9e958720a9eadf94f3fdbd2fcf46b658332a22a2771c2a53946df5f9f6e1c9b9947cadad26bfad85171ef8bb601b4aa91c5f5714c2b75e8533a1dcd59fde603ac55eaae40c27b31687f3c2e066b9f3de7d5d5c37a0ad689e2406d56ce16102a7fc6ba4627babfe2eda037a96d0a4f0fe7937842f043e78eead78ebad7d01e01cdc1487896c4bc89742658908;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4736d4c340809e4c3e1abbd058c830f3b2caa55d1220c6dcd646f7c304fee12c9658d5f6bb24104777aeedc475b3f268ca268e938563bf6dbbd2b738fc91fdfcbd14ae9807c507884c9930f087891d4cfd5c06c3d1888e079482b3beb4e1f2ac35667647cfc2be2c7b7834a1d739a86c0bc056c2465fd28a5ac7f165526d42c1fa82b7b1d0e07c5013d7273a9e6617fdabc7db0318aa1c8343467e8443ccf0ca2553405bbd0beaaade83255108179a4557e80d2eac81b769535321c3b980ef2e9e1a98db12336eb59358a6f109449edf76d44bb2e2c0660b145f48e4b57c0cb7897286f752600666404ea6e8a386d55bddfed9b4416dc6b855fe182f06f3bcc585535bbc04f6fe4601ea51be6d6ca82ccb2b5cddd5a4686de8b385ef41f21fc510b9a298a0c441955d2193c4dafac680e1de73693228c3b7351df8a7f6d5c254a4ac9b931b5af333194eb27cea01b45f30c56ced9075161904336ac63aefae16910f6aa2a31b899d6fdcc7fe44bd469265efa0658eb9f95252dbd859f9e96ec3de8a17ecc1f49f42e4e04c8ade215c7b0438976d9fa9e9374531479993e99131971a3ce9be31e54e5f2e305dc34fdd54ba286e868a21a2c41a4873f485a80b8b464d910f76508a8d1b866b9a52b665ef1fb6556892721a07a5a0ea1a7b05c0cfdb47dc48a81bf0ae70e702a67ff3468b658419a7c3f97db5340187418a466a86ac599e4825176493b9ab189e1ded67fdb259fccb46fa53b229f8d953d261946b22ff8f91a68a6e11ae30598b7ff0e6b17351df1dc3a8fb33813f6032c0bfc49c7ef3f4c18a7368332f6c28a362344e0a50fe4e5935c9cc4ca9eea7e057b44b6d8600ec8385293b0f584133a87f1959f31e718fd18d680a23dfc173231a0447f607604bf8362efc2df1ac7abb6850e650068247e8af739151bd6494ea4d7f02c57958d0277ab0268af79f7472b85f8a277371aa8c87aaae3bb59e50ef3be8c1a46343b25d7b13845d94d156c0a00d354ead58dcecda60c21dd048daeba00bb2b3d801b2e12384dfb1e5e1b0b8e671126e63840f5875761c8d19df1077f97fa8f22c95f6a13af6c84b0e945c39870d12a01f635f9de12b1c400859fdb8a8e0524953c3e4da6624114d21b89926517968485a870b1ac2145a594aec44544fee947f76e1bd238e22b49ad734ee67fcb339af990ace2d85ef8e0704900c0b1a7632e058793f05a58e4915be5fcd048bd6bc61baaa86b67009ce2a498b24c796c05b32c82b93530978fc2e92af23f7d71c2de63df9838cdd986cf943fa024b12e3442e641cd3fd929d29c847bf59202bf7770221595f9aeaa79cecb5f2af0582408c7b50d6055dd03a189c59cfa5bed86bae0b2f259a55d83bd077f99771085b6dc90e0758816269202a3fd99bb3a387cc1849d46df3967e3fe390a16129fc9337c910e3ca614829f99baef0719cbf4259b7bcd94ce2c993a687b8c65e831960002fc930297ba8088a46e035b02c76f195d266f74154820431d3f4af89ad05574eba1f19a6611f7987697ea7a1b562fd10e3391506b48599d95dc8d8402d86145cb63b99c954f370c52012041917e529c38efe996a96010914b9ba38c8acafcb90e55aa2cc647b6b60c5e56b909f4f3dff23b7b149b8f0ed5d0381fbdba21a874477d383f0916f4154e71ba4b8619260c49a76330edc1d633ad7a9891ae9271f5ed375cfdf7e45d7bd1e35815112dc882ff077486ea35777d9408f604bf3b2416fc763d142dc647b138958006dc4b08dd6602e31cae2ceefa8bea5a85e690035f7b2b4a4e4e7652b8180890c5d84d91dc5556de1c9ae3e645520bcd293bfbc4d7fe15016420eaeca4d08edd12fcdf64f5dc64beb20e03fd36eee1d495393798867f0bff707a3447e2c6766226f4008a259f284a15a6c34cec2fbbcc7398f8996b5f3b42c35859327bd601e468f77396534396adc3bc408406ff1497683217b2d2bca30e958537183a11895faadfcc6b640ea198042512721a6429536dee7f7a75afdc04aac7e7dc4d16354f95c130185d8f56779413b6961d24b6974a035912a17bbde2cc5e88a85a12cdc4fd049ade1c67fb6a4425fc464c3bdbca12538995a30dd2a92477281dcc6a5bd2829f44f9ccdb643bb2183bb442ad379e247d3a4c7848f59b54846292d351da34e9cbf82d7d54176d6addcab6db2837ab0f2bbc564d40b59f7c7510c7b3ad48e140234d386d6ecb363f063f1e3a231f80bc5bccff5ed7def8b82551772bf4452796105af5b5b983703ec2997de541bcae395bcc9161039e9ccb07acaf9c6ae1a137c02bd4725a033a3a4822aa5f2a0ed93569eb23aa7d005b0d00a84fc7ac1b89aa9f94cf8207b5e078ae25bc67eaac981399982d6ee755401944ec9750d3287e0db348b94941e8ef759b5f5de0f28c2d68e355718452048cb4a89d09cf4b0747ca699e98a480a81fca607cc42dc147ce4943fea3b318b108458c5d35fc532ac1444537bb7e7ac80c926ae5d511576f2aeecd3ca46fddee00a72285486518dea1d6104aee9ae249c80d1104f072ff24ce065e541e21093df38d732051ea354d7e49d72cace6ab5984d5eea470fda25515368b2e1bfb1d604c693fde3f82fbbb6bd156c3fb8b039260bd88f9ef5ee05b5883ec5d7812f247665c01be151567ca62da28d8d0cb450a9f5d7899da034d2f8cadd3723934ed59df8568dfe663dc106a54c8f639a2f4325413bde49417c7ba51e4e5e0771b20d1e9e08d76685d1d8ca96568ec548b9768ab63390df9c7acc24941558bf2e382ade14f1fd287a13574b356b04d4a0dff0fde68faebd1477ca5b110c3dba04ae49f3f4ecda51718266f776ef7104cfd939aef3dcd0d8457cecc70f05c3d953cb3b5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6b4a462c72ff07dfb2c76167238318fa6dff3e31a7434836f32d6932f1beaf17610af80cd843401ba4e98aabae883a6699815a32966c572452c3816d862b8aef5ad2b6a9d5f03b1479d1f4c740f66596b375fd9a0a599795545f8c9e8977a6073dd7a8eabba4f22c5d2b4e22c12a31d7e9e4e97c77c4ab20f2ee340097f335715747268c59598bb330ab051ce6a6c9c75278bbb0937b9e6cdfcc2e0e607fe72a4908aeb1457acae5ed558d5f000c31d9d540dd59548788680c064c3ed83fdc821cddeff153c7175b3687426313f4849857faa07cff8d24f8d796ac60f84711f4b2c27e06a90dc493843bead415355ce7bdc9e1c9284b5c73adb1d0b29133f0b9fbccc1ab786e89a3cb50bef9d886d2a6baf6f8c5cabacac013759ce4f42eb18d7eb7fc0387bc189feb50de11a36bb4827ff0e15c5738da253ce87f4d7f43c2ccf51e4c2126909a710a11fcd1c0eafe948c787a3f031b65464efb826020105b49f71dba9554acc1f75bfd5575155d68514b88455cd6bc10c9c5dab9982af424403dd3bdb93184c4dead44240c019c58522040cd9325ef9895c97d3167c87335913dd32b5d0823117342a79c97da6a402bfcdeee217e31a323004b7d6e4809c888616c8d8210aa12c4296443e9cdfbdbb5b41c6d9a5ff3192f78a077ee0566f2a5e95f95c1bf09882f68090ee65baed075165391e6cc4a16579fe5b9cb93c151ed9ddcd0a6cb3b7c9c4263f9191ee955acc3be2ff9b0dc9c1c4052d3f3ed9f7bb7954e1016ed2261584b36aa2146418b32091aeab174d12d6f75f249ae9ef3feb5cf992e24194e7fe300ff324b3be400cf8dc07cab3dbc5ea0feac336ca6a2823bed971eb1a918913c6cbd01b7b0236155683837c7ac35a29d0716fa3d5f38570c368d251aa5949c04a305d1f9d6700c5d9f99bcd13d3f11452476a6b4cc41e839bbe08e41e6159b129c82ba26818706af0ef10f792029411aadf5c42e5d00c5d0895b18465546e40c4d6f8fb202346bd16383f2101362ae0866c99434aec05102bed8cca3223cd6ce7cdd5a12b9aabd3e8c71e69469a50cf2f696361c14a75bb3b8a863470ba2eb68dd7d18cfce4fdf4077df5a812198884cb2b6bd5d76898a6a130967375f673cca684d025c4a711e892ee66839625eacb5647dd10aed98d5c8fe6c676f820d97a5378badd76a986a561ab2e80c0eca9939c887a45e2365f823aba3e8ea67344b203192a0d0c842ff8d91bb1d7545260771a1d8ef2d2bdf1f5c8e3b524cff67701f0ac8bb3b990d5806b2babc7a7a0039c0a9551dc5f9d064e7a0fa2fd1c57059af8589077455c72ca384e5ec4303375473bb7cb9b1d32190c1a1b887a8ddc04a4afbec8aa01385ebf8b07f9ce175f0ff5c68a6bc1aba7bdaef94846e2df1f60d5eae171ff5365cf0a2b7921570141dfba44a3aac6b717f52461c6cd6c2b1e4d7626e5199a06e166965d27256592df82353bcd8970f1ab4b0a13c7c965c59023f26579238d1278d15d7814fb0c8d119be94c1c2b7619b39d0064ab19ddf35d1b94f18ba784429085ce6d14db8951ec687e9c31fa72766a0c35c154748eb3af31222761655200753bd03c5c8eea644535505df784bb5346925005199402b6442c0eac2a4293986029b82c4ee475dae03b101d98053567fcdafffcaee58b4fe554a64d1eeae07f51585ca65004ebb9e53073dedef5b247301e0cd7869364c51d43bad15a7d173add4b51ee8f523f998aef11edc73c9c0b597e39f0357a96d1e7dfd2040de211d0773208906f70fdf542c1263d2f5bc5d47c0371ad4bee1f4938affbec5828f8299686d2c1a9f76ca6a728a77b0a99cb1b84f32fd8e279a144828580f78a15425c4e511e17231be555e29889a77ef9e979d0b9a9e4f8391f973df17deef87f644ea073bc9a34122feb4fb058763fa9e15335c8eb5d99c254fd39157176f3d33c64fdf3d4dbe5081f94075574c46945528e4bbb09808d0c8903f7ba85b1160777ecc82b6a473455948cc005c14354b7e1a40469e589a194f3e4fbdce7049b90bd687ee61f20dbb1230bfa2c223628244542f767628d364302efdf603e6931453a15880ca655ff242bf019fa6d750b78f55fdb9fe8c4d6982a703797c592b4141083d1f8d1e71f647cd38407068feb8a14f3e15c76851cbd5dc50164064d7a00b7ab42b10bda0c7c61d8b1f0853495ca8238891a1783b9a5273e316aa25c4254ffab686030fc3b105c0f60e5081ea5bbfbe96fe38185ef312257258ceed01aac681bcae3008f60eae7b9ec10a3713c750e13d1358d39578228ba06498d281c9a37a027269898e0d2db2c730002c342dfa46f9bd9908057de688f5b3d2aa6a00c39983962c201df7b2893a6f990f503dbd6401dee4db5e0e6e06f760061c925e91931301da4786572afde7077660cd380fa1bea01a55309aaaef2311007eb1cca49d4e32c22ceeb56b28372407c6063239632bb5c7b38591d2ab4ccfa18079ee7123c804fd55ba0c332fe48ef7896f595270e15fcb785f77646eb0de148f6040742cb594194e652f8606990da21ec0b639f3fca3846804d528793f941707e89cf11b78909bb03fd6c653c1036efd145c7dd02ec8034cd25a441ad3fc842ccba936b5a251b12e7806c5075e1e4eb8af7da2ddb59e9e50028d2d4bc649411948bf6b2a45889343097ae3dfab5e0627664cb412a301ef4510ce432fabceec22d8b43b94379b84c591510c0e180c14db761b6434e1bab67d6c4a1100f64bda4c2b2c1ec672a9f84249fc02715ae17674e78d61826f35dd856c5def9658351c774332aa5cc41cfeac199bd563538b97357325e3d54a4c79bae22fc937705d29e0354e29260471522daed5774599d2385c3e9f22be702fe6a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcb0f039186300e8dc28f7c9461cb528858d05d5a8cf861a3f742a25d5d50485932dd70a22a29db22b503d103b8bdc13cbdfd2185f1485045e2661ac0881c5718cc9d4bc71cee3f9d470813fbd9ba88b52746164fa8b7a7d0fbee2aab84175bb92fbda3a867f3f7f740b75136e35ea6595d3654b55d452f90d4297e4a9f5026b67f7ece5d4dc28c5abaeff455607cf8a58e98b23cb566a476f0d76c4ccfe423369136ffe1d5c61fa18849bd6f3b0ae070631378bab159041b3cffd95526df2728e3e53392c59952aab4c2ce5ba8aad3881de0e555d7505e20767aabaac6d3282956a8add23220610463669b18bd479161e8065c2e2705d398044e03a80202342590874792a33bcc1161868a792002995137573e11e9b6a9164bb2f99f13777dd50298953ed013ec0e143037c12fe509ae7a849e99f018e7650fe9c6a9ab70b05613197f99ec43d394edf0a70f8ea2a9ffd116bcae7b62e59b3e95d43816b13010d88eda9843489d0cc0ef4fec41cfbee211dc7d5f27b91552408ef120de568ab1e0301ecce69dc0e00f7eea2930ca321705ccb788fcf9436d2e53c55377e00741192ba4bd299dcc839b4e2828d4b9c74e1140f601c69734cebb9d2919d3db581294be331a2399d494920c719d429da70be47ffe2871215130b06aba113a04c55526d89c3b9c901f262f2b1b4dbb539162e4e7df7218794cf9006960db793b04c87df87079b54fb479a48f9630a666a6032fe1a7d3868fd12762c853ec5d38d7994cb2d85fda554a4a2e6f8733487e9dfdf99dd3a1aab28ecf30d69a5a0dee009fdfe6be5eebe63a1909232dd62f0d34721932dcec12a77a06361e37c981b982e60911e386db1378b30e4d4d1c226c6f04f8321e32ddec60912c2b66544330a2fec79c1cc47717581bd9e69cf3abc81d07d336ae0d0af00c970b3c0aa74830dc4bd6de73ff1263e35ede73b3f71a6b0074beefb5ad9db46a126dd0e07e9a80e490fdf48025e6d1e67c5b5fc6dbf17538169a3b2a5528ec0d02cd4dc50b3c3ecad4c960041d3d939e0a6e41ed9dad62707d9281565b93db72ee4d018fd20c897035995fac337258a28090d0f6217068f818b78da73c9543722d9c0f92e25d00eb6230b6b5b8f69a16530aa90530060c265499195c00985f9229a0c9a2a53c7ee5ac705c1d01af9c601ce18a126b7197f9332fb512b96e1075dbc5ddcc96ef66e2d20dbda739e9d423232ec830c5977087058b4fb68f3114cc57a2cac4cd999cbaad63a1f80da807eb806ae2cddec022bab382dc53ef80d35256f2f58da5f86aec65ce85fb6a54f29a575c2bf290a1eb425169c94434dbf43a9d50e6d045f7d910b8c91226331747988983582bed55d0140d52b150ed7157b07bb4fcfde4ed7d2cc093d3f52b231528bfe5714eb769c0e5987837e21cf35303e73ad114221db2d3f0939755ab0870467c6c9b54901e2eb890790459bf1181789189959bcb784e18b02e352b1d593234e7a5116bf76b9aafe8b5480386365b78d39cd48ec6359879d49837b0acb6e705072695abbea3b4bc43732565895bb6e0db7e759dad1f57f8a95677b4669d4114d0da7403cecd38b279bbf78aa285dfb7ea79ba68e49bdaa47ccdd213c0a17558c1bbd3064530b20d9be2801c6893bd667d80e36f87e48be9ad209ec5254fceaf00187ffd07e89f0f1df90f6f496020a661fca0cb7f8cf85e2ad799e42e3ce32623e01ada5d14b2732d179a51b6e885d93d4b13549810e524c504fe10e59444c9a90cf5ffdd5d03a0e38f7c84da3b703aa6fe6f51032ffab83fac3e5784edba46659bdfa65128d16ccf4ee8c78dd711df07d630aa95bb3e990c03856fa503643b174d15d1a01bb9df7516f38c83c95024bf2e0b3a82442456f8ed7746d4db2035ef92aab98d0c3ca3eefa19973d44afd6b6deef72b5721d93f9b9f9c5236590cd50aa009b5ebf3586c905f221e21f92e08a87b0d5c24c7e9de1105a5cf7f0217f10e7acca09e9f46290163fac7b9cfd7e18ad83852597c6e704e8c73672ace77f90f8413b517fba7d96434b4b8a72048cdf1a4a8c64f1e7f235735fd18717b7072de15dd6335f7ca9c6910144f1e2ff897edfb3c81b80112f90d1e9094247607d2a8637c2f985c851eeac24c51ac371acd77fb73fd09d54bac00809b0d2e36a09c35e9e7b0fe2ce291f572472cf5b0c0bdff284668dd2bb01a3895eddca8d9d41adfd3a67599ed88a6897970582c35145fd6b7e74508c113ca9bbd9d93c1a9f8798905902a9cb6bf645c178e740aef81948d679a29b8c7ee34a0fa748577ed3d644ddfcb631c0b6b7d4e8912fbf6cfcb5d285f2854e870490da66bb8353d2c59bfdedee5db6faf72a2d0866c86e476b597264d3576915f3277fc5b98ddfd16d8b026bdddfe632a647498647f5be208c96e120136622da90992bca9318307b522f5d1d99569defaee963e61e4d2aa9bc6abfef4800f05e03b1c710a469cd90c91a2ac90db4863c31638b3de2bdc32e7cfc9aa6830f5b0ef4538935ff0ba903853e52f34a8c0affb4c0f2292eb529c4c3a601ae02e8ed7ea8414e58ee2e168ccd5b5cb5513ee1a4ac0e29b1eaac97b04fd0cc7aa6a71ea181f261f31399ea682cad8d04b652e2be228b974fec1b1b1c111d81efe7463cf55b6cbbb5a969f4a46c059a9574cef0c9702d57537c167597de5fd488a7f9a93619bc5ca4a31255abdc629644fcf3673d7789bd1837f9cdc89792b32fffdc3ff0b190fc27344319da022935248f2e97b89081e399855740f774b01ee7e334c9e4d81db0fc18c810907d04ffd6f832c974acec165e0738c6b45d5a76127ae3a01946038c8de7f066c37913848cde98e21ee165ec2b1af3ae94287467a570abf854c09e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6edd02a5bcf1404c67444dd3a5914d18b543077bf440dd65e39f34b98b8af4f681b67ca47ed00c94e5c03cf9e8c782005608f74d6ccdeb98043a11ba1a550baea47f4d52835965cf303f9d38e82d38691f98512af87975c863278da6a2e0c8e613486f626dea36a6b7733e09b430c9775209c8872a56993bd6af81deaed26ec8fdabe6e91f876b7cc5b298efd4a02ede423d04f69609d39d3331e6a28972103574692b7ebe57928072da8f45244bc5f6ba79b890d4a3c9148504ace9c497b801e9c8964f9233815ac2434f4ead4203405aeb7a9b8adb6b749f5ff6816b8cf3bfc07e2a47e55657c83e16742dd7e5b02b15bf14cc822221ea2e161b7e4492f3f646b10b4dc90181f657988ef42643e1bd7aa5e0876f5303cc164af0068d0658140c4c46145a63394c62079cd21e8be07b22053dbcc740f0dac1a65c0aaa9bce545580eb7cb3272b5c1092e59a50d06e019a92a9218fa4da2bb8a0dfdfbe2f789291d2929ef498fb9f76466e17aba915480a0597b896c9c6074f934ba2128827a53925d19d35499dee7d6ca5d11e62ca9911a98174a45f6468ca7e0c1f5a26fc94c2c8cf77d127e9209112c873e769c5f155b8cece5ac326dfc4d32522d5eb585b281b3e2a185f9674a6dd8cbac812bee87d92e62d144897b88e60a72927fe2bc0f1b62e0142117b447c0ad5c82cabc555d682ee406cd85fb6eeef7385ddb4fa58127e8cf45c8fc7292da23e9b0e5045f30bd93199ae7ba25c7ac9a1930d1d8a74a5b5bace793dad5e202add36f6a79832d416f6af94e42285234dd41d8938d5a995b538b3354718f46616fc2a3fc9edd4c26e2c39a2de4683e42735b61c8f14252a0a44a305433717fbe9d630ec9e84b84850f56d9ce03caefd406ee20b7253515c49e8adcfce1d80957424527d8ab4e969693f504da8264f789e2edfb43d130ba5f53b6882947703bba8df540e04f84b3cd83a1e8fdb3585d4a529f8aabe46bbc708642b1730bf45f282c577d08d64bbf66c942d0370cdf31fb303793bf367b824cf6ef43820ff4b27d68164d868fb79cdb160135459799184cdc32ba54fe15a13be86c4d09a681ef1ecc087f2b35581e003735b7fca883668112146b5cb7c9d357d7dfc60370dda34b959a84b6f339343b8c5aa5e984c36ea4496b653750e3503b530a4b4effd3de19574c9a7340334c162b455f48c18492be00c18290e2426952af70caeccaa80fb98ca3ce7dc57ba5ed89a8bbfbe7b44f9afd7e6c02cfb922248d68f8990b1e47ad19190250ae0f9414bd8c8ff30ef1c5c5098f13f91686b0565c769299813ba921140855b86e1d0edc7e2c0f970b5df074ffe2e2a0c2733618d6345b683b00e8b40d58d39e2f0083ee032551f89280625b77e54a1eba5e047342b1e230fca2bd6a10d0aeb94d5cffa03f2d49704351adf3ad805f6abb0e30a281e0a82c5f17b6168d68845bde89833570a66db2c931d7b6110f616a9eacb85b910cc904c12db7e41ccba5322574ef5546906e534ca763b3a2c8dad256f2c7866cd94eb9ffd262768b59f02d6909e47859cdb96e5d9f263d06e232c8b514c8edffd3352431dbf30dd6067f4f976dd37aa820498de595a65e03dca669c725e97f43b0c7dfd08431ceb8d138c7e925410e6a3ade1260e9d5310429f6d0d7577fc78194aa14fa8e5514e7ac7f6b8c4c83753051ad024f677929125930a47215dcea37beb30c1061893fc4c7c0f0d004ef22b4782c5dad36874ca667a3847cd8fc4dcab0d4cfba3c90a5b97ac5bfd33bfa16cd2e1b832600ee43e536be6a64b270505be173a6f91e50a47596fd36000e61f32a1358dcbaaa41ae51582036b9a322bd055dfe584751e5ddb81988a2d3b45ac003d9b8b24fad8e824062680f300a2ca5bec532bbcef5b012a156596eafb9ec1e5e13a6a08b58ebefead239b871a2cbce8fbb5a8f57cbc6a0909b93061ce6d298856007b82c1e97f95d43366e35e72cc5cde401e9c736f2c4394caef45d38c538390ea5c63ca2e3233907bd67b056fa9a38c5273118cf23cb4f655f0c3aeb8ed8465141d736fade08d6a501f3f8312069ac2d9e1c6a480525b9ca56aa8f95bf35d03a41f02ce21330fc45d7c5cbd32502dc20e6a0d3ea0164fdfb81f977401e39a5b26c52b41802eb39e4d22fc113573309c8251e04639fe2a4f4ad731db04ff90cee4d66cfc03ba99f5fa71f73c571a07bc84e9e1999adad720dedb57ae551b6b02961b721e27f907441c9fd8767cee81ef533c9fa789841a5a947bb57f24578a9c4345317ca6931a64858f1a4014bf24ea1f426566b8211de7e0d23bcb85e189003e4845deb29ae2287edb67b935909900b80b84b175f752fc1f2067c57c6bab46d111bda218f383ac21c718fd1e7f874457aa65fe7dbeceef5a481917b6d870bc809b02b6d65bbfb38f0f24f04438bde4fe400e2657392ebd1e8d4f258c046ba0e97506d4e7c0a47bafe58742d69bc1bbbed8c98571993370b183498a06433d2d7c14276a7581ccb3b67060af80bcd292f1f0acf0b0f735e7d102c6e429f71cde21d627406f562924567d0ad8f04e0486009a9819f0c59a47f4578f44c285e5f0f906f1fbebb65153f3b1612ed2b71fdbe0451a83feb903c906b890aaa81a3567fa4d5281bfbc5d3f9863c66c26cd09b923284013b7500b20676507bb4205db9d2767eca707336d0a99b4ed6203ead4458ed7aedd4644329abcc41b3f819214f8c5ed0df3d09622ed760444718b97cf0863bade94e2b99ce483158191177a168bb9abfed19672bf45fa07d255cabdb1a727dad9b8c5a2dc6bd33fcb327459c747016c7c813f87047aa0534bdc78f4578c423e1db2ba0c13bfc8beee0990abd19373f7d1ae3d0c116ea9e0ec7c23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h70ff5916c387f73fbf786a78d8c19d31feb410b0f4a7fa3022ba24771fee76ac4d7c29f14541998eb70f0cc86bb6564df0e7da5bbe67badbdb1c07b7fde5fcd2da19fb984b29a0f79eebc31dc8912a113d2e3113134cf86b5e73d956151bcff8ab51bbb26d0e4efd52ccc5c7d8bbf8552b0e6843c6857f0f55aae5683b00eeb72f7c011aa1127322d1bc03d2d70005865358f2cd8b26498facf114e56a6a8fb0cf041d99b245c95eec0ffba6e52f441bcc6a6b80c8864afca85b5220b90c7df33f4771ec8c1c928e9a4dc109235495c269bdfb44d8e41f5a5bb8cc02c01d25bd809b66d519a4376256841bd8dcc2ff5731a0b3b3aa08fb8b00e6abdd576e7eb0bf3f7d0cb92b9d1e5adc52b34a6b1fc79c2b063d98e7bf1d9ec7e3b2410ceab05d8bf3937a1a80cad4ab903e3cc4ea332044e391f5eb84df3390640fc561b291caf4b0adb4534c1a1557132c7017023d0bb882b713e012db11756327dc5911aa0bb05a58f04c01653d24147c64edaa943649720ee0650ec720c610e32c8062f0204d5abcec9b48d684f22d9e8f1e7019d1f60b6d8ac8297773e8960a93f467e197774bf0d63420692cd7cf91eeb5bc99533f154adb4157cadba2dda37e265e9f209f96eeb4f235e8ddf7176aa86111f39b78d0ebda6498c23fc745b70cbe912dd795b5570e112bf89b5bebccd9b8dda19a16cf981f9c0ddefbfed78fd9a6cadc50e51e8ad10a192d4ec2ffb0a116d227af188e005990adc17b59445bf7441b6ea4c3afbc5b117b98a61c351d11dcd977097b062d1cdc4a3d3199bbacedc72e4de0a79bd8bec84179e57013cfc75fb4312fb27e35c9866c6ad7374c72719f5cfd0c7dd31ea120a38c2a992e0baa95d98b9944120c8953d43e532f35f5b5629cb78d08b425ff92e2a42692347c657f74cb892b00187f01c6d2d8a28ccbece9565db7f055afa248b21cbb37633237dd9cc6ae50553237777f3ee1e179a641849816123317625d4ad211d04b219f3e923a0d0f658a46c5763e29a0b01bd6e670d094b5776dd9cde4b65c3787267e652b8bec4bca0db677d6381ed1617b6d5be08bc48dddeef26d68f0d774a27c0f0007e29f0fde76188b967d3b0293d172d650ec00751f1dc1ac917040c1d6239efd7fec81ecbabf9509ba0f2856a94959dcdf91dc941f4a625b45ee2c8d3f78fa84470f4df4df362aaf3c0ce913f6561b8854ef588a3a3ec76d48326fda52994639c779e2c3fedced4e3d70da53fa2f6085f0c3307d1bd3a8219add3bfd6789787cc400da3e67c3de60f4ce8d4f16483557e389234a35aae2ead11a89529a0424b4d78cca8c6b971b875d10eaab94a3a54420a28f32dd430ad9d712f559a9d7816eb17f2d11d4bd9270b951353626fd391d137f259a25c0c268ce348e936b8f4c1798f6190df6fe9a715e4c327586bb9bcaa677b7471ac96567f635e355479bf81d06072a83d759a0a211e456d69513384e8aceae262c4f17f5a3f129759ab256d6674517ddc31abc2880c5d57557cae6d94b7f64ff99887d695f6d9dec94d597738b268684832c66cc3e668a28f2699b9356a4b9a674c0b26ad3c714724fafb2d2f7837bf12e460bd56b9769c67e6ee2bfae50260a48defe1b1d2afe885ffe85f7d420574e74468a5668232a61669d49fe2ae2df0c12c3257539355f184026fd00f763c686785a70cba2a096ec2b03207521b6c0ca2a401710926df9f03e08457a31bcd9dfc947f1e2e7925cf653d4f9dcde2159d432fef9dbb280fbcb2d2e95e66d79476fc702f9c27d4e72a91b46c2d6eb14ac4dc53042fd231c38a4e20920318bf457f28c2f6eb9a75fe62a0f6597e21788c3f6e3ea0886e0c80e09f20b558cb7767002203b1e7eb3a3ab4aafb9c69328beebd13b867bfc6e2ac7a7094a418d4cdd554b65fec8f46b820a202ecf69553b6de9dca07427353b528c45b50a4ed6beabafbca8f551a642dedb77438ff17189b276776cd5737f835608845cd8a322d5a0b8fa32693b7ec8d2e8ce846e944f9db8cf02dfd82ac40a2c390dbbcb2336038999d5a52f31eb7ffaa5b24cfdaebb599e74ecf39c6aa9b8bbc77e211619d77f64426b27c2e6f15638863c7d129c3cdffc4ef598171fb1e70f1617cbb74ae78e67759b5622e1aca22a9d228bd0e8bd836f61feb45ccda4c916e50703703b68d279fb0c9e905c96a7e5bebf28f1feb13bb4376e92a2636091fd931e6e7150ecfab88f5041ef60524c426756b8bc813620d106747192cec6e74e1050ff0ff7ecbf161877ad645dd19f32d2cef615c32f3dba4d37b92aff435e15e7bdc13d5b7b2c94eb1fe2ed8ea721d134365172e90555d9128566f4c8b8a401b2af87ca621a5ff300ccfa38550e39f6484e657c139c5a6678fe31a0d4f983c77b07df79a5efe056dac277efb6b2d67ec36550da78e2e4ef56edd321dbe5c6e1162b8b5ec14c0c851d1c68326911450086e4978546b484230aa756cc25c9e32fa21df9ae11711ce553dcf83e3e51672997564279fc62c20655365093a6d49e01341044ae154452ea2d2e166b1785d169777c88ca5a63bc62b6283abaac008cc3b2365b528291d7f8544e2669dbe72097848902fdf6e6a4bdbc1348e9959e954d1dcf4b8f912358d700174ef236a17f3f96db488d7e95bcf2acbeab76969e0715b494d5fe4f626cf822b9c851be8a56569e6c7d2d7bda053e938aaf9b8a194bb2d251a1f94ed087ac3274e4e60957785241276b5b89479355213551ec3e65f209d1900e10f6fe6cb8c812bcb0bcb23a9cb510ae1b3d2f9136b4387dd45198a56533c4a125b21440203b27c4c737dc6d880e517b375a45a9c105a7acbb0ae90a6165f3f969177b909a2c767f8de3b5f7621e805f3ea00095c990;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2ce2c42dd96b7b9e6a26cfdeaa6b90bc33d2aee703085b075b1da932397b2c40c62df10173e77a69e55aff9240344d39b697908bb7632c2e28737a10fb5a1c20b5380115b46f396c01a71e673e4b2b318776011ca0bc2bd6c72950b05e3cc221aa748fda2eff679cc0403ea0a9f4a6631d5449385f04a794265f296e02a4a5e4191d632637593e59d1ae96ccd51f1bfa9dcc5aaedf11e133e41a76afb9a7f93c9f87542f964791d12b2fc761c3ae5c2e4f95a7b35e5fba415d10e6abf479378bb39766cf3a0df82cbc9d75a3c128083154aff13924121a88ae931af1ef38a1ab9918ea9a40542947161a20f488dfcb182b8e2ef1f539bdb29b0e4d13022cc9788c90f29b9ea3c85479a66e7b94646f6b1b10595d550d664142c186a7f6ca1069ecf066238dae28a2386ab2b346ebd8181f92e913d01776240419d6f91c97c0d57500589cf92edfb5b82dedace30f621a184e1b776dd948a4b49937d9d1f2fc02a7627b76ddb6048032165cb66af6eaa663d5e83c96033a34e647e6bc73d8c3967d01168a75341b69d3b1f7dc573bd17a38502b487eeb658b18e4bfdc901eb5f88f7d577262d4c829c8cccb9f66c4ed546d8532fcfff57b8d8964ad9075d357d5dd9f92ecf5a91fbda2588a995180925958a00373e5366d9d85d764aaa26368cbc207da21e519b3de336b158e1b6367d723737e548097cdae937f0eea81ac904d1667d84e00fe89236230227d178ac8242700042ffc71e39f625bf06883b7672f463ac0c9da2e9da9c5c0bef89949f213fcb4777f2d6f884b7897f58389dc087239ef96be941f4dcfd164607577c83a5291f65164c094ff83038ea361469177a62e3ebfe0fbc9bea7d340463fe3f00b0e6fb124ef507748b15143c7a82dcb5960c32c4d5815d7f573b9394fc994e728f73cc54007c0ce7cf10c0e4a77d4c5cb81d954a9a3c960b67cac8e621241d59aaeac00317dc33f855a8f20fd23aa37c176e170be39a69c7dbba1c09e0077294e903e18fa1c70bc1f60c91a3c2d4f07c71f178052edb5452bc27a1f883f9dc210657fc6bc100fee1055eda49f899239f476e28d23fc43dd76d82ebe50aea1a0885372d6b9fa954dcb414a423c380125bb21e2ced1d99fdf6ca98b0e52771f0f9aab48bb137aa18caaa8f3c14f0eaee871d67fbc8dc8d8a573372387268e11665ee93dcdaddf2d6abf703e75ba576fdba1c41f1b029d534273b1fc3bfc72e412327fbb888df10ed42e2a80cae20622fc9ae99db6b539bda63a1e3fc6bb949e2a7d49466ce197a52f12ae9fba4048a3daecc0b2a52486241cabdbf4b08183a00c945031e720a470d9740e204fc806f7780f7249e9b23b8b242595a11dade5eeea70ee397cdcc0c6d6de7ac3e00f8f4689af04b27f7a0aa71579f5740ae660f03730c2c827416ea74642726ddc503ad35d3deb5705394dbddb90ab9816dc9665995aa2459f399cf1eef53e95a84249fd7ee15d3f83ec86aa1e8cbc9d66c8f5027374c546cbedb685af820f2e5a2949b36e669b03454b60a4248eb5c03d964941f8411c6c336a816a902a6c11e389f4828c86931e7aeaaa8daeba280847557ee55a1833ec3f274f33604963cb4a3e90304a965228b650cb605d3a10c816b3087bba64b9c520d2c542151c6cbf4099a30c56b9bb507959f48b8d960d1f7d3af17ab3ff4b2c6c693545a564834de98c70915509d2d4d3c06058ab91876e2e4caff294105769fdf0beeac67510c015bf5e20e37d8494ea82cccd1048507125c4ba59cd88e265524a6359d343d58e8fe17879d98a60e2266a5779784f043e4a77a78fb1368730c47299fc825119eb2bc86aee67750975397457ec2bae7c04b253ab6ddb3b60700833098767af9c54d172176ea32d9f7ee0a2eff1f8eafec20a3ab7e381e02ef42dd8b0a241eeeff6ad291a89fbca0ce9aa7d690e407384768084907167c819b5ef7f47740544e3f0a11422360e0354791a22770f65f92db4567ec000e7a893bae1ba0957ce4d6cd2b19b7f6d13a0888a1fd8ba352a19c95419760a5df99b0b08ab0e404be90602ec8392cd6c641c0243070aeb13c8292372cd69c868be872685ed22a6697bc51149e65216507a7877ed36a36236d3390112ed805f3377edab41821e13c3f7becb190e9f31e25f997e5269159e978d91483a1cc9831a9aac073d124fc42959a9c1a6b7d97b58f6363aaf38bd39c9037ff38ebf2293e6d4a45d7c99ada4dbadfec18dfac2ae1cf8f0fd929811472db4faf66e8c761b5a0bb3a622c488360951141c2db2ce9c0f2eeac633b1c3ec6174dc459f17b71d2ef9f4094c7672a57c003ccfae8de462cb42eb80e565a97e36fbe84c0f2b570231078c8ce5d5c372103037cc82b5d8506a099941dd0e8c66ee003a8d6d0fcd5533382d89fb19c01ba9b7ef65b1e6a1530f77adfb0e0df2f9c1ed32594e49ca0403047f83c3ab8dbefbb3b87bb50c506f34cdbfd94cb92ffa4dd5f796915befbffb34e28f646611e7f0edf96db9b88d173f6dca30f967647abff4b884419ba1492a1edd84828cb9c72925a633175273c5b84d23c68210b7992431905d522e84a3592ca11d38241c541c61b69530766542165bc1e3537fd3ae4aaf7ec02c69cc46963eaf56e3685612fe8e79a7b4d7390750e45a68a6175a76bda67242168620e6be2a301a49d00254053758aa86e3bfef8bcccbff8fefdcca2cd95910ee9bd79d14abbdf098e221890626ce52f2c6f3c065027ef640fdc2c25c8ebe9037b85cdf796e80ab1b223ea2a55930945190e13b5b6706e47be2cc9c6545993330b9657239cd85dc76f09f7b815b37e0db0b39366cb3c6bafdee9d9e30ecf14454dcdfe396057fb6803cbdbfc2147e9df9de6b1e0d616f4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4ffcff474b9b7c11df8e33aa8ebea71455cea2288e8c8b7a7d2d7999e0b88e6f6a1c9d880f7e48db3db98d73e3ff6859353aefe43a701729dda99aa0bc67e483f7560b32c531e36a5b872bd3d8bd4a76e5871c1263921cdaa832076d558c6f55578fb73963f8c7745a9e39332b91a3253ed20f7171b2bb965fe370175b7773976c478a27c427ff66747fcab2a8a2e43e56df1217d727df4c7a2b22916dbc33b8fec27fddcfbf99761042eef533a2c810c23364b6d626b3e5ce4c47b264f2cff87ab8389ab940b2c5237da2076f464f2168c4331b5e9863b05d7d336974836a672a3bc8ec2336fc7f21f570e1386773df7b912224b7fb2dec72cf688356a46a80c8dbf702892fbb16165ec669adca503c6e8ba12ea150d80c76df9e410c7269d5d72db88d102a578513270bab48fe307828026c4534180f2bd4a0f5dac1b391295658272fc90c1d210027fcee01c5366b8d95be2f9fa1b4bb2b2a3492dbb8bfd8e28ed6645802888f9763188afa2994a3258f587be00dd74cc09715a12038804b5abd58ff1789227fb6d8f5113965c47bab4bf6ee90a79f4d4d6f663d8934baad6c18234d832cbd0975c89f2bf9e5d315d4311d7fa33df383137eb3d8ba44c914f993a347afb4f744b63635ca4373bec9616d5d8f6d4fc9816d4e8d99eb87f48f17bcb2e1593e875953d67efa9a84af1e1981278d6ebd95724ab0048aeb7942a3b41215b9b7d2e8522c0842dcde6eee07fa31685f11b89bbd6a74acd83ddd229ed33e878928039d060429d6717fe12b655eb12650075baf3d269773c024d12fd06401bea743931958bbc0b925cd427181b1a655203f3e94e641bb369389e2336df41e61fb8d4d026e105ed575eba1484abfd2cb67b03ebb75c2cbae5a54f11da981e18657591dae65dc2fc37b96433f40a1f3dc186ecdbd9da8f2ac14b08b65e92e86eb68cbf0670e0814f3e5c7b28ade95c82397f603a489a2e3a2688f8f642e4f5e6cce81685f2b37916918fb4951c96391b472449b4ff5a2b48f8c3c49b8ea0712089d41f47adea1a9884b6c6096f72308bb22213bd8d569f9f45d8551cc0a238410cc2f722fb59bc1eadabe56b6442d430be17d364530f4a9d73bd8d0bfdb8ec0883dbf6c10f66d7bf5b4295f382eeba118e3c350c69a70bcdb2765b085d72f2005150f436445aa6a184d452203c8096b55f7faba6394185f1667f8a8877402c8574d746f633abf2099693acc4491ede7db715f11dc1341ea8c97e0331d5ed0cda79358851af6a6793cd4e644c28da6c0ea57cf81a5ac240709115b93d178ddef25b742b6dd5b651064242c95ae4c5083cbcd52304bc1816591b3d7080ec2de08ff7053b022622f69a30c9ae97d4e0a8e81162c6b8d03ad6d568cfd26ce4b479c02bafb4699cefceeab8c0efabdd2715cc5f57bfdfd4194fb44a702b7f2e5f53640d78170a25342f325373ec702d4a44506756403138f2107423380e3d1c784f3b0691a5c64402bb52c693e42abf5b4af3433ff3363975673240e4475b0d901a2e37dd2cebfd363f59c26ad9d98af93e6c0acd6023018d0c34c0a9e21ffa1078757d92340c6fdb09198cba834449c2dc5f9d29997b9cbf069df879f5853ce9c57f6aaaad86ef84cb6f38e398669a9077de4f638d7b7b968994e6656d03d4965981413bc0867f060ead7ddff728d6fc5f36855517984b32ba77a6e7f0e4b93c2644c7e3654119e60b5d93f09058fc1f38312b75a361205ec6297d5aa48fa187c9a25e122b8159119607ce7f38a3838c725ffbb83fe31981c115d02173a94c5bebf831dcc4fc33d6abec34f54309f234eee001030e06105276224f5bd535d9ff42d527e9f90aad43af6118115729772ad2767122d06aa3c36ccab2fd599a1ab7de2bd49185151131249b01801d424051f305287b540693d48ea1e1d2b372c6bd53f0f75bcde15b23524d2dcce170b91f4b916ea09dfc5afe6000118850d8270f8cdda07d5e4a071dd0bf723e198c5918357d5255ac4bf0f35f1824ee5701097cb52ddad1e0008032f6d0015ff0e3bb7941c44d2f0349035bf77bf582dd9caf25c3cfb0a8dd24c2b4d804895037326d45932d66e4d7133cf7528d535cfece6725d4c89d14e0568882129d9f4b81dfce3f708737eb9665708cec5eb87f475121134831436ac1d4aed77879dc6edbe4ca60e308e8e69bb078642d3e1f3868c1764def634ebf15a43f8e86c8efd38739c5ac59a3b8c6c9ed15d6d9f9c347d2acbd8b43fddf462e9d9031ddcfbeef53154f444e733686f296bc5503ecbd79db47f74ea896c9a6d358ceafcf6c3b84ece7d13f493f6198f6888c70560ba0993fd4008feb346040d0100bdf974c43ff11aab6e4fb3e086af829d29238a1ba56dc5795210027484d24d3ba21b01e0bf05bc198f54b8fdddc1d3f0e5485f8dad27fa0e0529b8372820d88b65c7769abf24bbf25e9b555b82a903d131a85591f1215e9be92ea571af2380da8d9a67849b834a73346f6d33fbfdb25901a434f414e947f2da8baea9fed7bcde4745a4171014ed4dca9b9649a096e1ced04ab0a2f00052eba9b40266abf04d821e87d63896b39db83381b50522d99add0ed9377b67767a17a2dbac46cf6598d9db8560ce29148d8c1daacfdbdf1e7a9d1035c343b7d7871fb71d55a8d04c867da70536d9c0a31d6dfaff54342c20464cf84087a4cce0491136f0a9f1a722fb22db6a775ea90f6326bd011ee5059c2d425c560d5a4eb96fc74231ee2830754356c5e22a825beec1b312cc748af75cd554669119c27070c8fe58b9ea0a537f6c15b0316967051b5c20b27df6c9e0825fb087fc1b5e5b3dd9c9a1385283d5b07d812c9c57be7e2b86447b16e2fa563b48ec8617d4543488171d38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h506b242ea28b96d7a1791911ece984da290e5e41392819b44fe1697192e3b471b0fe7cdf0dd6beb0de2b2d051475c207549202a08c22bcdea1eea4020444a754c62adc3455439838a34243d54272fe13f84a72a60022190b0da5962be57392c3e95a8349e66d4d9a62a99f8088d4e272fa5fb9f6fcebb1ec127b87ccd6cd8cb89717f1792ef96ca04b1cfd1a7ef4e97d5296c532a77966d928e63eaefda6ed1e7dc71e9b290c6d6708e4c471ac259d96405f08d3de7a3bc21d57687194ae3a9248de60da4a2f43dd3eaa6c69962bb88aa8e9cfc14781592a987dcb64ba7845ef09b63af554b05fa3c19c2392ea5fbda3c32027728c828119b42afd4a96b6da8f520be1af81a3ce10c4b8d136c0de84e1bf46726cd155aba012bcaf8ec2461bc7fd564a6a867954aa942a5465c738b266e656232d8ae5fc1da1a2da7a21351567df36e5d5f42dd6f45e704b68c18719faa82b50312ab090ba7ea976ebe3f1e44cb36f64f8fbb25f8268f05f80e1e8b7231025e19b4b22160dec3b1be0c19912423159f03e317baaa043e08bb92e3b760205dff3f4105263434a4bc5ea46b19b080f6441fb40a4bca6d930138d1f26fff4ed1f2bfd19758bd8cee3a68073e4707b323232785bf11ed62bbd6440dfc9f5905e9f41cd1f9d0adbd7779dffd5146bfff9f6916803ba86610caeee471f5befb7d6cae7ebfd65b8467a350e228f5ff6af746b202917c7d07fff865187925a32a18d27fdea1ef1bbceada75056492205c3fa71c159ea5c7a2b2beb188fc38a6da87c2d4dc6e53b40a9789924b62af67967ac8ee08eb2f88191bded17f20438ad2fe9c0b99136a639af958e047df7dd1fc4dbd955c391a8edf91059082141865eef24db9cc9edb97620b9a0457349716ed98f118c55cc28f2a89568564b692484f5ae11ace35c9ef9740f9d8a03c7b8bcb81d5503948502332ffd3e7c1b51aac16845b3bf119cc074df59c26e639114084659b072fabae0519cdb8742fbb9c0ab03f3a8a0a4470a448bd20470196f091366dd201639c7a8b9ba5a86474409e294eff243855b54ae215e43bdb4a1584b6845555011e94d8d2cf5b11b7dd2088b053097a9c38c9acb0ab5d53f4f042e4d1b7c55a2dfc6c7d148ccaa692b85d697b2d26a6ae8863146c003a32d1d9f1074fa881febfaa01913d0fb7d7dac0069e02d0def4165b31de84c74bc8973012edb2a1174363dc69319d9abecb577178863a98dd14e0144888f35af14cfac39d641b9490d38abf24860bd818cab9bfb2425037efc2f66b5f842a90e44be1d92f8c657d0fdb90f93027aadfd3b8843c28a8109a5dd79a1653d9c0fef1f07cdd00a25d4830eb8402e1a07434e1082a5026733f6e19e6ffec45d7bb80c2b52ef0806291c512205cd057cc135dba87e4fe04f59c0ab59a1acddeed7b4bc7e3455c9bfb0eab9f0a9f8bbb4899ec711aa72d414df55f93aa8c3c6035d7519ab8a35fc19e41c0da1f3871ac3bf489c858bd6c18ebfac7b59601cb6bb44fbe710964f641d1ffafb9d5d6f9326f5c559a45d219359be46bfe778e982652b805e4e508f4cd74a3611bf890b09f2aae7aaefe05f57b4f88bfb18906dc7d24f4742f1c3ed3d1cb5c52e7e2279e108701d27cb0d6125f67bec92a8dd36e9f60e531edbf3149b9b3c21453e209679b82b76e0516251ee3da394ce7d41cd98bd352ecebdb09155042d36aa969ee434bca12983b27cdd38dc3fef8f94fa6dee4aa16b0a05ae0284e7b1ad42591594fb5633259c86e5ed77d41dac6c3d91733d439341debfd203328cc5dc1f8b11837dee247febd9d7abbffb37e1212b723bf670c04016a9b87421289821471ee49ce743d0f05331ad319b20580b45200878ebdfbeb158d50c8f67ae87680b84498106ce3f83fa8da42a89dc445ed34924dc4a60c3d74f577b915e8e7c7a99458024d244d1546c3dfd8be36c793003b769f8d26ae84fb056cfe6a9efcf5a53f788c5404070634c584c9d8d508189662bde57b01fc4316e9e6cde222153e255d43d8cce5f65607c0aabf26ddab022422f3773709ca79cfb84d44a307908de5db4ed12ea8ceac8b22d4de4d6e1d8d21ea11b6c4daa90486095f1e99a99ceaadeadc935cff1a7d3c56ba86917e91b35831893bfc16a95ab78a34297bc16aff75fa0290e36baee5865ae2ecde3ccd460ed0f0b6382158bb7f078e99d362b388e4dc4dfa3c905c3cffee59207b7ffe28ba45e30c1b76c61ff5078be50320cba6ee4b87b9bb0e8e766f2680c9057660e1cd240c784505dee13379d6244c51a2be25581fee39bf99ae02aa66e49b0717c870eece7ba5703552aca5880984e7bed99039b4c92763f59ba0545696b728b7a9fe0e99e3bd904527733ba6cd205d08f764c6e5b9151eb29e26a2d71ecbea318a54e03b531103b58d623239ceccfb8a5ecaa6be8350c225e1333ea52b572382f8a9b89e109cbb8f467bbbba13d43f09476b6b1830bb90781c99fa433863ce78bb3b6a4d7a8b4a0acaeeb18125240ffba4867694098021d923c831ee073d69e43f9627fa56b566ee6de300a4cc2a7fc539c6fd33378a3cef1b02de96f48ccf680f7c7f68fff5a26460065d84d01141d636ea02c8f47e8d6601b6b32464d77a18e53afcd621e879946ad20017630bdd6d5e1d3b27775bd997d457bb883dfedc9937cf96e13754a93e69fb38ba463dcdbf3ad67ded5a786910f0badb41367049204fc5b1064363e659f389b0e6ec47349c07aef25fb3afd11e373f78ba7795d0500f7d92ace8d0dd5e8785116bf57bf562e4f7396dcf5bae93d7b501fb567f0f840974f21cc121125441d97d54f78bfe5ddd5b1734cee63d2b57b3ddd25c27e3c09a28a648dc880c1c1d5bdc82117d32bff02ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha46c099668b1ec1db194d678e4b96020042931c6ae7f91b5ae8a83c7e45ed046703a497d9056e97a7c77df0042e47014b8e93aec474f62169a624526499327be9a7d6271a26512e0a0af2bbb17c824b5475758fa44e5dd9ace88d00f8dbe871c6d295090506f01e606398979fdc1627791598359df4c55a606da4ae0f417bace85cb432ba97480cd95525d2cdee649cd68efc08ddd9bf4efa0e8093c8467fe2d008818c6d2317748d06ea523327ccfb3bc6395bc80c8a1b07c6ee87afd27d09b238251eff557abd36876861ea4b12a815814a20c726d409921a6ebf3700c14a482396d3122d5cc3be447b971bdf7d15f800b4c532f74a874df4c21b8990e8089b6645c0a7147e81d684327e97534e38879b169e58080ccbd744c5d2f0a55f652acf16b08f8cb11d210ef7f8ebbd0559b2944560c4d2c94c21832aba9e7b5269e9160a4fba04e96cb2b655c41047a0a45e121155e39003f14a4277d468d5c8fe042a8dccf8a1761378e67fb853aec1c920f006679e2bcde36e76820c411e704624083474483db0f846ec7b20c3efdefea4446990bd3cbcfe385163cdf5e036c0f9950c9ad1f6b093bc9da89c8916c29126476768fd1c850735b309b6770c86ae9cc0122e2cb597ec21bfca9785d9f6056e9b6c0274c967e8576828d8fd4429d7f085bbdff54f43994b0c68f3aea7e5d4cf03660ae4b06fed0eb5599b9b31bbae2ef0d851d9af4d709fe704f2cc644db0cad512c82d800d42c88d7e8deeec84a12fefd5c5abdb4e6582d9ddbbc0daf77a2341a530f8f55062ffd492d483f3ffa08c1c5ac766318d3789ab0c2a83f46a171c3e2a4b811ff6328588bd934bcd3a7c5318bb85ff6fe81ecea370f5c1e0054bd9cb1934d9dd1c38dc81893b5f6f1bfc8c1f4302ef718473ffd767fa061a1af43ca1800efbf15fe44bfd6a2f4887a280ae8263a72bac5833e0f5cf72d79f8a782df6599cf56333c1d95fdee84ef8dba7a62bde7b806bbdd07d413a3e1cb475145c3adc9b2493437f93db0137d1befe679db5ae83ef58fa92a19094c3d6784a3bbebcac6954f5d99d0ddaa6b77e250925964d9b8096f2ba1fd77a5589762081ba4546ce36f7e6dd6cd0928c48abb151e26b41b715db0774138484c4df6af39759ba7fb458d1d02133d39941a96a21545e18ef36b4c9d028774cf0c297429318e019d45110f765252822ab2e17f61423a2ae38ab48d3971c397723a859a6699243ee7b4b79a66fc43604317ab0caad337a2e95273e6a2da9112f889a75b4c2efbe838e0a50af1ecf8b5d55dc0cdd5818a23b8398fe89b292337efe52e46c0f45545d81de764630c12008083669448add903d43c82573868d5ad24d89aa9a25566a456cf4a2dc0295818a2b685881817daf6cc7df0e73f3cc9a857b6d3734a6ff0fb8a3769b0d94e95e560310e2af31169713add50e70156191c7e77345a1ba9b258e73589e3bf0888f64153cb352214565939c521593f7c87772b4daab98adc6d4ed737bf5e62ffc2a16154a2fe8097c28502d499d0260f255b5705e5cb29939505e744ce5cf622e9da351884fb5a8f35bee8d420e3df315e25c04efe5b118b81ec90c3846e16a3ad7ce41ceb4dcbcbbf53f754712395e70a96de2683be930b79913bf2119b0b6eb64cb220b2a84c3c3fd308747507fb2149d1e49dfe0393dbe278f23f3b348d778c1936cc3f8c56faeded22fabe7d320a1a43fea479848881db98dc7605165b20ac7333552e90c05b66a0bfa439ea55ea7b5e0629ad686ac1fc114742b245cf223e6ec0c74999a5cfa440880103f61e82d3cb4d514d62fb7e5cab1978702df5abe2285836fa6e53c8a4505ffa5f0564aa0c8e67a18a6b0853e5eb85653d7ffacab5a3989ed6f02f34915a7ad9a308eb77245578dd820270886fac71fdfc24b2c1aa771bd2223c1e87b83ad0dde8526017b1ef9169a70e6fe6ec58ea00d1598206774c20d184a7cdaa1e0a2906bcbc6dfef6df0ad7f4b6d586cbc1edb84531c1399691f1082d8ce6a44bb3ff8b6ad50333ceaf271344d8155d8751705096f54a8034b3e17fbab6d06a0d70b4129d3524835e3586ab5c37e79898925bd9fcd3abc079114df688c7cf509e0a896429f4ae77136027da768b4c0fd0b87d05a7e0314416c8db98a1546a85dd111a0d19160268da66c34d3d0e611559d492c584dfaf5d7fcf6de0041cd390e318e22d10d936d61e9ef4aeeb20181d0c129816e6b9653a7367b053079da2ad85d1ec2c39d8ee38fcb538b90b12297259526e8012cc22c4b2ddd3ff6ae9aa79d52d8612a45d90426a3daa87dede7a43e0799bfe67e3ef6ca949f0ff1b7f817b86021707cc93a924404b7941fda651c1c0e691f053bcc619cd0c8e1ba190488298e39083748779645d328a17ee266a7ca600ffc600743c4f6869c751f53dd458554dd6c87045410fa8611673f6df3250d92c00317763db6ee381e35ac77b5524c84ce37ff8ce10fb9c32b6ee22fab0f850e87d41e08c3805e1fbd488c91cd00858886bd93771d61696bfb69b5c14650e0a6399c899a9dbbd4eef97809f4183e608cf36f4c9abc09b093ea6242523834e27765fa11c340c362ae132af4cb7020c71cfe9b8f5d1e6311630e2ef763bac59694f5540ff422f76f4e68c1f940e7674bc22f60d8eb7e1ee2dbe71bd4a0d7af5c24d3eca445776fcc32722d1ecfd2872b63531c52bb8403493b8906ba890ce558f33fa93b549b69988db7b3b0afe137d430093e681bd1d18c5ea23607423e8e11568a661599c897c3d111f2777921eae0d554458cb4413d1960c0a1cd3fac7406c6effcba012219386432e709e852d9025028e326d7f16fbef35e64e5006e2df982191b80a78e64be8ac65c9393ec1e29f1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcb19330ec7216367a9f44ccdc0530767fec27a974a8e47b55cfe5d1dd69f62cd4ea2c712d03503a050937a6589eafe22e77282b361b6eb9d9323dcada5e65df83168fb1c57c24670daac3afa9fdc63754be7bd8d16364d7413d1f27006fbcd9dc1017c6279a05be6371e641d9519c9a18055612246424f7de9572057b089f706ff620de55ad7f51cf85f38d055d9fc0b9791d6c851799016b124f2db1bb599b19b9f586d6d7aa0d9c98744612aa3ee9fe39246181b652a1a07069ca98c0df4a20e7445a302031f3f4303a0a6022b996392bd9d9d181e4c062417da512885daa8a3e2c236d13cdff88864a66ba65c060ad54498c9636bc3f49dc3f381857b01fa6130c14f5211f7f3a690e7f0ecb6d5fc669f42ccc9518c08f87e6547a35c803ee8b4b8bf3164ad90e9986ab50168db5ec04cff5c59f49fe0b0de8cad03ff1d3a4ae8359f774636213c02d9e7699bea87bcae1b2cd09c30486f49754e8aa8951dbdbd9246f376cce24ea55500d8a400693105ea179feeea949f2202e178e28ccb4ecfc75b94b7b7b14e038759c9626098629b65d4386e8f9acab5a5a5948639c6140ebde778e69305359543e27750ad592c3eca37a9a8ea73f97251cfee9a6003991c3fb5c8361b8c9ad3f29328faac377dfc024494489cd305ddffd7c424bc7d8fca13d3169e9278554d507811325a8f6fe790159f7804dceddae92d84d6690271dc512782f54a55d9475856604409b7b1b71cdf6b7451f4f02f9034bcba8229550d23f347fe281b22648d270bd6715ea5209a13e53d91ca02f26024a00e2fa39846994c8feaa3a38fc216f57a5b32a11721f8eedc694a8e4a43f2483c6ca2d3e43a02317c833eed3571117b8306a2f3c5775df4f15fb7f26d9fd70ddf942ed968d741cd77f6ccc9b29521873509226e3da317dfd2a5162b49542b29f3ebc331927369cfabe5f75f8af04c0e4430fed1888b694441059da76b9673019cd20fcdcba03ecb73e06f0fcfa073b35033bbd9c18739450e7624459b2e9df83c8bb22b4411dfa83e93408de204028e21fadcd8b8a11a5a83432414628031c5e62a2fd5525f253d3cc43048171c54f2a19e85226999cee571cd7858eb4bac9235b8ddccc8d1aac10463c15d987d5adba32fb1cb20dc9f17f15b9811572a4f69a315bbbcaf212d5cd9b9ae757f4ef1b3c91dd386e33b6df67c6f02907cc17547d00d0193beafe0c17d986aae316b369e47dc4c5d275aee39ccc30efd60573c59599d3dadd8e6ff6fa524ede8b63e2eb26e54c10196a68de20d1340cc60e08c415d7f447be75a6e514140e29eda763f274a8d728752789b8d363ce47a68b2d86007e98bd01fea466a515d1fea5ec33179887488a44ce682ab3a7de821e9a36b30aaf391906e0b23752f0c0b2cb1ca98475eb0a63bf4e42867c7c665d03becebc698c79bab0425f5c0a7d03cb2d757008c6c1571fc249141ae30513059461af0a446f891907ed731e4b4e27cc3f68f6494fcb236e4ba9d4d18e2686c8d39bd55f8232db89fddf78a2977f9b7afe96ed68f103c5e289bc9303e3ca58ba647067c5d0a2c53ce3f2923d73c9c284e941f5d0ef62424cec486da9c8a3c4f491275bc07c2aedbce41173fdc6c161d7f2b5b2fb35090741ad5d3528f69a94e7593e6f975941fac5e53577e432e8ed81700640263377aa504635369dca420fbe68d88d74b128f531315cf100a7c472d3188b50e62b2b200c7426d7f4db51b46fed3f134c67f21d4f0c5d97d0abed5f25adde931e689b6196d7b946e6b0a66deddd08308fb6f188b22577d42daf18e46fa4761611c8d61e109cd319b2bee43e278cb4e3d09ebe59259db50917a2acdc65d88705cf098166a8127145c0d08a3335893ba22460c1b1efde4d203e146df04dfc69352ae358a4c7de890d8aea50b60756c935db66986b7a68812223d64c3fe89a693f7375b20b8a49b2c1e75479728f4e383b99d04ef9881e181a0974023876b95adadb44fa705aa2d061974517575f6c92703f4ba01c774c4c724095638a6b77f6fd71c6ee512dbbfbc31fb3a5e16d573b6e0fc36a12d753b259a35b26e84dde3740326e81707cb505773d6d8bab8033ff58a67c8f10b39737642d935b03c238dc59023d7a64e6fa0a6138a9699e615e33503e2fa2e4fde8f0fd3daee5de33d2d1cfaf455371b2002aadd877553f0cdf7b0b0accc59d324abdebf853e78d92d500e9561c06fa19fd4a0c909887aa10e3305dae1a71615874486eac98a855ba34014d996e1de4df1f78fc08492f2aa55f9235faa1bf6ad4bfc35c2bc019b186fc86e05d0e2bc645a49b27e2bb4fdbd749bf1f8dfffdea117d96ff058ad7bcd26103a94f3116c012eeec8996b783ed1d26433af693a5505095f8be3155ba0b96d78f14a4ac46a098db0ab6ab47e609dd44049b700729a657764b4933320919344f77fc1f5887725140737e6c631a4da3ba1234e35c6ccc6103cd2ebccb03941802dbd5497c45eb08cde2c32920060026179a7f558e2c2565ec3a0765372aebf74ebd9e5bd9774812058664f7add92524f62c2b82900689e4262a9d62c1872568872c9487c2f037e23095abedc46a41a28c954fe041c7ec9ef46c81e9e013b36e76853ea988cc4a028a89dba63dccd57c4389e6f07866d6bc81c34b6e3893879f99b225b4b15619181c00a0d600055a63280cb4e546b6d3942a49668ce4cc6ab3c094c5d490285f815392f5f38bd75bb1570466d6bf7e45bb421b839999c42cf2951bf30b8416dca1ecb8a953f551e00e62c2683ff3760f9d026b3f0a6a5a273a67ea1a6f03ef040f89d20d788ecd0c823f398e3f65348d1b02b136ac3a69a58c4e101124030d2769b44c6f5ef9bd00b1d9d975f7750a66118;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8b9732c1ae7d16a4eec2a53244a1939973a2aa81b77d9cb4edf9522152766cb2f3579563279715257c119b9b6fcfe17d7a1b28f3eff4272e813e6b324ed22815cb4ad047263bc3828726c7c6983bd9fda031ebabce24a48e30b1ab832e7505dbda96eb801658f68cbf7a4735710b14cec60afec473bee2fcf02c66c150b359ed601951f0d7f185ad193877ba64c6ef9dcdc618611aad8b3584932a1fce5a0ad905f2fe62d59027faab1ccace4034313f5a22381580739719f42d2ea37b96cc358389fabe989826abc40f8d1c99bf7a2e4a970b53d3abc9e9324792e6ffd450b96b6ec3ff3325549dd1f4643fbea84547699ca0351a94f4f7b8730eeba1c6a27d10743542bdeb3b5613b3f65274af61e574b90ea0f81cdb303476b7b41d8684324469c8aeae06beb565d30afc712266656e4fb50b5941ef5876fc9453190051dc1dbb5ddb1045d0f836b1c6ef08b561b28380d5204b9a3d52a4c3ab6500624b6f99ebb7c5b5fde1fed18e901bbc983c7b8649882ea3fd6a4334758f5958429b1b8d36576004d3ab0e590e1a470b1af6d052328c27e7311e973e15afcdbf023302dd32cb823d4de5340d28a5882a171f60ab6dc2f2b647c9c8be3e3e7b55832134380e8b9be44c3131325ceab430231e6e118ffd430912362ceebf72a6028085ddb41f694f6e541b50fcf01c95ffd2ffedcedc9d2334150fd751a6d9b2b22cb5c920fa34c206b93112a4e42bf035861c0655fb2603ad2f9dba1e5cd65c29f5828b9fae33f14903b1ecbced2aea0822a50b6394d91a414da6d5cf6cbe71211978e48a8b918921d7bd84444b906fb150e145cba436139c358bc0f9b6c36a3ad3e963ac13e03738c4aedf549a270019e02694ac01a17a84dbac7331d4bd47ea178f7ab429f4b1f6b9eb91b9af1f05f87589f3a6962972248788763ae75ae335cec1697d67d39087c4b1d7826a156e3cf722dd28c84b97c642a72d22f07c4b8dbada33de1245d17e7877eac2087adc644979b767ae9cdc921b48b4c47b749f53e187339da93d3d862355f2159faef5d5340f6391b18c4f7adf10781d59c24ee0a1f887611e3229ae2b281c304e91b8d78888dd915cdffab3f14ed4c3c6fa0411726158b16bb877e664e9e8562a79fc58a0fe956d4f4edb300264a5eb65d01a824b7d29ad8fbdc109585c8ba37495f66a3f64544f09c3b418d782b998357e7ca45b6dea7e58711fc7b092a3aad4f11b600e5f0b150ab8bbce634814f6a138baf5d0d6cbbc66030e9fc85496e445128129d479cc4f0d3775420c3261f67fa460e39eb36d721801d7be0a300a4014fc79af36ca18741d1ee5ffe06f6b9f477179ad84f63b237d447124a60d8128dd7065107015f9f0ffc3349b2062b90e659b6fe88b4433fc777d44d39654286d01d869f40be0910c6c6b5617fcb5e56edc0d99490268af96dca0987032a9ba08395de9f74f8ccd0a1c8d672af29a5e182795e6c4b7cc1997d60d928dc84d1624e8c8e8e29bd24060f9e3c865df7d8b8b61dc8ddae2e7d0bfe16de407ebba7006dfee04485eac02335c5ce034043d45f63666a6b59a9da7a2b8a45b8bf33f68490fa2058e4e19f7bd597958e9223f305767d2cc337190f9d6ad1fa97dfe6b39ead426b278f02fcde3e4279ae27662a6b02e1824e1ce4a8bf935f15ab93a9466e5fe04fc9be1aaeef50aef9aeb0099563b29f5aa20cb8b5ebb4e4a954d029cde22a53c11383d69a09f023c3d58f27317979727f70097c9919dbbb4d6216939085a698b80b119e37fefdca764efe657d64712f40d92704c16ef4b3d1718b90f0b44d3fc2d8484b9c51b7ecc355cbb0da4816f9cbc708e3fda7319113dbebc3c3919b7eb43fdcf76b8486e8b72efb98d95153054c5af98171031b73a38a70a38f7729195a0b1f8d15746993afe95ea7fb5eb41875aada799740c10af395d06f61f1d9fd2097533f9ee04a5601663b652956549d52fa0a1edb67a8dad02e2e7b24461d85688f1b0dee68920615490ab7c34a0fcd17c183a791080e997bd2a1233aa5dd5def31d9850449ba532ee4f90a2f1262a6a1a6369e7ad74a7abefef84a97597d23216ec6a411fb1ee25ae6073d135b422c67c1016bf1a58d35ac0ae368cde3d7da7cc8c523c0de1b385fdecdaaee54ab6de1481cbe83b07b7ed96000e22cb85774abc4ca12e11f19cfd2eb8574b4c46a563f10844b083aa334315edadba9fb37b281d63506045d5cfb203d7f9db8fc8ba2ad1432d3eb800b5d245cc9ace996c47b3d3b58f90fa5006a4c2b73b4d40864666f0d3df0569d9532480ca94255c5c332a9390d647c6b47e69694bad7c85f1c71b33799da0d2c593283862604ec4d5625547c329beffea69c0b766a3ce6e934be67054a400d7da9b99812fbe7c47d44588f0a7ec377c1510e908981f280811488d16b6fc8a717e75a562532eab3907a4618c0342bf26d819ea382c4195b8ce5717499c63a9d27481f7b499411eab187a58ae460917810b381f5f3d8daf96d3419e66ce813619f1615b16a6eafbab1952a290265546d6c1b7c2a8f09abba04511a35fa340cef1e706e0fd02c55cbb222b1bff9cbd720508af27365b5140ba76321f08bfe1383e77356a25677f2d7c101cbd57ef7f9abf85b4719aec1f98af2f8bc73e5bb16b10c11c32926ff412cde6b9686dcdab65a2b213995d456ba3db38df75766f3212791a406c64a13f4f08115c5de890aa1b228fcfc35d7c67bc9d0bb1c2e060d7e805f0b962fc885777726ae798f2464b16f0aa8befef3b08b4f7726ab0a676851be8e667b4919ea67d749f1f1a0a0d5fb9e8961ef70b2e4a5a30e2ff392cad4afcfa3e4128e79a8701bc5870f7f6449d5e74227fa070670d356f9d6b3acdd4f9cd69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2f415a8188a9765e0f4058df1a244da2b68823aa062c304a88ad299867de5686f6634c67c6941baec27fcf9e3b0398a86c4b3c14ad4ffcccc6145a677de805b449dd4ae7169e1b947403f2e43735b6bb33b0154da13da0ed942a03c531bec3e0de60933c54221c3eb942e12319d698de8ce3dc958b93f47a3f125b7b2cedbed95a34494625389f62b756e5bc262b22dc7d23d1864906bdb8a9ed3df762a755c4363a6f2a1e457d91f4763d848ecb0b3d0234a9cc19623683e7cdb1cb74c867dcd869b50b41f849b1b3dea693aa085508bf6a3eb3bdf20530f15186ee9b563a818e0be9007aea1d4fa981ef448c5fed1859b0529caab14b617dab8af9f5fbe974baea8b75d1e565608cbbcde770bfd4028ab89f06c43082380260fd4b7643f85f5e886b0495782c09c851092e74fab3e49e38273529dc3bce01cf0402666c407cdd9138c1a6cc724443052d230669eca28ab2988921ac9a0e6c0e852faac337f8cd2233fc20b3729d4c22b31c782bb1eb9a70cef8f06ff41adfee29f41c9e04d3220c43c5db0c03dead3bd3ab9d85d4876f6ad84586fc183c87b9d7cb239f15769ca980ea9aa17c6f8143b30cb39a9c55cbe52e5058f8e4370b4747f98aec05acdb6e409978c0db3a04588af09b4ea22ea1a5a3b694defd24e34463fe19d6b4488a54ef7db9790a5f4bd20005e99646792827c7acb28a0ebd78c7b4a48087dcd221df29ccf5eab5569f44a3e533b21ffe883e720f201f4c1a11dff7a87cef6eb869478f738613cb013c5d83ca1c4cf22cbfd0abc99387884b4bbe3d8c0e15a2b209e3ed3883ff324b2135e2a07a96b4df73a743d0feb2329480cc2dcf6cda59927ecd1e4b3b851b931e9f7c6e5ab20a1c7e58d19fca12a96dfd7bf85734e19c69e54aec4d44f84e645610a89e3d9306a9e1392961e323204917d9161cd91b393665df9bfc2b035b61ff47569f322b7a262f9f75304aaa3bb086cd50b93eb84acd2925f97a01fd8a5e1b6c97013d1105a8519bbafa3d1de9252344f81ecde60c231475f56eedb81a1faa08bf56470a55c2a072b022fb5f3d7f61ee9002abf2b38d7af4fb3ce29286bcce601da020b1295631cfba24d39ebb8ca1f84f98bfd7969055070e2168dcbf51550932349cb7459c994792af4f361616a8887ecd0ef39791d33e14f04ef6fb272a2b862851b790d9e2ae5a977c48b9337ea9ab4bc25b87d266acc95544a9cec8d6aa5cd0eda8b602faf5886748cf61c3ae87b7071a37e4629ff14e1f806108f5923d813c7774ec3f26edd2e59d448fdb7c4058aaa6c67c6816f4a4cf844f4b7922d745f0f2be8994d476f5a1c2e07d9dff976de6c7849a3ad102a79393fae81fc2014aeef04783e55d75c0061e561e4697c3fe91937df91328b826b68b4ae0e376ad151cd3817d28321829027451dceab851dd208526dd0559ed26ed228d612345125e65a6478d46854bf2e66774b5a8efdb435124bb7a1e0c1f7b7f2ad4f68dc7296ec8b00a51e58f662abb53919d2454f0544422b8b17cd6a32c0547349501378915a70570431d023ede7f330bf3f2feae53b7c17ce001a199a05d39ffa16e187f7a69a53b882825f368048ea010a8244b53c778303d0668ef404f276120906bc05dadc77066e1e597619289a01582089ce33049744a1390b2fb43a8d52df41e078d9eb092674be95f7f6c4dd290a5a43f21686c29aaf83492fd434265e83910e0cb7888965e4555c5a711ccded72b5f1ecbfdf5578165a21f89bddbbb9c54c6bc40ba3056749b3e04d3fbc326738bc035cb941c25119feeb75ffb9de1f3b3f5b3d6c383ec8e1c6edfccb752bbdad38716e80df9351ecece8a74c5bc482c8ceb6dc40cceb504151321c171a05d8c4f0ba447741153c9e35a6f87168fd3b129ade905e2827a90d5ba7fd38a7a2b73ee082c330d0326af97049779e3a52818f757375b485cac4bfcbb642f9d1dc06f6906211250e78d4a31068c0616c12eb6e6959c2054fed49d5ae0c15f78e50ee7e9cdcedf7c9a06df287e99df40bedd966493ec9e49deb5863de9d84bbbc8e22b89f136e85440e7c89974c3ceda7014e349651831b5565b2d085d12f40e9e2ae63046cd59dba65f55d4816f6525f9d00c78717b2e0b0e1f924819f675dc7d389c3d594d24d11060de787e9448bfc2d7a28e94ab3b05db4afceefea6850ef06af047ec235ac95c88bd14a72c9e494f3a05ff001006562b06cd1fa54e30d2cb83d5ddacfa63114af1a5c89f0e0aeb67a7172d67ad023421337db573e1a4c244e7c02b78a8ea2c0835561b9dd650e6907376eb458cfaad782408e40dfb2773e0fd2fa06fa2dfb5be6fe9a425c8c9512e780bc21eb07fdf6ac58fc971c1ef972e89d370f0ef3f0ec036e54fe3f94d82ae49c983fc66dc295d0889ab4c103fb854df42d444d06ae5c21d0e74a19ca6609d20392ec85c6ca4152707d2253b2058a9b8e1a7b8f8475854fe3086a611fad7d043084d7cf405bca4d83e7bca42a0ce2bdf6cf93b1c3aadf742e154c9d2b5a1cf9d4efcd208e4d9f6593cf142d21ba2b1e4f2e93ef34ecd8011ab91d5055e56059d5238f4c0544eb391e69a60be5b4268e02c23eac8aaa660406b9b4c2e51b6bb1774d0555e52f9131699211a70987b4447faef4cb374e6cd692bb7d559a8092046b7fe7360bdd2a63bdc3ec7175cb2e0077ffcd0dcfda1162e7005cccd91dc8845afaf744409de9cc3972708c13c82520f64087e0702552252a851a65d4ce9df8b1eef0cb72980992ea3c04b20d6bf8870332dfe72b05b9d9efe8c9fb110a9e3303675848e53918cf185c437ec881ae5b4ebd52d50bd38b63f1ecfff4d323f46dfb806bbd3384616df20a07481cff89d477ee2926fed4e4c31359c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h18d52c646cc9aba66d457a5325e0e1a95297df158944fdadb43ea266d1338ca4cd1afd8a0e23125c9d5bfe7ac3da54433f78e030d602786f7285d8ca2b019b102d33eec433059c5ed4d4fe59d50a5fadee8f9e3bf87da6a35ac9508c892c0c4323630840e49328e15fffbb9ac70c65a27603a3e6968853c04fee2d27485d51b38b8b5913ba16e1a8317d9ad5cb502170b17ef5f8f0d7497883430a4b112d6bf95040fe70d5b61558476474fe5169e7657ef75e5083f4db5a26b583ec7ec2d54f1756ccb969274e4846a32da7e7af8e50897ae306aec1f7e8b83312dc7891fd220e59baa3d1ba0cc6c4db8503a87dd75eb02ad6ce4f4ad75c9c41402a5d1617d47cedb5d4e300b12dc19ad9bbfba6a7921c66683f66e9214ede1efc2a2e3d6d78b878249d10a420811485c9207aee4cdcaf9cc43113fd4b3c68392e383823b6ac4045f5e198e4e5be3e9a6415eb3e6554b716e706c7bcde7bcd2f792a66a0eb87740654a447cddd265a6a21fcdb9b8c0982f95ed163ef042267a283b1f2e1c298eb7f656b4f75c49ea70d09b531ddef151ad372880a805519df4da897f1dba647721f904b7486c7f29e31a7321324994f434593a48c79603205930b085a5201e6e2e22f6a726cc73224a9003c9eb620123adb0d5b148e1c8eb9c60d923012393323e12f4ef2dc6bfe4e5233188b56a710fbb652923e599a08ffc616ce92fe2f92dba0511eb2354f6d931eebd34e944780b7cf086c15545ff01ab3a22d13b1325840e8670d31aa87f8ab0802f8c9d4bbf3a9dcd3eca459141282aae517156f3ffff2ccb1138d65c9f45bd44bbd43c7a215144788f5a1e761652534b61dcc8e5f02992fae1fd648975a0bc776753b32bd2405716ad1fea06314bf766176ece673ede42e772814871bfd819ec25515dccb614637663d72e509fa44943b4eb9437e97c94ebe8584066b16aee4133888633afe087584b5c38c839c9407fa08a4fb6bac5d06f66a22e325862f1ab3491fbac3ba216acc8862a9ecf003190c0e3977b55a9ed5a9ba1a5f2fc559703b5732b92272be193456c25af27c1ec18201b007e9707d7c47f2d239872e293568fabdbccd2491185170ace7ab97fa0045d164e4a9e08e813f0c757408623eb91e3114deb6ecc75248897b5b677cb5013d2b909029d592429c16daf8aca85e7a6222fb1042860d7d2efb232b9effd465be3d20c3a4690a1db785d9ab9864e4cba2545345f9986a3868384f693697a3a6bb2555749f36e5a86b0231c2b58707caa982457104d0d4eaf3e53fbd900546670e04037f225530f959b5a534e342a72d0ca3276c5609587d739519e414e8457ec7aaeeaa1435c1c993da7a9aa016450e61151fd73277cb0f95acd048f62abf54082cca9f0d6cc568e4ef8b4e4cedf73141c3a3ce510d99831aeda02bd337f70148ea65227400f4c35c0dc13b61ccda4c8be20e8617212ef6ac82543624270f1ab4389868c6c236e5e4004d16fa027465ed7ec58e75b4b77a05b9923ebd5467e73cffae9552a5791bc7b9a52c3107d9de3c750a4b483a0f6beb3393eb17ba6b8dd675748b133e363cd13891692c94a03d9240aac562f1682e2c528e6b8363994c3b826a5a0575a369ab4b77e60521aa12af5169449df27a83187514f3acf111fda51dbf8c7ca8e25abc146e4c2270e1c3b5364514a72843917f615ddb1f8e94b9cef8fe1a3af3e6e0547b2ee77e106534483d559b5da34834343b8067ac63a846fbcfc820e3d7f2a81f03023da405e29df5fd149b06f05602a9ee26f43e2220036c95ce3083d8e40098c1a9d457d36f9eb3eab442411319b53278bad0e654f7f75b1bda14ac6809596ffc348fae7913c7e5905b43582c9b95a3dd5bbd16e7de323d7ba0591617ac10a3d538b5ebac8f91f16ea172d85dfda60c779c2bc22d5ca59da008819fd4da7c2f43c5cfaabf8d75b7e6acad43c0a79cd54b0ed3fa4808a32a5878c170e4116572d3c570553dae12ba32093c3931d826818d4753c3e9def31da9780b4a63757f30499c6d1cf7747c7382dc3400833f80cedd276a13accad5f66b7e72bad525bbe08edb0055f6d202935bfe4ed3e0a6d27976fc5fdf94f8ab580e0544c3650f9e581953142f4fd194e677313931893c81587026c108412166c9aded286a8fffc9d134820f32193c3cf33b1dd5e0a3b6851b14a0fbdad314c86d0b10e8cee8785d1a34c90d4b50e7e70fef51117ed5905ac6e7fc56ef4956bd6bc880950536f5f8073299fdc08309a3197a509c4d2633bb70d557fa1d4bb8082ef2bb87bcdda21c9a03c1b25856364800a9d9697857b5b63998a9c2110c356c256e72ede7a4e4d0a7a908a249c4c6f5342d67b8fcb06aeed82b9d0ad14ffe13dcd634524f8206a9727d3b5d61ff30a91eb4ca6f99e35579d279015a8dd463d552f32196f9bb860c90a74be2a567ccdb4fe665d1cd377f00fe547ef4cdaad42f66a5a7e86d00e29ee021f825cbe4133172eb6014b9e3b851109b45d00528ac14a203cdd1ab69ec903cfccf220e986be183f6424f257588b430c130e3f887758a0189f4b79df72f78fcd18b6873c4f566252899ae2ae33dd7121ca78d8168c8d538798dc235b18352dca7df5a65c810dbeeacc57aba5354a7b3b9b5651395afc95466dc0a2b7d57fc4a3994b33438ffda47e896f3728755409ab37aab6e1f1ae6f76ee6b4a1b0ccf2a180884bebd7a2fd056f2663f3a08f55634e19e52a7dbf28c0a5b58357af0b735f709463b3c30a263b45989173a92064baf66098c237d8f0bfa49d5aa35b2df00b802c3b8ad104e290085cc5770fe02e5577d2c851bd39dca10283ed6ec53cf15462728a51ee7a8e9698e49d05308adda7ab3464595eb75b9787e66a186a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h12d044fddd65208c3bd0fd580ba2e268e4b920066a59bb29b0027ad12f4f86c49705a26ad621d0957f5b27ddf98d0e918ffd6ad916b8fcb369a2f6fcf54661c5b4b16a2ebd029fc829e4f5ab19961d3ffb8cd9c992865a651487d866ff88892fb3e56460f6c0be25c318ebf8b62c1c7fa261ca6ad408317bb2b7152bc1932ea6dad7c09e3cc8beea30a1f5c57a63550b089cc5b25bb92be0905b81b4d97f82631663f547cfe6ebf5d1774c3524a95f8d79a5c1cea094ab15d8e5a38404a377307381f3fd711d231f6efc7c504dada15a372417429b0fea496dd2874d499854ee8450401d4498453cd5f852ccf22e86489798b3264f2af535b66c6b279c7993980f7a84f857bbe798ca7621df0d453a5b3285fb0dd5dfb111441f3edba28801873408b16310f61ff04724c0287909593a399117df2c3a9b43f4f3a4cc4fc9564e0893a4dbbc98de4998c57417d4c1bd7a74d4ff7e5fd5ee156a18b363b12e54f0626de8d4b429de6f38be5dc083b10932e81042d42de2a6d0810713d74ebd5b09dfa6cff40d6e5d8124911878df5ce3d1e860461bb6b9df792b6089ef21e00b5d9e5761e70e3fd60fd52727b2616a4b2fdcabce3d207c4fe7f6da06057a7fc8d74c52eb6bb60328d141be0933f9e18819126d11db0ec7d7e4efc4b09a18af7a5e14dc44fc89ded281bc522d55fcc9a01c070d151979a71e9eca0794d81aba5c858b650268fa0c5e6e73f9e05f7a2ad8834f8e2f19907f53e0e546d8ad40c3e778e1b58f4f5e057571e2ac7b06d88af76cbea2e636c61340b3a8e2f85519fabaacee2c1726fc4b1ca622354924c11b6c98acf2c62bf99d58620eb69b855bf0a2ed2e7218f1aceee0adfbc8024d2ba208a7d9d4cee5262c60dafe48788c2c3446192f33d98ddfcd2b679b30488b343326a2c50ebf1b0c75340bc366c5b9417b84c48521e2b00f33f41ae6776c4784244e9026929821e25d4a59df88263ccb9a91fa7d5a197eb4ad26aa763e65a1fa4d64a591f8c7af1e99809c4b5c7b2c2ad8e77ac3ca2256dc5e93d6b3090213c32563e5341d690a3d75e77603fe984c23431179dc8d93ad159032a4303a0ea423e7d1c8359be07341da0a6c7cf095891e6b53cc2bb10eb1b593c4c2762a54a9207e742d9137be9c19af48b762b7358c8384c8d44188670b54ec52804c3590e56f79dd3460bce55ea60a81a04afb4bc2d6dc954935b8e92395c5824e2d1b0e027fb38f92766a424262ca0348da8ba506c70d025b79028c8e532ce53720692db5fd264fb980d192d21d233399624e85fdca812750607fdcf6e374eab1748bf7178ebf905f86606c2a029788c40b700352bbdf046682ebe950b3599b90d9bc5d88cb5791e738fb922f9e013d7722f6ed24b378922610ca62ff9b7f8bed6e435460ff7c1728c77a51e777acd575b70f34aaa1979ceb1a8f97d2db573d7f347f65870441940c256f852d3f3acbb309643d086916e454d29a233e23ac3d46c531914abc560c7b3041bd921ad388b6cc8c43516298ff166241cf12dc629e97b7a557a19f044ab21b0b48edad4e4fd0e61bd08a56a15d4ebb61ebcb568364c3179fe3e8bb3e50dbaba930b5d71ae92c0f9e0ee62920c88b2303e26531fa9ec253e2b80015e9aee8f1253f2575ff783561c42e21188549c95a0aa858af7d0edcfbf9a2683f5b9339369bb71e5f01d71a5e9f01aac6f1ac16182b40aa9e33b4770aa084b1bc0b02c35989af0b200aa3be275daadb651bd7ce4391ceb1ddd370f66665044a2373ec72c566380c8a91545ef510cb99291d8e87aefbdbf10045db51e8ede82a018a416c3dd51acfd73ee25f3198a5e7b1b18d285613421601815a161c5dedea73cca81ff44d6d9d0b2760de6ec6b19bab9fcd3a81b88316adb3f912ff7e0f11da3d40fc7ae8acf9c2581c8376eb179c6a258b5bc2da3e445ea446c7705c226f77d894cfe95ab71aefef4042ac2139fb390a6587f8b4a61e0ad7b2d2ff1d90c0fbb1844daab52f0ba15ad678c74345127158e0f9851d09fb65d32e26047915d6442d18b0553d8e8a6f66296b92e2ae1da36150c7848005ef7b40b5c91039bac730eb23ef8ffa17e51c26229bc94dae79bd7a1419ae65799f8980edd7dfcdffc1c321c4d7ef06c47c7684cddebb423569e082e1146913a62a469ed52fdf7d32abf513253651099719988945b076f66c4421a4ab5d2384ba8c3f1da271da90f3c1f00fb03d24fcb06dd80c023d9dddf222f7cce29343524881974eb775bd0511276d76e7ed42db00fe123d4754477ddf3c0fbfe6e8eff2592089c3abe7bcd33ce2fe1bcbbe9635f037e573afbf6e2d9ba70ef8b5d59e9fa146d8e807da9b4bf7eca892c10e8aab399cc35385946807680a3300e0c0f990bb702757ffeb7b07e28b46c6d48873d6ecea5f2dc00c005428c09dd8cf8e2724dcc9672b2e64f67518150eef54e7c0c77e83a0f8af2723bbeae92c633cb3d2eae43ec13564801b79f23f5ce6a0d572e2a910fcfccf4d12893c63acd13a2c5f0fcee8c2836a62bc07eaceec09c27fcdc460daa522e942cc57395253253f1db192a377b323b2f04d452077d3d847c85ee91a11cfe132aa76b344fb49060fca72238bfbc724266933fc786749e5bcf1ad589bc1c4091a9ea39d06efd850cb22ae8213bf762c13c79e1768b30221dc4c4dd93c68ea922e0d111300e5113d6c7f481736485a38b30189369a076467580be9a099f366096fa4fae51208f0a12a5ce1d256c2b3aec8fe855dcc826939c2fad9abe11295858db174613550e8be3a4d116f852233e259c01458328c541d630d9c4c67f8b863a07ed27704492f30fe50d17ee0cf06e38ada76057d14ba336e2f6df30ff9357c7ed8fb53f0adb53b207;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h136c8763ba112a5fe89c96a0637d151da1a1ff7602ba7510fb0af70c8db43930ffd6bbfd4ac91ee5e669af11c1749c4c0bd5e9ae37f16263e70ab2e782a5dc64d98d0a23675fa333c8ed721e5fb3c886707b0650081ad8c93e330b246436dedca1bdb3b6970100c29a52b63ccf85351539c2ad7bec38e42061f349d6824afe9dfb145feeda83493edb0b32581938b91634f5175f132ee834fd25587dee9cfd3bf99c0599ad30156972c7c0bc535c591ceac9e0c176469aca3370ebef93b46d28f1234bd0dab7e18124abd37baa0c34257c75dfc3fdee378ed9ba2eb49b1507ab5e416940b47996a17b4f5f629daecc17a05f4f2969424e6a2a21e798c744742b43bdb30d81e5cee5793028b2cab5f43ee51828b77ce0733147890f15ad9ca32900fe39b2f4b76a64a047f60ce0fdc21da8f68688d9cf2200024e8df81024635e9a7c8f15feaa0afe4452116362931401fba76b39eb1de72f23306297b9693058fef8cb7e80f88446b4dac923c5ddd50b10e5595320dda181fba20e8d4505994e0df26738cc8b222e35995d6114c936cc00988e194ad14ddb1f5f668151f3322a7106f29110a71fa9e4dd6b8395ce2f4ac0a042075394bcf8b8ca7f0294b576ffa7874ce1eb5a5278b05e9654114312594dbcd275253e4179da364b1c62fdafdaa0382dd10d3853b7fb1ebe1d9c1ebecca3d4474952bd1aa4302550ac5a4ae61d9fa4633ced9ceb456a5832180c1c1ce52226f58084acbe67cda998153af4976f641f35e9782ea875fc67b41595845a41f57fa370bd150162751ac3774a63dfddbb0397803709e000a352c987d7a17ca4c2060645fae3b49584cbec2189e34bb59cbe10ccda8555202ac8f7a977b32352e59f8357ae27b1ba59f6c06bc20d06d8eca40c73b8ebdcbae34102f0ea6860b01e71b205b646de5bd778dac2bc914cc27cbb1a1b696ed784e910588d057a73090487ed7cd08ab95ce06cf055707ef59963264e159a018a8f8be38f9dfd02c8185122092bd02d6071738b7cf42a5b5d09abb23341edbd7d313b244f35a5ae73872d6aa50d621039081622ae5c0fa80e30db0441cb08678dd7b6d9be08393113f247c52b7fe643a2a9e681c05a3c3b5699312d15782e3c3fbdd3786158e1171d93c55ac2349ea4866126fbe3e325f5db30f1af5a91da1936748838ba16d3447692918c34faab40082e444ec5baa4230458e80bf4d5a1873787c8b0f95d0a43f0fae3a44789eb0e9e7f6d5b92839df8bb7cdf4a352e6c6f4fd47fa4770af84be3f933f37df77917d355c53e0f92e85523fe46bbd41583f370bac93ed5a9025786e514b77730c098cd437fa1cd5361bb6e6601e272786f17f6524c47ab2a18df3b9f1e3688e72951f6b6cbd487d0ead946ac15688821148fc8c9c3bb5a34262c19510213dbb988c42117317f23a58ab9e3a7a0ce2612f0b53a0b3e9651777a247222587a7547bc10e14f6749c4062dcc0e97d127d624b5658a3d45ee6994343a4c0ed3d648933505fb132c9d2cf2500655a9203c0c7ce4c989aceb8a140738aefbdf3ba746d79da2f121f20d822b3cfb95fac065e4e13bc94facf312c6875e136f2b76c87985a89bef1f516cf7234d9baae849ca7e5ad687bd4b1e6ca988ee228372fc64a107c220ae8379eafda74a37478de9a0881850210e8e174f60c543c6a9dd6de18f830e9a2d91d8b063885b27e60427a71d09e4c23982aa7cb15f50e097302a9e21de08be56a750eef02bc29bd631d244107338fbf0788fa864370c4eb699836ea8127ac08fbd898b8ab6ac7db4bc3d1a88eeaff3fbfc981032402c0ba2d87d5dfa87a1d2584c2a56b4cd3d80559f76f38602822f9e221ab3bf9824f58b41619d6e075e91c8a0d6457029b3dccf8c52ab3a0a5e51208b0045eb5d6e424d28a0a7551e951f015b4a64a2b928ba5361729b4da2192737b1d746aa7fd088c2a88cd066b584ad60db10dfb48a75fa02983eb4362cb13bbe44eff55d1dc6b766e58d88a548ffc022deaed7f825c98be871c70084be1cc831868fccef379e65967f6f3b6577b1dae8d5162de61ce76a61e52f501f410e61746e9d930e65395f600f1e2001c48ac5d30d2c9dd8d81e4688e17c8dc041f7ba9c911890c69e8d2d15f08b018beadbc07615812ff18c6c058ce8fc9e2c08aa0ac28eb2afafd931b2e5f1c69a4b4f500f822f476190011e79211178a70da34cb70d8a306df316a0b1a5de323e6ec4998eef01bdbb46aafc47b354b421e0bee4884bab379c8606d56c4acea717a6b39ab8f5d9fb629232f2f393dcb0aec2f52722d942898e1439af486ba08fafa5c1a0245f057dae36ed1d3c363ee85a6af740757e6c0cc91e85f3462778a5b822d36f4b0ec9bbde5bb932d12c1d0131d3b86ebea0eb3ac9934119a895c18cfccbee8ae6f62a0e8ca4d3d8dbfa9943e3a6aa0565c5c8da49076be73100f91835dfa5f4bb8b284dcc0f6d5e57384e8722f244608fbb04589542e68031c22b295b80e36798ddae1e80264f5869669106f80792048be2f6ff0c3c3c2655d796024ab0f95e6598be8b1d6751f43f8400e824e988f16740f9195b48afb59cd2ed0ad474787c801b9d50dc91bc421228606ac8d45442e1f6968a8faa87b43ed3e5e8e2ff726d2b2a2c985483e567355de55981627fc888eb9db65e8d7e8252d321147c382b599f305cd8a783951131e3fda997bb4e35e6ebf94fb4549fa214f44f5cf1f27e1ffe1591608bb95fbcfa36a0131ceecd05c6851aff2d82844eeaa1be84e2217063ec12fb45ef4d39a3e01fc23837430b0cae907966aecd75fbe83a87b6716d34df088bd49cf4d108f5a96df4b1e6de03c15a2e8af97d0a833e41c546298a835eab2224de3481b938aad0cb4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf56bb668a93c9f83f788fc372f47012f1864ae510b12d4bfecf364ec8605ce475df1fda5e447344945602b7c4db515cec456372a0c9b6106bd383af0c54ed250afafce5d422942e04c275546ef98cacaed818893c8cba533ab0a049aed3dfc9f8588ca0702bf1521e41f657bf944c1b8f60a8655df19090547792b9811329eb6c35f3c2f520ae194bc24f3925a48dd2e1c337ca8be79f5a787dff5abd24d9ecacb78b1c072f7342793984523c4fc1cfcf681c1f78d4d9d585e4141e052585b4072b4055e226213429990a4cf56db25ba1b5d5c0cc90e3cc99baf6c074f370c41b9a608f217882669d6d26de46f447fea850bedc5d59a50e8ae9ec720a6c3bb83828319bd5e32d6b11e94ac55bf5e136a4db2a4b2a8a028b30ae45769660f068a382f4993794ea19dba2fab6930394d74867c694a95bd047fb37bf5a792d77f0dea379e992292bd7a6be5e3b9acae4e0b6d497442731cd15e75543f72d6c0a39d545d93af92acdb7a81161f06b7263a532d668444c68008a0df4c93647eaaea85115acecf5769bb7d72b7715f9963f0c2e321412ba784ef82c57bb3b4e49312271b475bcd1f4a4da1f0175fb80e394a7fef3d873fa2cc8f29da88f731c11285d23e9bc75a03cf0a9790d223ac58cd66f890981d7b63c4fd77fc7bb16047f72882b863e65c657a9b47f049c8b01bce369491491aea2b99e125d2469e77a4cfb48a94fa837411bfb9c7c4b712df402ba8a9e7a98a04903bf7769f11bd8e5c99e2ad3b90dd13d8449c8a5b527f648bc846970715dfe85bf69db931b93f8df8bf83b96db8abf231554cba1d4bbdacb57c24643cf47552914a532c8e793e08bee485fa0ef29e5c5a90f254c4e32943bb98d0345e7b2625b339a2e8eddaad6f9d317490c001b4ece86e4c76d2cfc62b402f8b40d02a7a33a6cfffeea47b07774bde5e016105a82f2b38ddbbd47bb512a55cb0e62df0f9f17e571b04fac9ce146b226fb407ac4a47276e19be839b771c5838233eb49da39fb792e7a1207d84fd8011604bef6983af593db91ee09700646db4d4700b172020673c25fefbc5ec20774a696a313809c9b451946d0c0433b170a4ad8de985a6f9f16b2049cdad62952ba889ea5f4fe9ab8c0d4c30885245b54d9d75b2dbbc99fe21e99c52c6e23b98171c2dfee2175080eec566d67c1d0fd348c84e76dffa4cfd18947f1c4fac244b8122b4cab0bb6465a34e2744aa21528a78392d9f83a807c11a57569dbb69ac1346b665473b8f426bf073f6f84a30b977f7050722309db1cb1dd334213c9ecd476a2e0a6b142b7835ba59554b78d20d2062cb5daa2608a6282811670f061d33181b92a17f45c1ba3cef6aa1f3af426f160d1994ab4c4aedb6ccc842578a2eb3366c41486d30b7ec5d41b320f078df1208412b53500d0cfbed43ebe37101beb939f99a0137935eb8cd10aa0df201e32451ac7464bde4078ebc3c988a54668e547e2b7e7512132dfe1d0ffa28898718b280166cd18546bddc93ea2f187f048edd6073142f96a86b26ce5abf448e03bdaee06525bb78bba74f970f8ece659226cdc5f7f7f2363e602487430c11ea62d40e5c3a251a9c55362bfcb08d4ee0a2247f9db4b3c08f91e24d1d3f722035dafe6afa39c642cba25129a39d3d47983a25c5f3c567fc3ca79d04d00fa72048924d8d27d937c45ee101bcc8a1ca3d4f5abae17b0d54c3378cc116568eae4d702471f62b12b980505d30d0ff78379c48bfd929f85778de911dfb29b8e35a737f6dc0f9c8c55b379315d9c6e5fdd6e06fe97c3b5cf4bbf970ff6934f8e18668ae3b7f0e5d3c1fd0b9cbba442ff6130ac2d0848b0b5b8cf245036ed759df99b900b0462bed9167ce18d0426982f75a7989e2098700b24b899a5c82844625df7a1d149f1aa661b1413ad85972f370c227d6089c1c0297a7e54c61334bffce4a65a9b75d6369f3cc2bd03c32592070c8468d6e714711ae88ca200d89e2d07e07fc60f7a0a7a3687659ca3cf20990b441e2abe3e8e61be0e3ae420d79f3bbc17f606927e4efcaa74bc9f7e37e28c9150f83c7a845d001622e474b2c0369e0821f93bab1030c8cec6eb5b37db60a0fe321782fca67b131ab594b505db58bcf03c858887c86e2873ccedc7061478753004605556894bb0c2b771ed11fbce94984e2909216cfb9c6e7627b9e9c52cce4f71a24eef91658c10adb97f4e1823c8e92e87605e430fbd7031147fe8241dece6e454de12b72b30b439baf8a23326c830fe0ec85f254127cf7b18eb57978b37cefec52156ca9d2ef594a3e6ad2559e2d0b20c4a5a37307561c964eb7cbbe773e926b59e392df4769d3f2345bff7c1678b8eeff1e7bd05097c7d6a2e91f53578b38f859b7c631acf1ee364fbc12a4cc77bb7416df91c0787dc0136d3da59db0dfa20065d0901bac703155d5ea4f16bda88cd77d31594d17acf74db4bc5eb9cdd8ad9fc52ee31659c8d9f3565dfe4fe6c7c4068049e4c84ce570361f6ac966d83889182f521c3b36c2dfc9540a6a9f43d81cbf26d66052173520818a740ff1c465fedf2b1c6170dcf0d58c2c29bd561b5c960a34b9ac24ace752a6eccfd2cf1209f10ec6d526737d31d2e7680d3382ef674ada97e0cc7f9d35fbbc95f484f3182fb0ade124d06c6a732c987ef2510b9e83498ac84ae3ea2c901250692cf690c4f1f83a350e077a749e2e7e711a2d88599a4002cf034b309245f51d1556594fcb1d2cf1f55659219f93035443a861a93e34a49776de1011ee17ed3e75a6bc7f1fd0b9bbdf5074db311eb12678e174dda85e51f38163fe52e0bcc52584be90bde5baa1bc337e1004067f891cde00835f09964d4e0a6219510b894c4b79e839ce489456e83f5f72025b4fdeb44293;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1f1fae2b816b730926d00c6a2e6fdee192e10d3eef4dcbbf0f1f607dd14dc026a57c3f29d821ecf53056598d0a83cf270aad1d20e564b460dd25bba444320662cd118f035776326618f3b418d74c8c6f6f239ac0709e7fd8ffa6e3c35757a520d6931f2663a8f330672915e739da0e1ad465aabeaf9a568e2d4d5fdf47eee2335240d40de9de1b5cada2513d6ea48dfc3aeee41d70c27cd1190289a558b3afe4b008b7a3ebe6de544f4c913666f0f71f0572ea77a06c2a95e6babdcd50f80f723bc6c7929464eae9e0df96642125299611afb391cc8e033dea5007954008a5e9bcee7a0ca74ea6b178794d49547ef44c20f03c271de92597eb5eb7bc20edf8b65b7095f31abcfe7afc8112128e67fc4532529c9ac86bca9d33cc01c4df661f98cff55c518e27442de19f19dc26bd3a8ddf70ba21eb01ab8319b3f5c1f136fc62bec717616b48f70b10c704d52d93fcf99fb437eff0afc03094404487abe4a702b28e8543283ca2f1405969587ee1e763ddf19896e29208215ff535a4f5589fff09c260d8c5db54182cc4218535b863b4d1b8ef46e5293f0e08b9ab085d9f1e13d6b8c118d8920f81f1af4544ca0ca263672663bc1aee80a262f2c777f034f148a2804e2e50cfb8706792232d8773680c72b159594ea3e0898d8d9c696ccf033980d5e3ae782e7e586e4264d7fca4d73ff3e19d6ee041e042a15672ede0b33fdfaf2533157b2a7ea61f6a3ad8d83f522c783858d302242f28c891b029358fb9a449fb923b3a2e4ec887a85f8367d34e758b6423d1748fccdeef07961b9dae8059fe433d21a897d29d8c445f64ac31de88a660ca0dab4364c18746103268a79e49c134161f60ebd148d70e96a692f0c5f622478bcf9aff6484fbfd30091b6f75f627ffa11ee3f7ded31938a0e1ce0ebd52ff3e02b5f2c0329a72016898bd9041c0258addbf76c153f28dd883935e5e7b31bab7d3bb212a9d8a56fcee0592834b04d9688933f0c52ea1c83a913bfb39b212e3d01ca308d1d1b90a93f319b18799464a0712ead532f4612ce7a75d13d504c4a1fa067c9780a55d63f307368bf24cbb5913a570254d170b123a837e2fc245ce8dc7f60ae6b275d066bf150a9d06c1e34b67a64ae381fa33825d92c8bfe7e1c2b7e8d5061ec76559022cd076269aaab121218d98ca4b64d8e484411aee4a374e73faf8d42dd78b4d79cf2c8d2d5e31534839e01ea229382198c14793cc33dce92a3b238583b747a49572192b2ce344593a9439eae31488492172c09840ad3c785d94724b06d75386871837185d90e093a9a158bf55525f76b7bd50aca6d0c79bce0219608d9dc8aa6632874b5068c3930e25f54e08a3f6d6e13ac89560db8705082e697cb9c2afef456b630be7dc00475bd54c41af6aef8ca29c9062ec1dd82df4b4d699a2152f481555898d572a332775d7dea15eba7beb11671a0a4f9848419a27cb1fad67a798849ab61f45c475a31166e988b5deaac37c12fb1374cd14ef05f2fb9d75e407958951b51b7695845b192c6027be04eeef49bfb0fa1adff1358bf3605786e8454fefa914536672bae21ee36021837eaa60dcf44d9ff137a0e51af29d1aef56a0f0e7c9ce2d26a7c7e988bd1c0638184bb82503931396465275fe6a431f28adc0717d1a399f5e53d79d7179d7fc7eac998badbe1fbe4af278b4b625e6d397afe5e4055d3983d466d83acd010fe72cd40a9e76ea192299eb121443a83fdc8f537cad205ba9c6fc6a128966f06a99fcbbfae7ec287b8595147b9cc1205761cd7a6eae21df8483a5079cd6ea0dfddbb55a24f4eb3d5a8a4d0c64fc638c21fb56d50f99cad90c9e67bffd2c55a253b47a4a3f741d1128d90e8fbaa12056803f5da7d904190a158a8b5508207e0d93078501851390e123da16807f6ef37a8143eabbf5ebfed70a3522fac6dda4544e5d064d067065ff8edf30d394b5bc2f2a1875e5e4cfdc92d3276608d487d15e000f2e5e3f746a3d830388d89b592169d1d24b745fa2e8d9b56aca90114db078bcd0db2b76c19752e0cd82402880acc8aa7a22427c7a0d149b80736d1678b2f20c232ac415361a7d6ae0e0a2ef34615bf0f66f48952558fcae61ad118930fe562b1772d9fd02cc43c2d4108c58b597c048d385ab0988aa4a3b1a27287b8cefe10c2d91e2018797802dde2f0238577db3dc955f8e91eb84dc4792da20d45fa17fd005334bf8fec4e1f03edf02dc3cfe35c64516cb77a28314b15a7655ee04729d59028844a449dd247f706d47d1b66712adcaac9d04a4a6e8e9a6b1628efc77dc6ed5bb434e1f7d489904fc03204658e6916eaf536e5ea76efe3c75c2aee7fab12d5e73f9746dd4740f36e60353f243b2f99b4fcc5d136432bc497a7051dec074a3c80c3f109377b804ce50f9bb6825de3b8c3f8baafc71e82574accaff9bfa6008985715d0158988f1af6756965e01f7e28c890c8a0c4479751a8f94ecef9544e6fd4c6b12385f232076c9caaa149d2b3d9e1cb7c4abe43948e2d28ee216b312cc53adefe585c9fb602088caf05134824a295c13d48bc02e9ea0e8f6268863c37311fe673974fe6d1176e48d2112b7ccbd73015e605e578fadee0ec242f1393bab4e472817d89a21256c782a4ee4cdde23bb2a33800936b60e49cbf64f24d6814803d0ccb200469f7b7cacf4e0c5aaf172ee245f8870eee0613e3cfe389c1282ba8ba59e2bbdfb205b73fb3b032ce939f40906676197974ccf2c768bcee6259850cbc934bca545f95fde1d1ae6d121954faafee99a37fa091ea533eccb0a40298d157a99eed6b8c439af13c7412fbf85da1ad7da97105c42f4d8c23c2f261b24cae38f2fd604c1fec91d49a22c3a6857cdb72d820ec317864b89860308ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbc58d4d4294ea0aef308f7003f75b3834749da7bc6dd9b2d3b283649e6d8fba9a0ea8bf0211bfdb3ef2c5909c223e01a02a2f19d5b9afaa759354f1d9720c6f02a165217da80cf12b6c1fb6f33d88b04e4a5bd71dce6d568d7b22932d9771cd8f6f8cbf22ef3e1944f211ca5bdc117a031a74b86f919620866c78c5fff5f92ce84d8959465682b8fc45041110a4886ffe0dcea9f5ca82b95acc8a3db37d61e66707e5793e5ba1e281279ae6f600b26c3a92a4ae4feb9a3226623ad08877e9a7e454c716c7e9d15a2cedbb71a700c6ec02bb3d8a4f767b631210adfee2f5e6d835db15c998c241fb52b5bb04db13dbee6067fa6f6de44f5da89fdf186dc041abca77b9fc35669a0aedd24cd32a042c8a93aad3f8d390b18f3fb16acfb6d6add463d7f43164ad67ba0ba235f30f93868fd31e726b512f4fdbb30c06b4f4c5dff31f188c5388cf4cc2189337ad38b059a14efe5f0ab5c20c71141bff15f369cb594fccc2187b4d066f9481d6824c548d49288ad78e0499f2ba120aabd15fa8a933983d87688b1f07a3ddac1ebdc899aef5a051f90d058fb14b7a44d9a20c509cbeab414962c426dabec15deb680a890dbb889e695dbf468fc0d3638be0e8937f691dcd0fe2ebc8b717ccb0969f6fcbc509a1b33a9821f337caeb631b4d2620444f3b482ab1459d63313c210ccfa2cfdcdc1bb0f0833796145b2913d86031b2d75aa7df66b9999c9f833964e23cf9ca0635403631a9a00eefa2b802031fda66e5778f0224ffae0da1aeea18771e8c7361356ff4cf312c43d517470ce752cf32489b8bb281550fe982a1a60ede75ba1a75008f3b39e7ca680890bdac9e580c9a8fb7f80749d79a33a5667a9259f438c039d55f5429c73cec8513b3aaeefb0de85a6f9378855f930b37a3a7616e9a88a5d492b4efc96e3daa1d522ce394d6fa88f11f9cec5105a9cb405a121e639196513b404f86118d264552ff54c12baa27ce29f6fef71c0ff2dacdb60caa9236169f15a72e4970739ec0447b3e341fbefa3a1ed219ac1755b5b4375ecaf69d85f103715d456a36a695c60235aecb29317bc2db8589584ac983d88603fe6a11954b66656bff3085e970e7d556719c466f99d8b49e3c855de5d34ae3ce7ea0565b8287fd3684ee30d5e2cd7b29e8ad2e2dce04d3f07e65cdab71ca554f3eeb2dd4ec0920b1c7cc7d162dc40f26704904d7f5bccb1d181a79f291d29e50962d23b787412337180296ea711d463c8f82094db2a899a27be669dc8d127d005e4ec25a037f3c91b6d7fa64091be2823ff77b02b9cb534e94055bf2eaa4dedaa47be9769b1d1c5f282b659dd23851a67d16f3569ecd7512a012048cb0a98eebdee76200c538c9864963d0304bc6c40aa9fdc893316d2dfed57aeb822a69303541cd0a768ed16f806e5fd18f47565e3560581fc1820714887c6d7533269ea1a59ad8533c6408506ee44533cd8054a2906d58561505a6e12009e2e55bf3b7267f65f66524bacaaf5deda41cbe6b5a78031fb80b8189983bb75ac2642e97372e93a88cd144f08520d99dda3edbb9da66ff5b59170797a669646f671301541c450a9447478dc39a5fb90d9cf149db603e835870704c97e05249313170c1412ceb9084e9ed1b38fdc51fe708377c6f93d3689dd1c7ab6ce9aeb139888c3fd18a3b3fd2484b2f297abdc3d45731e532f6717dd5e9f9d8bf537d8b3ce0a66dc7fff6f015690b49c901cf771365131228b17eec046ad3252a6fb085d4f16e9436db06c21a7c57fb561af5c840f04c6945efd665c3edc1fde9ff691d92d1d2c1591c60579e3411c3fcedb10f6f0df8b74ced28d79dff0942c68139b4e9df6c3d3aad7365ab9d1cd89c8062dd74c49b4676bfe54006ee46ab041618aa2cf7589310df744b882fbe2cffb2901623fe75b1ece85d7bb69b8d9d4ac9e0442fb33e747e2aadae322a3d10396e4482b1143070d56bd457ac186db0e909bccb75af5c6c9e186b75d406f1295ebbbc5e0be7a0f121205e87ee1ab6ea0f0224ae7fbe2b2f8b6f0743267ddb752101bfa9c819da72e24dd05ad26e189c14496458fce4beafce29349611a0f615484033dbf84ac3ea1258b62e89d71585f1949ca625ca006d9bd156f3cd3912bd1191a49b716bc7defd700a26235719dd3af31086da7066fefedcdbf58d7d345934c59f16a30a6cb406a91c4bfef26694273ae4dbd6e06634a66af1b96c351f17d3da02256a4f7d2c76bbc094ae763dc0734e6eb6b4d54c3e15a2f4e37416d6197915fa41258dae45441edb6e4a807f0193fe0c80d96861be1c1c7cc4c541ef42ab1e878bd71c2bf085c00bc9d6a41405957d8641f358b0c24b241e0cfdb8cb53eaf8ade38c7c695b463dd7ad13cf3e94609c9466b6bd61af329c8e5a88e3b4bba38e4469923756b18b17c23b479ba75bdbf8e108211fc53b1abdd640201c980d782bbedbdb7ebe12be38069ae8552a374a0cfb24b96bb96c620cfc9ad65a53a5dbac106e4e9263aab3d31efa7edce7c750a194becc4e61fcc3fe9e9bc9bf9680db5c4338d94aa495c4df1e8a54998e5218f7765b39895268ea84dbe6b924ba1b4908e71d8c8457f900b1b32ad2100efbed7d9ef56bc66f19f103b363cd2f51ab08d1eec4ccabfd9766ac2da4439d4550ad230bfc1f0eca3b401fdf73660b84c411be5399e34f36e788dbdfad429dc9cb80df0243ba743d7d796521d01a0b06a42e0c1d2dcd43eb8bdc58ee902f784652d70b56f57c0a636f386357ca5a28d7683613f23d4eddf9e67e3bd57bcebcb79dccae1462cbb8e887021bd058f4eac224fdcbb360a30bfd16aa58f04fc1fd1920f28bb0c2b32ca182522d4e8149701ee1b57b1f73e6a813ed39735a4a1d526e6efa5597ff2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h307421bb67709e3b42dceb81572e1a1eb81fc9a6981620798266ab92cf9326ec31282b4bba5756ffee8cbe0d0db2c2cabfec3674e9debc1a597f3673eca5d1fffba63d5409d349f88a6444a3aec4bf154cea6043aac964fddd042ff7509c6061002b95568017ad45e1673e70369685d40784b1635804d429a5fecae7d94a0d220fc63c9334f721ea0427ab66a17f8cb858346023de362cae1bdb6578fc46d90f86e4135171bcd699e8e76c9a79179b25ea491481a3d1027314d296d07c979bce22af9fd7911e2b86884ba2467b5208cd82ed2f37bdafee56b49bb8e2997cde6d2b0b16c4fbad4e6dcabadb538f8e691a74556283a44fc35e212da51045fc3cfc77bf0b788f33a742d183470508c1888e2f0b25d4db381c879a0252a6cd900ae15a8c70aacdcc141867b53043236fa16b252a58f4a96c9d0c67e7111f9246ae020b919ece898440311aba3afaaa69fd5a7429e2cf59d357feeb37557270001859f7eea7d5ff32a438ee88a986ceb50e4b92b08a9021ab883d630898e56be20622233f2337690e9d32a3e455fa2abcbb2fe425f9d048b7a05023d0e1a98392de85021d0ba957e5b3bb55ff751df6dba499b385aeb75ee40e258d7503bd4327636c05b4298f72cdb9a4ce9bdfadc68667802fda946b7ede54fc35179e14219ee5f4452abf460152a05c9f7c124b4069cf5b64326e0e0d4262176b695f8bb0e6fb1f9c3ebd7736d3b903a37a184fde035de1b4af50ccb6034bc4ed6dca8bc8da6d65c140f199181a2be22da9079b3308690b363107a31eff14e61ba5d913827eebc9d0c78ad73765a59a2e6dcf5d04281d36308b434546d7ec57b3431e821bbfbfaac659689cca2d26295de682bc016f69f16c37c86c6fb0a9a4be98deeb42f681466e5c4ddba7c385b23f6c70111d9020dcb92ec00d6f6fadde9d538d236185744fee429c10db85b0aac12632b1699dbca18f38808680020892d42770198147b6e04a2416997193541333ab62961177f30035b86c08c6f6e0f8e4a33bb130695873b22a1b6391e017101ab31c2e5f279ecd8ff13b91b9c0abdb7f5b62dbcd83f417716610f59d29e6dd54f911a9a31e3a5d3487b3e14e46121cf940c985bcdd34c727fc11f928567f1fadeb6d9efb9d56add68dc967830bd7e8a11819c28255be99e754194dbe3b03b27d3c1919ce78a014944f8cde5611491e8801fccf4a6b517b96b5b21576b2c2cdda877155472aa1f7311dcbba38a5a0a89f764d23f48bde67ce4541e756eb815eaeb717e82de7ca5615f988be0ec2d88b2d2b6b79561bc7f436e0a417158bdd070f4f26a3b8c845556b94857f3460c6ac6c0f44dfb20483f8e1e560eb2dd3516912e0ee527111dfdf4dda4c43253e6c079595bbe8a1df9869b98c5f128777a4cada553bdbfa16fe6345dabb87c10da65a834f8dce0a628bd76173cff9804ab5aa538f7627e0f9835a90c6fb57a7c5fad3d59123148e78f2005e6788cac609720d304eb298f1637ee0e047f32ddcf6662c5caf701654b3a13a246fc9f694838e957a547e33fd8b691a127097f105c189e9bbd686675bd89f657d31d3e695577276e3f384c2b1b24213581c8fecb527d8c8e372972a6bb1f08349fbabdad86d38a5b2eea2486e6d305fabb7db88b1ce1f0ef4e82a08b737dbfe90067a86df510cb535fc26234e49f9c4f50ca88c2932079e5dc49716b01810731ddb6c8d5593276bd0a96151f53ed9b8867929ee97e1d459c4a2a406e8dbbdc4ee3b0e173c29b1966f1288e1a324a2a340d2e9890b9876e65ec496f890b449cda3ecec9ef71dde5a9043acdfd771b359d6baa11cc365a103f6158421eb2364a978e72891adcac48f81d7c16f9a133f47fdf45767891118cf14b088ab6355fa65e57a0ab873cd474c8d6ffb29d47d891d738070f58014a1667eacaaac9ac2b3a0c56154e906c0fce75c5538e9e8d1fb0a0aae8f08f8b765ad37635d45aaabea22127625d0a23bd82e0cc2a99cf9d2bd5cf5e0cc495807d75887291966a73a1da1b719d948b8134c5168d23effb2225e6ae54298914b63cdc431f7c0cc51eb8e322b0bddb3b9acf4dd0d30c3949ea6eebacabeeb282e60aa94a40d1dee48b50d907cf47878cf46332c4895aa4a85082b599d61e03ecf6c9204320c193cf060a930b06acc2870cf4e458114e65bf01fc07e4ebd1427cbdd01cd14e821f153daa9c78be5d27a80cba6a56cf1765c848d4d6d6d71ccb8de34f3f15753a77e9d38e0a67acc909dbc39c2e9fed3069fa12ffedf1c404327de111c99f5ded837c34235bc4d18db47bb09e028d684d42b880dba1bc9a5b55273a22145e3fb3e50136ac0d7ef5dc21e57ae5be888b36a5921151db6fde8a4db4c2168b0480c8566f6eb9fe6ff350a7b9788b4a5edfde7cdb68ef819a55c412544a30b0f40dbe7d3f4e1ae977f2d5356a720daefa0cc83472222186412feafd8cafef3c0848c37649c11d037fd63772bc19645cb2b8107271f59b586ab5b65924ab50e8e5baa31602277b697e059ecfccb67f6ddde83ee5a17372f7f869a91f6728111da2832ecc85a2046304d6c3fb491be22a62b252e36dbef4740a75f9f40ea9b669a60aae760a488c7e4bbeb624e1b33adfe966737cab6cd7956169f7afbca30f8151eea1bf62f1cf435d2873aa70519ae8dd71dbb2f3a2631547e97b805720e57cd2d9a538efe374b6e87c66c25d32eff7b67ede730ef3710145c7e553b9a59f16533095e04fc3c06428db4a69966b560987657194e4502841b0d9baaf16432f33f0d7a08d36e9832400552feb47d748109f5f47f730709dde1393b7c6b3f0645f05f1dab6abd503dca1e4fb67d63b27ec33ef64de30c5ae63957553fdd2d954eb7feef28d3743bf938;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he866940815cf4697d9e59edb926203d8c13671057c2155bbdc171c789085f1c2bf2b833322ef7f2b1ce41bfe37b6d660708ff74c97a768a9addddb3aa5bfbeb315b58e6f765d456e83fda928fbacd6c7339e7e6659375c1025a8dfe6b216d006b4e60d967ea600575b430c1da8d56452943fcdabe8d62caea39f4982d0fc2e3c068addff194a5c6c52ff8d55263e338e1eccac54a32839ae2c52676ec2c38c99ec138130b8cbaa88f523344a3c490754f00e6ce60b167ea2e772bbe1275c33743eea05e99c53b40b373b176514d90d46b884c3365b576446a3e0de0555c8984745ef6847e05e8b9e3139b04be5710a1f127109f2f2753140f584c436eaa09c883e515a117a2944cb0a0f555b971378b14e0b4932c5557ad788efdf53ec5536bb4a757cacac7a0aa743a4f8d0a2f240b961e9fc6836585cb87d374d0bfbb230fe3865c1a3b7ff91c163cb47cc97621e1b207e78b51195dbe3ff7515b90ae6dd08fc9ade26d785b2acff6f56b25f8563deab4a91b98fbff61312bda7929a7b919878ec362c5fcb867425483227011a7c988160dda42427017a95d3ba50f10ee26b8f163a2b738df817dedd5834bf2a6c407478b16c0795d2d99fd7b31f97ddf192f18ec349791d15df31bb9076c31b4ba230c62313436f687de54381fdbdd750994e912281095978069b501de73e7ea8b1f9c692d6a7a1933325fa3f0d50181f3704f61171ad614e9b2b1ec309fa5189c6177deeb1162d0229fe2ab6d809e51dc54f95b1aff78de3ac065b8e3c94c1b0eeec28027accbb7e566489eb5a99946e67d5ec1ed971581ee76be5edaaeb9448963f79f27ffcdb6e7cf8f5fa31117873058fa7b67de902773cc38d0f845ff1ee2c7ec223738048cf841a3b2c30b3aa792711feff0e3710ebe819b3294d70f225e58bd26a22c638c6a1577f043fe18e66fe9604ec81db8fd4ebbd9db7e8d314fcc4c04386e6aa8d3692a0ae05662f4b0efcd338e3ff5e8bc8b1152ed99d967faa311fcda76cbfe51f8434bf90860e5e07fe4653d28aa78bd25c760d46e8af7f98def59aed75df23070c38c9a95d03b0f49cf703c306a6721520e2e8cd885830985b78af9e2d76964ac0d49270e1f6f16ef9e5cbfb2041ece4951c5f7b69a5bff6c9d52195bc1ae9ca01c05e4b3ff193bc4180fb631e542d359186bf230c4030a99631601d7e618272fa8d16d16c687991a5eb0feb4e74051a1316e44444fb19ad47c8196e8ff876ec5dd09d2e7427b60b5456f84627dd87f55fc1618173b5b6f06ddade56cb85b4f9e64c924da4945ed8139f0369dde9e55d4cd14e5a30e1bd0cbdf60de000668494139915b66f37961e6a65de19e4a80ee6dacdf5d531af37420e812e9eb0ce86f9cdcfac061ec4610a6f1c8e574aa0b54aa15254609492854e238984ecbef8c1c6c7789d7aea47a2aa6e5d2002662b4790b15077ad9a52f3b3cc476992955efe0c7f765fcfc58d18979b2cb0a795fb94d8410e1d8a79d45c45b32ecbd7ea31a76b717652d394f9eb82b91dfef186305272b62e342a4b4c774f71845160168680baeba9d6d2c0ffd49c0cef45b1314b312f1506215334ee81c5970faefdfdfcbd5a6b34eb3f3ee88318d442b1afea6355b356be7e59fb3fecdf9dece15086d6fdb5469d7ac0aee36d961f8b5ac90ea94c55694b86569be3c42e10d71ad326726b54533dcd7ec203ae89dbf1c4c4bffe63d71bc062b4ee71f17455209a7cd808275e41c895a116dc423c37ef5cb507d4940b76df38f3eee6edbe34b0367ef35997c0dc9525da7d85d3a68974ccc102fb1f428456ef84d7305d7e2a3f5f2fa0844c45047b88e09c0d78ab116f1ce44d7328a2cfa3b315a1e2f8e3d7988fbd388822f688b0a4f82c9c33ee3c33fec84e3e282ae56bf6ae23980b1d7f0755c2099995e2b5e0f586e6dfa75ec76b7d0daf56ce1f75f2282804e5b99d82f180a930e9c8d97db31d9ceee6683e0b10e02fb9f01dbc27aec707eee7d033c0fc88f79902aee68a452f7d7a38ba43f9c930e43535e32dd111064a9e0db93d453d71a594d4997764f13e62099662e1ded4bd1595c4fb70a5b2f78e60111e7f2a2fad29f4eb4adab97df589b8cf5d9d750609df17a353da92341b28c035f8ffef2a79d70b738d03c304904cce532bb41f4584ff795e895106625ec16fe50574c3b553d886a3e8926b0312f9edcc9e14f22ba97ccb8855b0c7153ab73824e4018d3879f82818b761f7619a4c40e6ba882e7a2b3ae2667c711000488d855c714a87a3321ff3c181a44e69512d4ea2b444601fd5080b0a7a3ab59a8b050e2010bebe01ab43cff7ee6e7306f761508a4c8da7810d584bba93661205edca02e6e1e6a3a78f053661cb9276d618a8a06617a32df680facbbd6e5b781cb138966130237823d77755cdf4db4ac7b06741e8cbf78e8a2f2cf8a91d7e22b907c3567584016c6db4fef55a05caa1a7dbf1b9686ae601f893c2ab10d35bced95514beada5bec48b860e773972262c134c7da317b5a0757bce9ebf153736591e286bf6454e52ecd5bd3290bc82cc6ecbfc6e31323cfe0f82d4de05c03c20135e2212b9973c9f0c419d342bc773d554f338bceafd5627cfedbab228afc193a889c12254087bac2e883256b0d89e74aff0e8d3de0544a6e8216ed57b36818d72bf3d938eb29f7cf0e4610eca61cdd73693c35e1fbb977c006fa8a8092ae8f13e800e9976c209057c8bc2c1c6eb1b1f51b4a119e9bd47c92d5a453df8d77e2300e5637d9278567c56c5629f7724bc5bdfca986a0268dd30a18df6f8aac6bd1bc7ef315439e2459535bfb34353a466555d8f7b5842fa91ee966476c3bd9c4ed52f84c367d88285a01bfb27101d65ded795750114ce5a071147;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4298bfc9b716a378c4bd845daa28aafba2613d948093d90a032a1fe5f6d9cee3106402219c60a44cc27e1809a5ff157ee694bc521561e6e8ff8a22ba55537c980ec59f9616ac4e429cb0ce26572d27c3076c94a9d08fdadcdfdc212e6ad3747396ee70ea217aa713dccc73e2487b7c2d6ad80444b142ee7090a05f400d70a24861464558998975c57285907323e94830eedbea31d9061791ef88b8de0386ec918f8a32ec4f67debf9f9c3dba4ea571aa2eafbfd0799062f311a0a3d3c3887868c27cd01d6f4adf8b32e68692628c6bb65434426bfbb85be4fbfc509668cb9e0a83f299a2087c77050acecca575c761b6f4f574338651eee585c40d4368fb731aa3a0303a658f2f4bade4c606e753bd72c316df29fbe45364e47410396162797fe595c6647c01f8a6aa376e838ad3d17bb94eea1bc6af7dc3161b6eb0d322532fec8c52d2e503c54163d57491ea08aa59fe7f07330ed4b9c9fdfa45ce92dd85947b51693c02c04a6ab57a926e23e395cb86b854bd000a3dad5e594b33ce2fc9089d8d05a84ad1d19ee16897ec46a7099c29d3340688fc1bdeee63280002246b6fe3b2c6a265554e8994913597bc98d1b79cb414fd5307e752812130f0a849ef035a590166870b245499d2aad22b62414496260672a5cda411de9570980c9d3194758512f2660a64c6d6ed893d0569092352e246056e8f7ec97712c67daab69a2e4a7151a749bbfb5aba5a29e0d8583d55205ecacc3db20d8619053265118b6f9fdf2800fe496b9b4ee9ffb9f2c8c557ed7587f8b47bf170b4f21210934ed58395f9028b6b03c7372c6bd9b466e618e4e49c1dea42105dbdaf23c9f7dd76bf36d09a361077686564ef17513c663665010bc277d855f62812ff9e4fc4e39d03151bc67f0691c0d45e43705c1ad1ddfb82de7fd9600a32f8d98cc8f9a06585642057b5e42e08a36fffb0bb7beb1635834fc5570dc5f4176fae5fcec9c03e0142d55fe8e6fd73faebc4cfef61ab4da737660c86fbb9b7a7da214f254c45e20d3944bcd9a0fb482bd49a5edfc9aa269bc1b9763530342fe39e60e2a544d3d0e44d98914d3a62db99ff742a2b8d76a1faa894a01bf0c72fb58069cefad437f8fad8c80c375b230865b97bb626d2a6fec7372a30b92e68f50a0a78bc5af68265f3e327f969d74284dd18be22bfb4bd2e6caa978e0048fd007c1a1fdaa4cf9adbde43e512e864a2ce5aa61b9ba9196ef08afaceb2c0b9d5af13433f72740d637bcdfbe63046eb9e074fc0c14931790b0e81a37df273d94139791f4969a790485902850ae8a812e2d12583495eb31a9f096a46c9bf89b7b28633b000e1a24dbdbaeaf51b5acc281fe44da251a32c527e3c48e4a9e71dbe255e3ed52ad00f7206bcf920be5d6754ad4ab11996a8ea226a577e8a8f93f820a6d27b6e9bafeade8a6333b06802927759d23d2de1d2af24a528063eb9ba3f8ead8c8e96076fa7feb164fa45607f811fd127cb2607656aacdbb7095e2516a09faa2c1345640f7c2cd3ffed3a69461df92648ed2b9250007c8f97119e5c3a1b26b93620205692e235318e737fb4696767347fdf6d9d104a2951ac87fd6851059b8b3b0f693c0506b08c6fc5ef60bb7bf195cd6730d3057da3d41414647a2dbd74072b0ecb3c5c7bf011130346b4d62b9f1c6459403fb2288dce7a32d7a069e3b6e53f947c105775d97ee639021f7de8a8cf8200a5f29f909d3febc591f2e2f6efa7825f97b5624919648a19e8dd866db3d3fbc24c8ba02a802c38fda13b2217b197d4b5f4b2ad5154ca914940c4fcf41686f91a4b6204d50d255d523843d1ce36ccbcbf1abca9ce524a257f6ca83890ba2582f80db9c1bc03552b87065b927327c208458fa85621d631ed516c8f7c9e8b5db1df805c15a155412d7841b009c0743897fb050aa2155ca2548beeb15533337a678ff89cb4f382b79f146605cac09672e3cfe30d30589ec084c410b90177b20326d2d19445e9aaa0b00693820ae0919917f7c6eb477f56b3f3bc02dab4b4441e93f2cb9e6213e4c67b49db62f8269bb58083a76659ee211b5b13adfb7ebed1d43d47189a37a1e259e3877537d09bcd2d6d6008f585eb1132969eed77fd3717ee8c7b0c518bcbedb12d547a0b0479ec2fa36390ae037a319d05ba2e7f3c432f2eec439c09bbff4cfa047ce44f37f9e39eaf90a0909b62a76f91e72df21ddd5855525416b2162c56377efb984c8dc2163f1bbc5cc2e6daaa6beae9a7bb49ff40468f697e4611480d24ae10858e2024808a6693c5ef0e7adfc47760ca774049cabe3111c445d616d44b32a599ebbe22e6ab3950755d6c2631e517c82f35d525c3970cf4d6598d87ca3454d077645904118e803eb3eb40dc43699bb31c92ef3de502ca91e3ff831fc69a268efa7d70c6d4ea77e3f531966d232b5c82820c0e25aa241ab29f79c9ddb4cb70e7e506dbcce3f1abff633a0ac5e7333c6b09a32fac31bf8e6cbd053c9120e101bb4001f130f6b1a1f3d567067a558cdbb7f3279b728ae7bd9bbcf1da35fd4738f7072c774ef0bcd4058dbd628579c2fa06ff339f158db2b39a37d3de7bdc179f192605314b1c7aa74537a073314d3ed7df4559b4aae2188a32a9872b31703dfce10131b3e42de901090022e835ca7ebca7957d725c323a73cdff8bcbdf4039dc1f452916be2c3307ef09e928514cc93fc1cb4f4ef3e80e5b0aeb824303acd5a48cacb58ec472796f6199ff136b2093b91ee7b4b1b1924c5842eae9a7ce00259b0a73fc971a4d19a75020ea576091028fb2f4989ced32f3d3de0f50fd486152c9b1d353371433693c031f290a446c165da918500cf6c8a569cc58b47ced8dcadd5a442fe30c87ef40bf622ae7ce8b87e54fe3dd1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf9dd69d800feaa6b682a66ff5bc924ae43a1f36ef458c1ca30285e212e080c6bfa48040b8384a845340f999802a63942bbe5bd4779f626ab263a4c4a7eb9872919ddf509edef0be4fded02e4fb5202252fafc53ffc94d68ade3d26ac165569b65725d22dd7bf384c13f203bd2cc99acb89713a9151504da938c41c8a777a13db0fcb9f37b421e318361661d6a75190fa6d66ba343847e237eb0f32bc195a35d2dfd4cc6194fb007233fa25b37356c2b834cbd8c94d6f0101193768d03428b6124854753bdf28768990092bcd9526758ef4580eb02299033f5edcf42041522400006904465390eb16737b1654ef336599b91b18a7b29d9a2efd27273a18aaee8b679a47a99e4da1ed1cbdf756ec08382a65ff3a5718b2047a5f1c79f27a5720d690f551cf76f42c56d171a66c19133e7f926b0c612b45bf150e9276fb2a664097faf8b31de7befc24bbce51d5e28f575a383ec495e9b651f5ad7b2650337a06abfd8becd0d7a4027709bc1f73cb9ef7e30e3d7e312e321fa31cbea3a4025aab361f7fab542881eadbe663b2c1b880c7151ab064020330c5a15cef1fcecd5f5883796768f3676eb00ce3d0834cfe05aed404a86ed8a4fcd9fcd67d9db0495a7d67e853faf8a44d68be5fd829429cc3218f9cafae909044b8981638c23739e6dfc1feccd67cc970f7be6ded8b80ebb776d9c1bd9b7f533eb4ac68761535abff22858833bd8c38784b90a07c6bbf2cda2d175c08ba64be89deed23b0bcb99ff3633955f6f2ffed82e6531d936ce6ec7e995f1fb4c2ffe126d28a063c1b270fb935e80848dc719ef44d9d57edece443268cd40db1987ce27cce0dc90e5e03aec094116176a1f8dc44d28e485c42a8c311760a37cda1b80ce29fb22ecd555abccd2068a53fa5ebcdf5688089b65bf12e46dfca745da8a9203986b9861af08dbde04fc8e794e04bacca570e90fa8b0ca24434b4f822bcd288f3882ea3b598a53536a136f15ad45d768c5a8ce2f35f0673be25f842f070ab7731af00c408d83e6cf1c88ece90178cc39b4f542a882e03b9e32db476e27bde53ef0643d782edac762a2b1beb5dbdbd7e962b2a19f13b3774d283cdac6967e8e6f57f54f5d1f3b2aec3b52e0ec6fe08f8daa5e9264631557a7b041fb1b024e65651f365743d19ca56ddcedb8581489d1e129a6287194b7bd073a86def83c4aa4002f326bd271abecbd81c1d298e50dd6397c3303bbc91637ad9da3375a9d7fb325104487269ef0dac65f0ae8d0ebf54d777fad3260fc19854e63383f4fe11a36d3a9043d22634d7360c549fe9d1532f4fd70ce3c484a8f9df9016ea9cae3a1606348356baa7ada9a25791a19fcb72116261ac0bf92e4cf9fe5d383ce37c50c13d91ffa65ea7478bf2d07912157d4cd8ec598ad129eb8ae556ae415d435a2082906b75c179db0e056590546603179ed6a5929c754a98bb877d1db049f8fce57699f8ad317888bcebaf03acac8aae2df5df22a85586f577acdecc8f390c73ce2f168ade5beb94b33a6a82ea4baabc4f75d7114a74ac2bfae89a50394baee2125f75681ddbb51b573ac707308462fca1f66b88eec2c6c5f6b53f61f6695ff47c41149d7255146cc83b1b2ea2ceaeed35203d5307b5031989ec7dffd9f67d0d927abea939bfee4d2d88a8d5115e5d0c37fcb2447ba92f1c3d9854654af3649322fff00c55ea7226b16eec077d597b61d01635581c78cf227484f648cd31fac84b38b3e62e55a5f5daee833591bfe417d251a440c57ed444e1fa076572c4b38c4ca0ec7951a442f1859dadbe51f4489103fc385b710b25174733fa90ec43dc75ef6f4c3e286e85b800a09a221d87a0f68202f7b50f1114708eef8d98f4381a8f66b51bade4f88d0f2d46ecde0e57af32ac091c391da1d3967bccbdd499ec91de0bb41a2ab2a096a893408688aaf8b47b7bda97a71d77b3b81f41c431a55d452861cc88ec16a3e8abdb8129f9a94938735b21b06df386323423b1ab2d179f90f47dc9d61b59d1c3fb277a9d262df2813b2c27586c4a5f7780b2d756507defa9b8475e1cebe67e62a95e1de350c069644042c2627a7adbb33cd03abab29da5fed28b2a8782c2d12a39b0d6febe2ec66ddc9cbfaca7fad783ec68f67547ec79c2929685bf6bdfd560a4f87872ae956e3fddf09d46ed7bdea702a3749126f3972ef07945839851284aa283b769e65d4a37799a0706d907cb299e611a36dc3058a53d79e1332589e10ab0db2cad6f419244f1a330edc77b57d0ed526f35d72616e9d3a5bbd0a22f0372ab85d0fa0933621714c5934af5f23ab7f0cd701d0b7d5dddc93303aaaf858b0caeb9df04176446b78c097c0e9fc182728bb5dee99d68c5fb15badd3c3af5d841528f3f191cb653dee3245b218ff2b05cc9592fd1fc96e9b2b672c5addf27715dbce9fe015bead9e1c14c24f8c1ffe95aa6236409bfe0b92bbbd55ece8579e281b32bd60740731568c4723164923f0b813beb9b31192660c1f63dd0b8c70d224710b369b762729c211c09727fffc601e21d52ea8ec41223b32d12df72844d73e486a2688542e57031bba1664df9e2acb44903b61c0f5d19e8f9057f54ed3f76a806042a499837247d7c5c6429924ccebd83ec79b4541b678552f0855c0d5a54edae25b14d7f02ac379e803bb80c17319ef624c0743d0b1ba64a5ac618b1fff22f57ba4bdbe8476fa967e2459bea34535b7801cde66b2320fcc4e5e3abe23e5d5b08753def6649d40853231daa8ebd6c0acb6794caf77803639aeb911341066c62c702d644d8686e6a79caeab55ec864cb0b809a22acecf52ff31157c76f56ea2a0699b99686fe2477dce1b875b077f2111b539aed3375993451695f9ce7057684093ab3e292a0a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h741a1bbefb04072b93e4a5e29a25031ffeda16716e38b1d7748d2854f413c9c37a2fca4c174a8ead441780531d2af197e5e6d1c3cecaae78a89b5150b4517cd24164c859c93e76bad03e710375e0b87a4a148682d2cd0e2788454685b7dea3bce99d9f5bb8beebc2995cff9ab3c78d665421cf2b57e6dcf1de9d5b48209d2d4322bb3ec131a26d29e6320ef837abbc0d1b81651be3adc4f362c8b5dd42c73c5fad8a2a39130d8e1c0a4c2c3b180f129a61629cd51d942b27183d47ff3970a9f5ad0138b19bcdcc838bdd0d58a063b5232fd7efb40f38f1cfa012ec371744012187e5aa7e006b14506ec37ee47d54acad7782673cb5d64b3000270383cf95b6e93f8742bd9d416ff914222cd68ed5d4c225fb2e52b95c1e0b042b0dd18d14ab1e430e3cce051b0bfc3a857fe55622aa773bbaa3cf02192aa0a53f71ffedbb97375d3a89dfd687f0ae1a04807072cff120c6bd962af7aa2fcfb71bf67f7a103f031a36db05578153da272c75c604d9eb48a1a71d685e72fb48940817b3064eea3854cf10806447760fa9f6ebcc82ceca63a3c7241a5d3e9ca922fe61b3f6b577a7019e153e3515ac188678af49b545e210d95b930f86d08ba717f099ebd51dc092399501b94717b1b364c8508a38e79de82c79dc8fe0c1522d65d72ef95b470c2309479ee66b4e544c4dbf0f38f9e88d6a8d02e80d92b8429de97a597c2455c669ae4710b95a03ca76dbf1148c88dc38110bf750002b70e447851f787a0313a26a025b3645190f1e1c4d3cffe08ae9f04266ca5c1d48f266a341a4a3eb6b30323b69792fb7dcedc38458e362346fe480418cdb971cdcb667ce0bdfd6d0c6aaf7145264e0e500ee095f7a6e4896c6ade59d9d66b0c489ee9131408516d98ca4997da75f68f3b48d496a0a877b9998f4313e20cce76b38fc6936228db81cfc4909cd20aeacc3b538a5b468adddf3b0d5d9348f8f8562516bf533b0730db2ea1497884a5415e9b0a44b6827d9bb352e5cbf4a2286652095652ef5e7f1d6607ea115400907fa39cb1302b008d44657ef6a25e86b7a92a8cd9d0f00e60a823b29b775dab7dbd94b6f3922266687e6e8f3203a10064d896695413b5395e0fee9bf2d28ac91fb46a3b2750f71e3a4934ef6d10dc49991e9575fa2a4b0cae5cc69c338477e77bd63fc4c3d05e1d8966858e081d9c60dddc3a80e814e0be5cc02177443ebe5585ae095063acdb76bda3d30420809a516f06f998d992e76406cdacdbc4e990079646d50463c638fd7396919f131bee67f181525f9ba600afc3101e764ae81ce1a82cb3cf61c763f78e4b72e478aa6601fc85cf84eaeb1d342f69d3e57384d94cce260c49d7df6b775e98b293e3c066dc73a499e9d139c6d9cb39d3b1acb72d9865b042bf9761a88671e0c0cd935a6130589ca912872efda3391308af73343e5fcb59ff92edf84a076b7ac640281986aefa467d00b9bfd0c1a1e6b6e4d1b2760671f6e1f6ae13c1d8cd27ae5f34f3bf646436d2c18234636b2135ca7f54a003e56ca20066c06b70e074a7e0c45d1b8c81ecf639e93afd06d6f72d8182ed780d2422b3e7143dff5d66c2f9877422ac49b91b55024045c523ef50725e8cecf6c504329cac3d1b6fce77e7b4aac5ae1ea94ea8656de147afb775cd8533af7a675c3dcbc8ddd925b007c861327e2327c38442aafe764163817befb5863927d7e330de92ff30afbc5074172109ab645a668619e9dedb26f43d836cfa93ff2b4ca252d47a942a3f8434a9bad229b19202554b19bc41cf85aa7e918f42f2c6af615f9c6b8766c6bc7da9ab8b1a93e4cac800237932d31b676fb3f612fb954b5d46992c7d3afe8e7ebd6d463a65d374231dd8953c2374f7c75793ed174e159f73281b9217fd058e307bb7941ec306621ec0e1af941a7616bc67ec93db8a31036105a4209867117b894dcb3dffd9cd2acd17d517d12673e427f379c5383a8244eac603bd56b7bef572d08e9f63eee9c1bddc83ad8a83e2214c474067568535fcb0d26a0194111312553526329d58697602c579cb968e7bcc0bdf51c8f26509e2d69ff92e1b03b26cbe565c70e1058dce9a6560ec1b90f2e20e382a6ed8a626deccaaeec0e55ce48ab13ce3acd02ed31fe8187a43b639e3d26f1d62ec80ff69025485b694a7283410e96750d18283dbb44963e7296e8d8e81d1365ecb0792f9de8326634eee1651bffba1f8ba37895a47726c1d98f676d780e62d937f474b2847484cb08df7403673440958f2aba2733d63c0530ec0832452d2ee8ac2385855749312f86ee01611f3eba8454d0accfbf3af2e7bb1e969d6a22a890df7143d1dcc29cc52c44c0bf0746949f345fbbd9142c0f8dc514d6b375ae43b5cd5f61168a78692d8ad3803ee956ebfc67cd1ff11006a69966c623c40cf0d70d44d33cb245e5050d4d6aedccdfe5054b651522a426b7e259d5d9eed6181b725172294733cbf7f3bf057e0c8e8de03b111545427eabb040959ec966d1d1d2159313e30cf69f509379e2c6c13de7f41769427a23baf71cc1dc7b22309ba4a34a4931e9e5ac95b36f1aecb62bcdefc9f06bed41cc987fc4d165ecc3f27b2d860e60e8b89161225c503769d8eb823de8ba3542bab1f70755563ecd807e9d94ee1bc74b3d47e98d958db3d1460ed7e67948e94e3c885df9ac04191b3b5eb33770db3d22aaa41f8075580f353afe9132616d016bbee72771ab0f49fc6fae282bcfd7580822b882ccbe258a2591672ae8826d0923012c29cd557c4ad68adcd2657a4038998e0cfcef72ae749855c668a3e9f740499247840f5f9c98600ee6a86ffe2fba198140b368553ce15f3b0b2956d6121a24a76b287e191f743d79dc3848e89cb77243b2f33c2b66594271;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h81c7fbcd5faf166c6d14c9eb731f1e4ab57fb69f93e4766ceda6c244e6f7049c0c063c188da81a5b2c51c8ca8f34879587a9c926781a5aa899a12caef0872cb3503b69a4aa06648469facdc69b20c3ed95d397da284fad6d42c086b2ed1747a1f920c233fd28ffd706bc65d86c7ba9c4ba6aa34218e3f0769609e8a570781a77146320987a59b605a44aedcb6a9101927f760cca4b68c47f30e122bbb89e03637df106a84cd7963acf986a482b54ccdecd97709d66b1cc09467dceac1807a5aeccd025965f177c876e3101c4d9714db66d890c12c1130af289b52d00bdfe6eb53e66e4f09b78baf7dd3d4533c8c47c97dfef8b954ccec50d60a42309e8cefe535ec9eafbd870cfc2021d6c48e1ece48cbe9e7af5f5718579accf677ccb0335d632e6d78c0b262e8f7dd6249cb182429122697934d6d298bad750e4de92d121fd81120ab9edf3041e87aa734d13b2e5a57fcbd7a289cea88c66f358148ef593fa79a09cf1f649893a57836b1a1d4afb8b143e519c9dbda1071981b28a7e5f260be82a5bd0f16dd4634a8ff7aaf2e0220a05d623ca17adb6a4c5c508cf5cd52a0cc94442682a45990ccc4bc40504a1a53614f107acecddd3f4a8904c41b240780d3242b0e311dabcf57780c57780b292e0cc6fa4ce185c3db3e21c643fab5ed82436eaa56e394a93522730928a138919a74dd1824f9386b47c1358a04790410d84f9b093eaac0717aa6a348befa7cc20ee2f4cfc2f9ef108374397a3eeea63a18b609865485eea6ce2f9b738bd1ac03a6505f8f86ff0853a0f99ce8f055eb9b1a39fcc379e83de05e2967386a624a347892e5673b8112d0525dfb1003e04859bf13f8ef42b8daa81ee19ce22f88e26848f8c9e10515e02aeccf4f5b81e0543d5dd610729d71e6d0bfe0e3955ca132f587fd85bedd344c7730daa9bf670f55b398bb2ea7b52311fdfc321674263fca5ec56a927e5b60aed88c014f53df29abe879007c6820e5b06e159de12f379fed4c0b4d2572a57c91a9ea546a7b011507c65a4d6ae44a3a4188500d536e90e7be85d94804a9a091709b7eedc5c67cf3fc74e2c315d905ef2af5da8b7e0bcf93df76d23ebaa83624b5341436bbb3ca0c082d213ddaeca73256f887fc985ca9a4b8c3a5ec21fc66c8e9998ca0c594262b20ff48351c92bb9e0201956d26c01708d33f9b96e484c0a771fcf5fc5683e15c3d365ea72674ee7f8562abfea390a8aea1b5ff721f20d96fbefc21e3a329e411f290635b967a8c27e05ba372cdf014ee5df5c49163caba20ae922fa9579ea680ba204bd9c8c3d57f719be2aa60751a7d05cf1c8106a599bee353bc8ab64ac0e2fa958cdc055bc7aa38b36c21900dc4272c1cd42d113c0ff475b13fafdee09a5d6b8df71fa629d756311efb1a6f926d7ce280e2f9defca783fe2316f2b2b01ff2b302dcac49b12146e0a68fb336be075f17ef5d7a4395d6fcd41e074a62d106b620165d861133a7493fb0da11b351b383fffd5f8d2d82a2f9a08cd5b53a88f53b02165b6d092061a12d40041528f6b608a395e1967fdefde62903e37efa8172de9c308d53a315f7b78ed32fa0f8011ee736d222d5caed0e4236dc59acc0e0558fd2ac181fb84721ffcebd71a21db44e229090e5c4441df0865a5fe51f22976d4d3ad7d51dec515f3aba1c56e9815188c018e9cd1ae4cbaa1107c0a83568efe6857c48ba730a9a2bd790296f1b64c8f29300ee22ba94032603b457e21961c203aff22787c51f57ca72bd29266ed98f1a90246ab80fe11a416f054338862490cbde530a4858e4ef48aa42716ba3022383823c1770b424a7a3b6b1f640770106508f2120c457f33f0b9a5e93022c77837bb4da927e1386eaef5422149579512cb0647ed7108ee82b630167caae1af15689930ac35fa1009c3482532881f3ebc8463d213cdb389032578fa6daadbb6873c292607f3a9eb0927b908f69ab5cba96673754b686bf2044214bceee6aff5b259c43809a585e752e89b37e8c8669772bc35cbc43ae479954d9fcd037d2a48503cd323368d689447dcbc6ba016ef5b41f8668e9780915072cf9d0ec3c6b6be418afefcd87da524cdbb7281abb373bdac16c8238df86ace37ce06ff650a57a38a35476da45b5c65ee286c727222b28fe0cba53341470e563c461137eccecf1c877e33de59439892436f4309e123e6acd70046538e500034a70382a9756ddd4fda19a13dd2487e6218a238680b0ecc34ea4495b59d7e2607cb108870b07bceba98ce4d1670d73ec69b310f6fa4125053c5af35f72910586c5940e36223b2cfe674da1b454496167286497bab3e9775f73dd454c98a12cab6c44479144727a7f0df78f2a1eacbd1dcde549d3ddd0a9650bc53e0d2cec2a22c8df17970dafa3249e2683804ebab67914a51f0adc6df2792c263c1eaa5756319ad3f5b2436a074cf558d047ed105c67cdd39c1791dc25e5c35c9dfb4d5fa3eca009153de7c1a6783dc240f1bf58fee09f045312cca01793fa0ed1bbcf3b0fc6cbfb9110300a6fc306b08ab60f9f84b5d4d2865b57a616cd66e307b1427ecf2308d95574a7a25a98cc8a4fff68568137af99b9d87a11e955422a3a33761a33595440a4ca3b927945c70353daf2f59bf8405f34e6bb2af2310d75cd4e9f4ef16335ab5e668270c1afa1542a78b29a341c226c2541efe356f2eab85f8c003790a8950be15a14b391216bec7d00a28f36da1bd6f90ce429e543d34d967344a08cc1370441bcde56721557b064049b54ae74ea889aef4e3af682bd7c26da2b7dfd6d02f097f95c7fc6830f894d7fbf5312f106ee8414f2dab5f8928cbdfad0ca04e2194b473dca45a3bd9cc1debf366e43f4d9ecb14d443df4d03cba596de1deca8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h50bf85fb2f8b80bcbec37a381e7c73ce9e70c64c2ed84b20770d67996b52d50752533a23ea47b36cab15c046ba74d033597517e55abb07ce40f20c9f9c4a7859c6cd1a1b09088574a2969625f15adaafdbbe3f3ba7aae15462e15f5b57faa469078e26c2f22a181717c026680a196739b4cfcac88a7e6064dbec8a9b6314c962f501705424e9b44f599f76f992ae196c74060940710685832fc5edfbf13540308410af19b86f6fe634c90eb883dde3701813d8e1db8b3093c15f2d878695121a490b20d7b7780dd64de3dbfb7a6eeda166ab8ed30efb9cede7db4d541a84823cbeb6cafe48a9b30cf6ddce0a6a9336b13826e32beaf3611ac7b86a22e85234cc9314493cfcd557c33339b710cb0e6da05933224dd4fbb9ed44f5003ac823ea6a4b11a71871338089c73f8275391acd5c344551e3e451178dff046d3965b1f5f9b1c1fa99bac6f83128e2062fdf55585b028ca95ab6689f3a82550bd9489eb7de9d2bb9743178053c55a897da79218f9619c0a0532de63109366441c1f868529a96a3ebe9be5462460686851fa3491699ec40b4ca94e4c7ae09c9d082f0d665cdbb7f26358adfd3c5a6fbbd7c0d55ddb9fc7b3dae919b9512ba3620fbbd1b302d5bd67d2ae95feedd41eff4f716ba891ed2d189bae4987fad3eabc5003e5d5140532aa5b7e6ae2f069f8d8a6795c3a75a418cc206478bec7b736a213044ec941bf93be8b413e795f0860317cf0e042188ae22f7f40a7de50177bf52a5fafe8b389ec76553596735c55dd699d694dcefdadc29c9cacc8927328f08de38d65fcd8154e07ab72fce2b7b1ead2a57667e917fd4c085824b2bbeb8165b67016b6c8aff5b9d957677e2c5599dbb08374b5529388ab26806d06030aa9ff1772e39c4283d893db3d77883bdbeb345e2943bb0fb58cef6e2fe78bdff6b966b2aa04ab3d2174dbac6e10ee783ae368c27abd0112d80f0e71306c8515f24eb91c711c919e47dce4eb5fce8a1b0da1f5b37148cb35cfcf89948d2c028319b0ba8aad4b5da2bd7c10bb523b70db9622f4ed5d2b3a261ef3922bf108f6eeae778cf1423b295dc938fed9ba2ba62a3545c6d7bc0083a883d8afaa45b01bc40ff5a1619eed7ae3610cd7824f0d03b76f5553ab287abbd5b8296592f3509a380985f77bb7dfa349e524e3d9af5a01619d7282e70c5925c3d84996a8cb50feb11f529b59b4b1c27fa1d381d8f4b1f1b11dc02ebd736e7c74fc33cfec0c52167eebdeb943ef3ef11703010106e2c377bfaaf7578b0fa91de3f69a87c30c162383c877c822f14a274d411345a5bb073806dceeb48aee394ee6e37bf675a6fedee039693dd1cdce511eec5858b2238b554c91f42a4765b076eefbd610ed7cbfda76e61e62638ebc43d675622a8bcabd96303e33d2f940b55de337739abbc5d73fe59f257a4cffb9925c0b1e60115ff6a7cb87ccbc4f897706746bb8f5411df01164b01d9d03f480eaa9554240b7a1ab0a330c9a8ac244117a19f268c19d6ad095198f4676e3f6768ad3d0dd6048e249a91f65640bc8a698f02552729e310263f44c7bab9ba61f43337e4f768fef7de3de9905d4cb7d14170e20a9e4f4002d708ff7f81eb834879d9999acb9c97c0e5babc4495fd305cf34a7f6d5a4196b802e742a210fd64b2fe8c53658a9fbfa4c0151a75a3219492e50aae610d3ab98eefda4406b05d6c2a3da7ba49e09f4aa2e03c27a979951a9f2f7b867ed9a0fdf5931a9202075eb056d90b9f5b9676a29c32358982523f5626a3f181e85443f66af7f510e5cf0e64ba5f021bf5d80d88e926d09f4a41bb2675cd45d8c6b6841fd877289446deb4d8070bfba0e030793a8a7ab1a65e4d9c3506e37ab314f3f46fb0f2b49a9eddeea65a3ef26021e6ea6b44993a3492f2559e9b66633410fa1240fd8ce97e24280247a62af95c98def15017a1403e3b5b060891f11ebbfff215788cb56c5f0c5a7b78ba2c1934646944651c5ebcdba73db50d6035f6851ece836378056a1db3eedcb0612e01b6e6fbdca508b207980e59aaca54ee1079f730d94c4bb1f19d63c055cf9361bd1daca3c121ed7b4f572969ca3151fc5909d9094df0ae127dc373244e66106961d94d3a55630c0a871998d2563f5bd26721506ac5a41ef87ef9c55e1fba5fcbd7fbe3bd83a2e6ab7d3a73a40cf4653f37c5acad4e33f83e0bf999941f0753bf793ec13976723bc6949cf0b307e3d4b760ba7e53565ad825eb22e132455ecf9ccb3365dc0e7a738493a5cc6afe926987d64c50f1ff38f437e8d384817f1c27b60146b6e1eb39f5ec49b17d062df5da10a8e3f85162f5d67f9563bf9598a2f552a2bee2c8639b0d5243e984d322103c7185844d8d4db9254e5cbc00ac0aa0be482e3bd3910e22e462b594dcd834466beb60b109a9db8fd3ec16c50b4e4266da7a8857eba8bbd02dbd2fdb56f4e63d7a9fd000431ebd79c3097e7883d00d85fc0f1deb32426369645b387627058acc9860ef79ebac413ad451550a4622cf4d4d5d657abd3c526df76a6a2ff3c83917e75c1a24d31ef7b9c01e4e66fb4699b11303b90763f59aa2e4f812de275dd20100421410c0dc6a1851715f9352a76dc1577106381c879fa37299f1f55c3ec0cbfc2d1da1b672eec1300376ba29bf54fd02843c98a4e9383ce99a583cad8d355f4c8122272e0f55b975acd4a89b08b270908ce8cb0159c6c1d4732e009e714b1408ad726add20252fde1955fb567dd6d8e353d3b433c7c9fa8504c41cc90dff148e5c1c6d3c0b55f91676ed4e9f11d06f65dd64d02781660ff9e6b0915958459b4f126bfa5814ff6e080974be67bc334502a3ad428c6ac6f88f701adf298b58e9971897c144ba9d100550e6f13c6fcbe03d5cea730034;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h97af524b24cdb98c6662b00ae5d777960a18ab3a2f10cf95a83f92366ace9fc8bb85c361fb48bb19b904f9ef4332d1a8f5f68bd1c0d870129fbbb6b9ec951b56b1e77550c8153a033e60f90874b10509a594f5dbaecd991880f75f3faa49c972530a3e51b5066899ed5d570a81be1d76a3720e04ac364e1885ed2448ed134476b4c234b53162bf54454d226f1602b32b45876d5fe323063d3cd986af447be58021db26e401166302f32356d71471d494e14ab5b5a021cff98271cb7a407ac8199e36f3911e2cdb0d1df04c5618902e69fc5249d46ea5510c1bf5f6359f782f211f918d524d2cefc11c2c157e978138c287705e077ed5f56023764c644f0d27666df01a69ee7ee90b7e2a818eb35443a048e0306d77a0374d301f18f23c5c8ec1b0c8792313753b500916a42249673f22bd99d7dd78e7ef9f08df1f6bca4963a29119f494564fd68bd6d6c3ed43b261a30e1008b9eec07a13f662ba4598d8d244cc2a6ef61a8e21ab0d29020ce775a245809f8f88398e8bcf67a2d9e27e9acde8540c228114b0182fb37ab2ed6b15bef9d09759d8269d764f4f11465d14d6726a631e331601d3046b69e32ef0d37715cd184a3aaa6e13b64c0f6b0f71d574f1274dc42bb4b8813de09615099690c1dc9b1c6dbeab0cebab8a557f7db005839b2353f92e5600f12baa6b2c0d64ea350a0fc245061a26a291c5e123bf2b058280dcce09c482f22da2bd9ef233e83916e44f4cdb8ce62d9f466e8409c1ab06ba46e1e2d63415fddae2aa1be894eaed84e48be232cea50d2e4fedd7557fdc83fb5fa999735ab88b554cf3d285304ec21d97c39557be994fbb6b9e1ad5aaceed3f2dd32c3d398d119cd1f374c59259efd16999101253342f70a7324c19622ef580a8fcbf26e454be290f3349cd5931ac8a9c35519090c3007519ceece8028998d319b0cd5bbf2edf6367bdfdd5d9d99d9541acade1479ea5fa0734e60aeda2c1a64f69769bf42f645be6812cdd82a2522ca48665de67b7ccadc92881f50be45c899d187caead096fc645c9df69096034658f1b735619f80f04c7f428e6746b9c8eeaa4110eb70317fea2958051807f9cf18b25324f89e5d2fba1cbddfe7877b67ee31578d556a230db37d6607f7f39867d0c60ecdfa82d07aafcfed66152c99a31c3146f81cc349f182417500733259567ce3491a096f8a074b7d99abe78d7fd796417b70daf28560a6dd55d12d083177abf4ab365c9009e3dfa562792d60a17507d746641dc9b6f08964443c1b15c6320d6da08b809a5f71bc301ff571f35c3583d06a7ca294a98cf0f83ddb7c09980b0a591df30390db5f0b976d0a3cff04b3b2a35b479d0f47cbebe72c87b600523411f875c2d72873aa17226f42486250a33c613c855582384be5597e5021d07a062311ad10258af408401c8438373eb76acacf81b88d3f44bb8448cb7f00f65ffb9117befa8e6c4d94b684b7705c7a1c8d8aeacb6af412018a7f1f80da26cd6baed2aea6c77ff8428a805a4c56494a9fa16e36903eb23f85e9b65e3c068a149bc38a530fb96cf9fdf7e9c8e1dbbfceb4fadd04002a9009f75e7e6d450622f4a50b67d504f050ad338ef01ddaddb60e06d623e51d21749f769d23c23aa37d1ca830e9aa1b46877fb6cccfb5fe87f84e429107ae9a1a85a64c894d6a41ba5fd5fe7a889df6c56bcb7803963b341ae63b79f9ee08383ce9a86a03434fdfdc4b2f5fc2c4cc8c7c3c2d729ff9034b896669bb5323618386dffceefdd5de8bbd7bb0207ef9b4936efa7909f84aeebd3e3c1e42885f28872661097a3b84db343d39578fd214df64191bdc6d6db0d08685f7ebacd2e5c2fdc48202139237b4569f6f79d470803c2106810f007cd6086177391960f43e46f6ebdc4501d5cbc506c0a723c527a23fda0b7170a5a2196b95b9789acfbfb83378cf5d03df045ff28cfd80f8ea6f6606f41370f375aa605748e8167e731085f4311e67e17221c653cc5e9607aacf49c06a80384ddfab6dce7510a7a34043bdcc6feeb636ea8268732c8e2177b840edd76c352f02c11e184e48925ed89db0d93842e87ca1767b4384b74eab0ee5a0c2c731a0d34dab9da479f3a4a8acbeb3c4261b619623358d6b154b9da4922fc31baeab7137de33baad7ba69c2e8aeb626d59238ba58f960e6d1381abaa6512e65ed36bcdfc042080b8d26b2359602ade47537d15fb8e38816bc128a8852a0f3250328288220b687fb4a54976bc3415964a3e8c957eae29307af386533af6cb3b6c9c2f6d472ba0791b427bf9206458fcd89707804d4646126d5317aa4240633661a1354f26a7e00e21276ff84d1d186fe6162034b41209cc1ea887cbc3877c43dd6cf1e661c3206d4fc097d60eec40ba3beb4a12545806fb7b580d46ae9e9b3c4123e297263721089ecb9302eebcc34678669146cefb4857dda80c60fa400bb046d518c1243b0ee74aea7b3c96cbadef92bf5a7985d036ba1a5d12d9a98df02e4c3cdeb4f8c6032404e2d4a935c992a1e466c289be1c1ae21621aab6c6a9cde4f8651aa9a63fc3cb7db0e7414d5f6c6312dc3afc54166e14ea64de979528cd7139b204c620fe5011180f8893205d6da37f4c9a9b966845c9eb28404677755c64e79b51c6fb160c10a03f2ab286c8e7d658d0dbb47d8c647e33c1ddfaebdca98f236616ca9a5709795fd9c5d2a1a72343b48ddbe2916c696ff94f4d4a2717d34c1e9c6919dc829a3cb04a400fe38bac330d3a3744ec04f6c1d0df6fdefcb7a70de05f7fcf4d1743dfcf7ad77f131417295f7d7142c7b12813898d4d98524405193ae69793f2dd753f7fe0057adbdbd313db9cc5f29830682f1c138204d4afe384b7d26287ec6a2ce3ff3a0b6d637dd650b995f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7e68b6e7095e937ff23d89b67edb97a743e096c0bdd5e93435054bca8847a1aafa6fd9fa90c945862395de7a910929d734d9e04037ac1e5ce6e28acf07764a081af524ee84ee5717413ec661c0c09bec359d31711ba16bcf816e9383e8c83b58273b494f3eb39c0c4b6cd12c301dc0166b7aaac20ff2bb6da63ec9d8af2c82621a043cce1c940ad5ff7f44ab958a6a27f581c9d3082e0bd99c396377c9dc69bdb9abea20d568a091720559df90efe8e2172186c7dc1ceeb7e8088430e5aad57cc728c733e20026b87d7219787e34b9849a5d546c94c45d1a30754253a5c6fb1601860df70471fae6c878fed97b21c8d181a6429cc46e196967f2ce7438534196043febbb32d0cd5458233ca012c1c0357ca19148fc40cd68124cca5f2de33c6758be687293a868b78e69699d48310718f06f9f6752c658b85ade8523b2edb66fbe91e9334ca6d9cd78efa2d2785bafeca4ac429104395798e202518cb9858cae913bc8a9c06cd51d9987f67fcbe866d1a89693b75edacd968a8b55f5101fea6d1ff656cf369d4dba211027f82648babb795574d40ccf55fe779b0fc3b001697ed199863e8d19c5911164ec182408d6256af60d4f128b68d5ebc38aa4e9cc5a2ca5d9b5ed6d173b7783c7022a0c420b81b2f17e7808960b60f26b0e130e2cf731e586314b0e3eb537674eef58992819f0f6bd849f8a85113fcbdb6fc8a7510ab8ecf88266c1c60e1fc949cd2b0e7e41d4962237596f6671f7eacf18247ae4a70e1513fa8f25769ede33d8d8332fd806d5ca64d75783a1056425be74f7d3fa779873d9f13cda948a7b69440ed35284480270ef78dd5d994c613023b8f0c1bbfa6a8b83100d4c58b6d87ae20693380404060ca9d9d604c7b2748e8ed8aa63a0081efff9162388dc1441f706b2905af948c1e7f7e9b5de298a3679968149f5c6db478eb3766dfe6df75aa685b41b8d0cc40e681f5c7089205291603dcde32280b00e0790a9d666e22ebf0546c6c72c6e9000e89244574da7316085f9fe4afa7b8162f9dce147b343a5e8f8e2a224fa072a78302c99ec57bc6cd8bd3554370acb5546755819f276aa318f4777adf72c87f507d9670734f2f7d30f63577cf40ddb747a8debe32539cc80da280a9ac418f634acb90968a8a385c603f3f67ac15d01f9a6c6b228a0f1a386517a7931c707ce4ad9e38396379ae386a2427a723df7f807c2c9f0ca95759ac4388d3bc62c34d4865480959c1f111998f0d794bb7c3c039f9811c20455bba2c9debcb01093b93709a551072e9d12fcbca4e2349c3502b4345cade719adadb20876bf3b8164852b6b9c1df29b297ac4a833c49919b1b32683a8635166eb7737e076dc9c0984fa0372eb0d2d8df01a0a6b2c872e9dc59cf6d1482047c5fa7202c1f9898de5cd2c2fb39efcb02ba2022238664ae0100e4e353bd0d4729af8b4184b4c2950ac2e0e3b69ccc43923dc98fa0f711e7bf64806aa6eaeca09b9f2479e3c3105082ff91b20fd36cfd5dd39c3f4192b45b3073696693921a2fd6179d695ec0fced6651dde3c31e25742f16f3be9fd19fa040494d0e1b3e2d6eba6934af417608d9a29285a9c4b28193cd63ef47b2be5d811716fe54d81f00a9c89f1d8febb0d3864463ea18aa0c6d60e5eaaf76376bddb334842cec03c5a63f846898e9e374257d7ff2b336aa30b051d51ce7bde0561fc4c091b6d32dea4a30b700351ecec39dedd3770ee34d6b35ea52f0791c091393dd360f2f3fcbfb06ae06b2b7e5f3ce9ec4d2e26d85ebd74b20e5b0933927d71cea0573acfefa533be833ebff49f123496e2251152c2826aae1e281f444a750d95e8c3fbbedf9fa4db4839a0d9c08c5434bfa3fabbcf7ade2530e736d6a2045c9cc2f1fcecae1efa2836cb797af2dd0d7353136ededbbd5a4502f06bd58f95fdcc9d1cf5f800d51290ef9bbe3ecaad778aededeb9d95873fbc3b3e17331fd610816e3270c17cdadcfbd002f407fe9ea8d05e88b7602f28bf4a2a7910dba89aafee0b896e71db836a8693b5e150673001e9d71c053cbd313b67b269e0dbad5ab5dfbcf9d986ab32ce2052619975539a32cf982034d547dc97bc296af4d6f50e342d0064525eacb30805fd1d3b0f134562110f9042d2a4263d54f50f7714d87ed151c3b1dfa697a90640a515041cbedf63458767d03c5f08329c5c069772ac97b21fa204bcbdb7c34cf8c51e5b76a9a6bb50580681576229d239e36fac5b5bf37fce6c6040f1e0332694f41c1a596edef72c9398b09e0d9ab32dc34eb3200cf8e5ce528e640b6af0cab45d9fe6c4f7db39b2bb2f2d882d3e862af2b2923567a9c2535d722e17b9005292cafd96a4c6691aede28012cdbdae6c04d417a26cb81237e2abf4f43d09cca4ed99bdf5ac5fdf657a494132d447fc91f04d3f597dbef74aa7558d8b31b808f65e3bcdfc4fe47d59493e2de538697dd152648ffd16812d7e5d80ceede7f334ed9181c5ec9de8fb88aaf574179ff1b14a1d0965e7174b87e92d5b8eb87c73789fb29db91114d8b95a18e85b587f0c100a7f4993b2d82e6ec2f57df3bda74abf58c911e92e5eb44546110f09a36b9e97d734cda08d6ceed958dd25f0432e1095edadce18d1315b22b566d0ea7b46cf2926a124497bd1b42e797eecfc84b5569e27f6046772ff3794a4b55dba87618a2a7b189d45ba13c88d7f15c287b8ac115debd48a4eb636cd537981d8ed6538e2363cc078207e2149f63afc0ff95be54cdd2225ca01456bfe930ceefd380f0e98feba7963265907a4108144fbc130cd326e633d2a48a670645ed94e9de2fd87d124dd9060a57f187e6e1cb472faf889da8b764c15cf38f85b5bb0cfd0eff56a2d806c135d3fad993d12129a6811de8028c8fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h16100f4490d1b894a6e4d2366a860e85e8e6b118fb3b6136cfa9b02d67436edcaae4a9a241896d54cde05fd3365f61843cda04776ba3c4c5a054087d53caa2ac88d8057c3ff88d00918b607f6f26e0c6c8ead3a01d2fbe4c70ea8d1cdaa2637bd5ab203da73d42fa07377cf8ba86dea775c987f4ba77976e7e48bb537cb42922ed2d23b7c7363cb8aeca9bd5888385a8af7af34572cad5aa3723f247ce65e15e100e9aca632f734697465828d837eb72160c4e4b900d39da193c6b65dd34e29031ce2e7c133d71b48a4fc5234e7e02c8cba9fb660626cd39934a7a2b9961555fca3d89aa50be532d2b136e4a957942f4a8f4778d8e82a90940dd22a57bf0a8b8aa31287e4e57f8e4725824756d0dc24e198650468655ba1428d26c6e286b067c0aaacc0b68eba440a36265ca943564e4dbf7ff5992c589192a49e8b1009bade0ef43a8be60e1612a4e563f01ba58e856d33c3aa07c24ec060e740ee7263ab3141ee66a4a68b824241af959db9e431aede6b78b6943baef4dddecf5f0a1975226784eb091b6fe6269e16400747760b04c79bca9801ed7f3ebbfb1742684ee511be77f045243a68b8a8ca7da9c5985bf502bd02e62ad9c594dfb350b630fab22f9b1e3000044efca80835fd09adcaad78d71d01c1a0f9216b25bf79440099872d82b9ce39b6e91eea26c59cda5bea90022cae6c2ee8b84d92e1cf18ca288b5ba7e21505db58f9ebef2b7b5a404a676c37bea99306755ae4d31e75e260aac9954406ce4f8b8c9d18e74309566ec053ce14746471b1a36770c4fb60c4da3b59e8ab647198a0ed81c8160039d120b39375ba5237f5bd412bbd25c9cbb5f408293a970485bbb5e2436217aef66320289b2e6b191835eae17c4e49c0f175da50963c9d1d37436828f5e84fdbbee8f596f2b9c536471ff23c63c67c84db4fb259d293f7753759c1e5ed4f1c653c0f517e3de6a878528f3ce33b58c986a1e3e1218fd1dfc6bc5f8461f1da5922895681a9fd8c0bacf0a480fa1c1fd86c3531d7a496782358378722cd5964e6ac28c83cb7ace43d8929a59c544d0577f07cf316a44475e30fc8198866debb02868e7829855dc66cfda292ac533bb8469284e00659839d1125a17ca2a2410e5a152d87d8bbf58752aad4217b6f8d81fb8b3acabdcf90ace008e823a0581f528a7a4d7ece80e0dd4335d9e005bdfd46facf9c1abcaa454705ef1b75cf0e03a5668e39d045c8f0375094a3ad8d50c66d608aead7dd2e636fa2bfbeb26b64b9bd039ddba62883566545a04a8a09331a6f74a58790b4ecd02708dafad9ac47b4fd2fde3d2831946a0f4ea618b86dbf6d2bcf62f16753f59aa7a3e72bce3959fe6903aa0479625a533746f81b109a3290cb21bbb0d4f65319d59fccc6efc942b2f438efc7e5293697a0ed182ee5323c27314f0ac973ae91cb81793896bcfd2275ead610faa71cb8ba2c97cce01347675b52d3a755b38a6d999040fd16101d4fca83d4638bb83846d30203c7753454e080a518bcdef76ef6c3c63e9512270393e0e30d7c4cb8c29e8d81fd14d45deed4e159835b720a795741db6022e899d2d67d9a0834a7e0a5ec870108835d32f1c02517a2df715cd3e76319c44eb43fad0d545c3b7e4c98400c20ba69cd934c2c009231712e346f672fbff36b47508b882d99e86c3ba40928ac6c8ba8a38f14abdee487a45186ec64584c8d43f67515cd917292ea618b05e6658497d0ab808d1a8bb8c7041630578f18140d93dbdd11e2efd94d7c490a4305463e0def81507f9ef287fe090cee62820363594400e622703f63c0c79961ecc98320154b0b554b01d38b93dc12afd52c2e863a15d29861b67ef60de7092a394db1211258ee954c001dd85435b7431c5c84c7bcf41f162817eb5808e5d374fe5962cd737d535bcc3e53964da3756dc5aba98a6ac02a027b1adb7e14996ff5a5c0711a6640618621d39fd5c2c91b5af4d17307bfa0615f61cbb421659133f40d70233522510ff2017152572363ecb703685c331ffdfc41cf6cd028a289a34c9bdfea70a82844edb608864c2c2993901a5710842d2e9601ee5b66503b0a07c47055d6f752fd23234410eadf065705f05b58277ab5e1fc221da765299ab6a5a1619c23de3ded934b5c1dc29da5b03492b1943945296691b320b21c973c7c27b64d072796c12c829ad11e9e0ad28afb63674ed00f993d85fb062675fc3dba0b966c3464a57f980e8faa4886e864978375830ecb9d0da291181044a1fb017c9f480108cf73339b9d8f8f651e0e9f4a260919ff7cbfa87eb9121cb11a876583750782b8e512486ffd66bf592621b72f9278f262b2ed0bcddafe08660de2676e276553ef9e29755e142d72c5a2c0c714fc6ecaf2f88ac06ef6a490925776600d04aea0fba58bc77e12dca922894d8dac31187f6c88d95b440c33d2cb1e0a9a2b37daa4e711b3d7df24ee91bb14822079c4d5d0ac72804c5dcdfa70bdc3af51ed81829505b94f9c4968107087c0ebba59d53293ee6398d47f85f73b884ee2db225130d860acccc4183de3d80ab5c47689e2ee722dad57fd99b9d7c26b27d9076827490d62c04fb650b2a9c9f4ba8a99a71a98a3187ef5df1238b1bfea75777a39b82976551d9bbf6ccf16cb699e1280be8bbd123269fc01de7e0aabb9f438400169a33815d94482ff6c6aca0a8c0ccb7da7024667da792cdf38d0e7fd84c2e09f9439dad72fd8ee7a75f800c67ef65bb37c931747795b9b26993b1c36f18e0288783219c0763d65c36598eccdf2e65d92ad14ce383aa56908f8d53b59186c4a8a21aff22069446a4f42a9e60ae720674a361245a1125502ebeb65599fa70c99c2240a0d13177847372e8b56537e9c25328310082c72bb7ebd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5c4fc3c839058320fb86a6cae13a1174118fe9d0b8f483152ad131a0bc673da6312b7c271260ccb00e5fed9287b99c5ebf33a7eefdb6e3ca739a42b2ca87216e61e4d2a3b1f7dd93e0a6dc4935f5a78c719e40196181ea575bed7cc06b937e1820fcd10bdc9bb769aa1f419e86bdad7ae2b9198c5338794aa23e9973d17d0175fed6fc76d13e4ce3fdb2db6b394a8d7adce26ec6d6e406311f6a6c5062c880fbf064906b6ea5058ab56dfb2fcc717000567730f95d1cdcc60a9a271fb1e0e30ce1b4aeb6019eb0cd858d2dc08498eca3d2486ff701971be53bbcbf1b315b72e6f8b2e03ff0b2c383bbc5293d98e81950e64a60dbf121ddd0deefc57f5965576f29e5b989e753bac32f7888969121b21484c72fd1a0c991a9c0e16f265f0ab9b8184bae37161464ef9baa91e1c34bd6c97379e1a1b118e2861749c8b44d2a720b5a22b71545c1fed3e306b4da04a20679dafaf39edfcd80a2cb45a4e5601cdf6535ce0a93abf2579170cdba58b3ce5c410ad8ffc5a9ca6b5ac872922de0499830785c78969876edd8fe3be885575e7a23c71c024fd5d45a8d4b108419f9703daa5fb69398b7634e6411a35ec1d3a0fc320db5e2340801fa9caf2336dfc5173a501a759e2acf325f88cda3631793b2976652908b220704b3a1e952672d8c72d7ddbfe32d1a604bf31e33a3851907e39df1c6c23457c67bbad31876a3327900f58d7765e3a23c6b3a80705e28d02d69f29864196e235efada4526e703da8c37ff08299d284878c2ade0618ae1e6b32a58c70cde4bbf49875cddcfd25bf2cc5892afaac9d5146cd2f13d5420d9c45caeecad6b77faffbde78b5d08e864e99464667eb8c56ac2736686adf00d5053b9db5b5925c309499f1587bb1f73ebe9445dd3fdfbb751ddaf1dada09d9cbd4511389a97bddc35bf3f79773e274dc6625908f1ad59c4bcab12038ada04131da6ced114ffa6afb9d2917a23886fd221039a446fcc15df00c98bfe0b4dcca9411e69bbad6da7721746e5304ef93645936a5200ebb4608e8f545a97cc8438d01fb6ad6d20124c9c33bc2f2f1827da13e04643af06536c83b6eae64fe6e2fc2b61bd0664ead3f0329b28f2965af31e3216028bae1e06e444cea220449820cb29921424e39605159210e66ce21e694e2ace38e55e6021d0ebe36866a96e629ca68f80dd7a8e3ee5dfb48fcb514dc1edac71b736224775b9c3b39d92ec82786326fa9a0d2c908ab0731304e2e730f71fb30fa4d33d9f594d4b38ed058a21996dc938c1c86eaf1ab10898df75f891439eee32819b1008486a999e6df97caf019688cfb4e0ce29c131060e431111b003fc8058ba69fed92e27ad7c121d1bd9a94a8ec8941a8d65a8489e3981cde2eca2b138eb0fa9ba02aacb1e4284fe9879911033dbf3482f5b44f53b9a783ade2f970614828f03a418ded2dc3bae6d6de7100527d1f3c069ddab44fa03bbc79a28ebd46b5f797f604c11c7ad97265089ba4b2e83de710cf916fa1e2ab9ff51ebbac9cdd5a606be31fceaba97c5fffe9fda79b9e17783bdb6fb6780bdc75ddfc6805be02ea5e59ad102274145878cf8cdfe0a06ba166d02a3ec4eec3a00110d53b8bc13dd8d3a22dd53972ef409928e4772c4f7c873481b37f9e28b4695e202abd12b7ec8182e3b93804e1f985352867ab5e8fc33ccd4d6fa651867ed21d22ca45266a7f3444b0ca18e0bc0d9d47911906dd1b67f11ba5824ee2655fea675ee5faf228a544975c53357ad1d28d5f729446e5dad829ea5bb7cf415ba03a0c8e556b7aadd5d7c07eed0e0ac1d9887f6259660d8fc0c8098f17854324c5d7b45c257def15249d6a2b61dfe89ac1e4081c27af8396448c9e78e01c211b3b41b8479ce9dd700e86336bf9d19d301fcc88b247436332e9b14126af435e560b1b53cb5e2b4f1df7a3b82b3a3f85ce7b52e627964cf9a766d5f66824613081ddc48cd97810994dc8bc0dc7f5c51e401548e0f1527cd8bfd8566faf5cb789e22151174e513f5e958ef6c8b5a952e2be3e948a6e6e05775c6ee1aba152dd549dd385345b3e8ecc26772266653bf82402abe0ee61ea5e2a48cd8a099b8b3d06e2f2c8b6b30e75c56f825f2a0c0c03d8afa039715a41254b67d5a176fe7d1a07be38ec72a99ef977ca76a896c8c2b550d25e77b541a33ad240784ca1266183c70f5eafac0f2a2b55a567c6daa9915ab97ed99caaa3155b13aef236f0f5176688497de03ef92962a94d66ee715be05a97707dd6aaafe135bc7823894643b9ccf2d1e5f3bd756385246f742f02fe03c824a8f6f89637a49ee7413ea62f3d5c6098df13ffc6410e2e2c60bd8f6b4b28174f5068d465c324f8de33bfea8b7cb4ea983560022a3394b7b33a016438ce0c25990740f6a11fd35d8637e8103afae4da850749613fd6e841af3cb581df9b5de4589e8dafa9bae552cbed4af0e9df36b683f7b7d67bb1fd49e436bfc23b402dee267424cf102f2007a1656155b7b22c8daa68f2e9e31fa372cad31d669197604992c9927ec07e9e5427c78e040ea61a300092c28a6f09e56889d8feb9307fd0a629c6b4c0f8f3470c6c7b0bc6d11a64e40d44ac018baaec2d9980ba133c4ff05fa36c43225e3aee5454c5e9b1ef446afd875c5ccbfaf3bac619a4dac89b7f5ff7eb757fa90641c42f1ca4fb589b6a38ec0b59bad6014b86677449253acc6fa95ead42186b468c0eeb02c9a427471822b374f9187efe1a2ef4e30185a9de9387492925becde9e3732d0f0502caf2668fcd3e56747d4cf9b76acbf4f27f0764bee7fac26f32a8ae7b5841d1fa97fef52cddc48526dcf0bed797821fb8acb426c164ee2d7203e271c2c44926c668932afa62afaae24dbd5f2bcc724f2c0b6e01e279fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'haedf4a103aa1fadb7f2f57d51392f8496ef764447aaa89021ecf7702d47d649cfa92a1bd904cc5cf7733d3122daaf18e794aec3c9f946f645e8084f66e7e9e2a83ca0b985580ad98e658e505d15f587dbfc27a83cb0da9991c6db4ff65e9dbc141d58295f75a2d5da55b4773dcee3c54b81ff01bd60225fc1adf4da48472052f2b42ea920e190ccd3199d140333d26270668edc72474d4084a8421dac68efb23c0df86e1f075f4dce8a2105fd8d0cbcbf41d18a1d4f03a5271caab062a3bb197242db3c354c38fa3cee0a736cf4925c27aeb616ffa132d1c72940f0bc8ed768d395a4ee4c0efc8a693dbe5d866f11b0155389c56f7c7fdb0405699188f36ff3dd3810a8f4d0ce1c0050c21c246a5f04d5ea846e696b26b2f2105cd4d3f9648114b08b913107eb2e2aa1599b1da831f95304d8ca5b0ab7af451441a1a43d6baa2db5bd2e55e055c04cc4345d0094311d308251a5e0d89a1845a7fad20273d7aa404042c0684b2d095cc3bfca1d9ecffda7099d99fa88d25350a8ea7843bd6e12d3d92daf6ef59abbd10ca56811bf1e8bb788b2656966043cd0e3776b24de20bd4b03fc0e5db7e8ceff92d1b2c8d152cdf217940aa5c59ac20a7b376b272d06d9717d77193af1303ef61c5005e0131f6d85231673fdc6ea0e7a558bf4e21c22542ab4d23c696bcac0a3aa752e3233ad7f69604d8a7c432f8ca6ad4241336917deef26d65dfcb85f329b74958ea261401cac3f668a5a9d365377f9d4cdc8f965e97a2249a945efcea49995276b9835f5822968327a5afd04d59b14487255096a99b8b739e56b6e4eb606e7fb5d94261e9660afd83362b7261d452a3e0ed627fd2e0698eac050ac8640ebc5710fa06fe3e4c2d18b5276d80370be748a7e0d169e4163d2ee1b6718ae16e920e7a2ea38d394cd22e6edcba15cc63ddcc05417617699faaa77d8cdda64a06816fd97451b8c10aa14c24c5b5200d2506fd8f2c3ef52fd55e1d86a5ffdeb8fec75a380affd4d2443b0772dd6ddef8d0ce138bf285181595dbbfd6252d5cd39b195ff086f59e9d714d8992e44d15a0498307839abbc2a29ffa7f42cc5de39761820a0c1fdd7ac73f572ea8bf1b3e9c7ec940339ff880a06bc136d9183b78df49708cf0ff8be8b018d13227c5cd354d68d8af84361d6473155617d9e7a42e7955201a962fa8784b915e5eb8b5d8ca5c142af265c1fd2f01d0846a56fcb18a6c26fa657628f55f9e47241cf2baab600e09bd16cea2948a2d41872895974d4df942fc01302b39c09991b8fcb7b2137bd5391ca516fac454b49bd03ced23c02159329d0991c5a60e8ea06b900ade6f545e3ce8ee4d7a10b8bc921426b07eac0876e1a8f41e9c2c5edf1d46c0bf74b5ee36a5cee85f493b24c11d98645fab8f6636639a986386d869848690a4cea9925280c5634b5111e01eb9fc5f047b5fc6f45ee43e27b01317e7e50c7dcf79ac1d4a7c0f8d3998380cb44325488dcdfbea7f109359f97e70e45661f7ab1e6268de40a0938ccd5e4a006ea7e905e8022091de99ae16539661a829bc78d4aa6613abd7092f8f88760451602f95e7f9bbd1d74f2d678566ae3c3140eca323f9f13cf4307cff2a35c462bfa093fa3b0bd50ec4169adb7f69f73749d39bce5f9b976c1d7b85015a0ec5f217d126dda927dc3876267dc99f013929f4935eb68404d38e60b3ead0440eb7d9632ffa560ffefba83dde0e15c01cc08d64486ee45926da02c463dc359256822912ae1af6255a0f6351a0e2c733159907fee9c01e57de54d5d4c9026494150c3a78b8c269162e97ee42ae58caa2d468e49b54a8456ed6f5a8a1619fa386aa89752fd70f51aa6f00e95499a0eacd9677ee92e34ebc8b0816fb02fb1235f53b4a178ffc803f2aee7bc7ea7d7a8bba878c80450540f42da57de0198744b167ba919364942483987628ad6651e465d73f05e2c229a063716c805374ca5f6e910d81ecd09c667f76d6652be5f7122a6bd5a118b9361e716359e9f973688b364a141fed0e1ec6283b103ba68100168d1fd656c9b16b8b91783ee812c8e65e9a2ec648d3beb8b95ec4e357c35524ba4a1b7ec4f4dbb6a38b7473479dbd1b996330ffa4191fad0fb1eeaa234054279731206645e09e4927edbb7fa864f5c4e30142d5afd397178522130f50ed8985ec079f1b041078a9ac4aa1f24055adeb3692052225c35ecdb76bf91bbf4d6fc02aad39ad5f0308b62290614c5a1f9e4af2b2c24e1175c6c0816f2e939e9371c5f288e890ed51ad3c5c7ac8e171260ac2342eca55833b54bffa135360a1073471cb686049873ed967e428385e0e4c50c87160e68336df4f1c88a7fe12f32e9108207ab2b19ec7a38f0f42b0e18bdc1f203b6ebf077d3f512ce123c47dfb934317d04be44927ba7c9605a5abd206504267d5baa0d1c83f6533acb0b838fe92cce24db76986b5efb430538f1093141a8d6b1defc51f7536b521edcab87178ba6aa42c0f3946745b2679f177898d31bd18973c0229d63adf148e6a3e52c0ea07729a86b7ef3d51d2445310c57d0e4456f4c6a66af8a641b6fe42dc6f708fc5f85ec1c077d7256313b47b1e1514ff1b20ea23d27fd31c58c88091634581c0cd3e6a0daf7023721a0ce1e798d4f256180279fbfe48ff9fd8ccef8e46caab52f854a0a03882b78a0fcb8f37c1a5be00e181308bbd1588a51983a94aa6cfe228a0fb2cf666f17e067df1a9d45f31bc7926ffe04f6005588311736bdc27387fdfda70d4ab1a669f60f8344ff9f71ad5910299905a090061064cdd79972d2472098ab8136b288e0d8f105e2a94eadf0e0aa6c8926223328313f578d75f4fdefdea792c43c54a0157e068e9f29909c03fca531b5327c782090c7fe166a960a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h30acec00427b964e4021cb1d70267d31927cdd4e7635ada62d8ef9cbb88ade89e4a89719a13ce47c88243be2bf58461fa5732d4bdba95a8b45314fbd517b5abd2fbc17a935f1d194bb63014af8a26539b169afa97df2fa746bd04624a09e1d9834e1e28df20919dbd0249994a7e54aa5f1d65f2a375a64ae6f49c708e536034aafb68712c2f27beea2605576c290eaf2d5a4d2be739d16d8106568b238f3ff568ea0c4dbc053ce0c8588a49dfe5752d72ff7c07888ded5c51c58d89677c6f92582c4a8977b05fd4931e5d77c946dc0de9eaad169d885ef769f1477240ac37dc1e86c39b88ff9cc7a6a90cbe0572741e4a45baeffdfe23778d60aa392a168fdf2ac6d7a13eceb408dd7c0ae24f76fb36f766400b2b9b73378229891a9304c036162d847912dfed0061bb9210469796a06b26a932238606f3db913f61625055a226c18e303e580d8873a572320eac79aec00437cd29b9059d0712b29b91bc5d59b6ba046500093f07aad3477cfbfb68ccd29b8c1aff5bce9bc507587a2be1de8f1a1fe6bdbc76569e2a7813db38db1650ed46ebb2d2b72f8e075576a10a6e9439bd80dbea2021b6511b8ba65738c8e878b54f8db281c6e036e8e67655b314120a53d648375c608963eed39d4be5137fc541f91823b0e92aaf599d43217cc484895a073c31ad120f068d335aed3f96451ae646a20e8561739a6599b744540db130d62071ca797098e66e6765cd01a36ad71a798913713a6cd16a26c1fb6fe661c4c25d3c378fc3433c1e617157694e3754970925186c5d8714da1241b895242d83c9f9f887c6a8a54357fcb81960b236124ad702de53dc1e33899ee01b1d71c1355c3f8629ff4607a4d7c66bbd110db555cbd99f690cedf18f63199154040f271f9b4029806a433b8755e7482fd1f80421bcab8ab1598828e6a8e24ef6cfacde9804d3d60f29a7ac7f8b1d31bd2045bdd1d161cc87716b29a8a312ce3e61100b8c76b63cbc7887f8331f2b37ab00444a5105a897a3d57c82c35e5c7f5b745c53789654fba1de9eb8fc9287f80ff37f650e9870c17bc623d69e5551695637d7b869b8d722223092a60abc904d25d1c411bfe5131c1da3f416c99d0976c82cffeaf018ad6f0f97c68bd00bbee91c0ee731b207fbaa155219a7bd99e3e155db5222146acc8670ac67a74974d9da63d4c4a0576abf628e36ae91ac3838617fab3628357851e6bcdf5138f7e61ae18a07710feb82e62dd9eaca638393ad878fa6b65cc370ad6f0889846c06790dda2f138ccd459a4a6f614e067ef61e29e978885df9a1bbc97a1e539fc59fcd15f561eea0f30703a860946d2069fb693a733ac6592b573e85398125a2166c5a9e5c2c484da98ca872ce713663f2650f288eb86ede7b00b93610106fc18fd6f86860e406e6e3bbec7da729b125a406d959b82fde3a9649993675d5f4994fde37145629dc129ab4e8a828694dca92712b91b7fa481dc627fb950fd0557869b7abdb5699d25288af286707c31103a4bc81d1febf4116e361f26172c58b9dabefa12e7cc837e7e5d9792598f74ada7a7ee0b5d4e264edc1f646f87bf8fd3ea56401e383763433b0e4c2cec1832ac79127dc3502226e046d6b6e1740c7ec065c7382eee3ffb03dba9a577d8970a1412b747d03d89fb1045ec61318b1280ca8b34f1bd18ed9e4dbb45ecf344c1c34110c30d16f400a5ee1272a7bf80322761348ff79b764f8942faef672a5845267f9f892e52c506a3a23489914b5c4f6bf838554513af7fb2a4a425171559b149d38c2244e350a0924137beb78660f7e936a8c2231b2c7c827b3bc8c1493157be3af027bd24f2dd02134f989d73db07d4d49a335848f8db28007324f35669e5828a7227f2d54fe83f74e204560355922a46f17f3507748fe7f51260a5dff62f4428ff656f059435e17e55436bc798b7eef571a8beb9eff96bab6f715de07a8fd509db3d359f5d015b3f5efb19edb44f714748fa224d5d53ac5a9203656a691db0e5779da4d977ea62b850d4fd6e4d698aced336ac9dfcb14b6b3a04c5ea421012e36a21e903d835eddbb51bc9dc151f6acb4e87c2bd997dfa4504e39d6f24b7db03d167a25831595ad1694360323cfe566ac29017508cb073aee51c02ab1b7413fbd48f9ac64c333f687afb24fd34748048bd480661d272a8aa3bfac450daf0dfd0469a854f08afc173f297f03d100325f125e199b3920dac4be330d3ce8fd5be479c08421d7e638a1136fae182c92620afb93784390936801084c2d580eb288ec3e6f2a3cddedb834cff24b5c3d2669373a9d7038393eaea5151eed48926f80596fd17c457a31b7761030126148ec732ccc6c00178962e4689ffb38146d58b6a28145416ea38e5efbc5e9fe78c3ca04d052368250928f88dd40b6ba98683472c60173bf60d0fabf6f2d278faba53f7c7b7600e404e0042c494c7d59b6167994b0ede5b5c6b2cbd9f414faa52e90fa57e126d8fa596df9229d34452c87e2e79820da1cd2d217906887b85f7dd21cc33914bec8c0edcd43d9ad16d0b6ffe44ff7419ac1d4225d7ab56dd2f7e2793b82bc760fc43e472ad3817a80f282b24891c3730583d2f88575cbfd37557562144ff0adb83310e21f6ef74110f2d851ba113529e8ff58e254f525fea2086f60f767b998172e270c7a5c8f0a90d1a0dd86d957ef7ad88dbf9038a15f75d8451a51ac18efdb1953a4603936bdd9367a5181db4778b06e1acba379db1ec62f60105f385d619564b1184fabc17da6b007727883fd485c7d959d6abff831432d099c36640e21f888e25aab632a76d7c6d7d10eaec065e676cd51d3083f8c9aee2b8d99a527d0d158f665637271551a8271ff8c3c84725a07b1046d970e1e29ec851;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9fd563be28fc86d818f027a0a0532b9a2ea81a9a28b2d91c91fce207d62bae2e1aa6734e4c7d67547fed1d86314e02e510d263ae37ba80d518730a73ecc0368ea3fef40ed6b9bb4fa1298733061d3aefa5df44b6b85939d9c433f29a06447d134ad1f536ff2eb6168b516d783d0ce36a0befb637aa5d3cba0d1c945257b51d4f551599d180c458c7e7db0d7e0870dd475225693efbb6778df25bba8ac64e3588b1142f36117c876b3843020c0dad88ffc99158b96cd0c086def8d41cfb7375bec3246d4ac747a1c9474b9b916755dad82db30bc0591f7379c546338d085974850eca83935c46201cc8106cc8e68226f61919e21e99e41483d03e199903418d921a261e818d2cf7c8970ed3149fb4b9931a68cc4399c1d1e8aa73ded686dc7a70a0472e27884ae251269f1a236caded52cce9621607ae12356633b1511753f61363d854bc3bea3a30f7d0c04bdee12992c8fa69a022d6d066ca1c6fa12608ba189567f10dc4a6f2af061be432860e4ab75d83771ffe7bf37d1533bf2066c4c759656d9e086db9dca93a22052b73dde80018644299130840ecc174a4d054a7c00ea50ffcaa089875ee9505d31c28a1919ecac917fd9c04b7188558178ea176232e539660e7dbe6b878d5bcccda4181044aa30a5071f49760051f4079dc698590a9cc5674efbab2561d3736a61135bad8ad27f487f2a1e8bdc2fe90cf6f43563ac889c53ff1e7f5c0fddc6fd8c0226d3887c76a06a2f4e002e3919440ee8d25aeb54e8aed4aa9faf3d91b073b6a68acc6e1bc0cc285d2521a50cdc1a3d1f80aed50ebb1c737257077e3b2734fdc6e039443d43053c225aa98bd1c5a2ca947c1b4f81d7ea116624c8cfc1e9a8a4778e5ddc22555ef4b0361214a90362a731ce7cbb15bac0b6d3ef87c5c84366a5ac3bba817823641219f9822e5316cac62a7e936a2c306605d6c5f277972354a7cb1f17b76dff9b4485e7792c73d441e3ed5b1afde7ebf1295f95a3329d8bf9d8abf2b08398d7ae3ab6e6fbd92cb0a50528d554cc9ef31e60450fa15daa9b447347fdcc2bdfccb9d276690d35e04fdc864d7e4e5dcec17b0da0732d4ca20106028921d1b94bd7087cd6143a0ea8e1efe27fce3340002f13966673bfe08ec8658e031765f33be7bbbf536d46b80a05f0945c5b99bd7663384d96455633375be864b2cf2f9d4370037b8d8195d7227d29c414d241d4d3b6f6fe83588cf910adda1ac9a0c27a1d89820df327059b45f0a865a9fdd3055ef75ab09e59cc965a59557b8050ed6e9717b1b8355697bd0c6d5d9acbb32b4049b87259d2571580bf6d486f93193be7b93222c800227b6f7cbe6565f82b05af07b7ff9df7527a4160911b12be964aa30410073fc97eb011030828b9af66d13bc04d53e04fe6e616c1cd797c1e1f6ad29d92f2e75dd039cea5e2dccc4529dff9b2ea889ff16bfdceb361509fa8c20133505f9e397af4d591f8255080c7263b71da7197d199b587a9f1894e41adb1356d29d1946f2d7bf28835d98ca18f332347575fae3b02d73798514197ecdc6347c546d183fb5b7a3bca86067baa18536e6183bab15e9aec3fc387a65f9e63d54250f004cb04746bbbbfcb5d9ce5aed092d4925bc2019b13e1b21936c7ac3d534c69a60704655435a6b4e5dfdc55f74ac71fc02db856eb1dfbefbc85b24f2f4f039a02e94649a9c4e61f98e0b96abaad353a138ca76665b774db6901537f74aba17776cd4b25d88b4a2ed1ecc30a9724d3203da1a8ceb3c560831dca845540748a55c10196136335e440c5bc9fd02031d86ac40f761804cbf2f971ffcad0883115f374d740654ae580a29f3608aeb98ceec9e153b861bf8dd7b7cbacf47e8b68f524e3dea6eb55060e780d9cc785824f63cd7d2b1880b2e0f829112a9425131748730761d41f15a72bb7736c8a26aa43da35fe38b1077bab4527fc995da58d0e24d95cff6cffa71ef40c722ab6321c9db3d1d7096c56dd83a9cf6c6aa23ec5118266d1ec38d7b4a30f89da2e3448b4a8fdcc56c85d04d6099fe88774a8f4881fffc0567e75967f1cae6b6f11f6cb0f37a4ba13cf418ab03adc8bcd0440cb7d8b05cfa09e2ee3effbc54a5668a802205263ca85a8adebe11be70ca2c912a30558cb612de2557ab6a168a8c3a7f5ba0083cae20d876ef1a63357125ff19a52de1620a0e9d5989dfe198b49fdec7c60eceb3ba9d18a8f764638dc0e29b662b4b989ecc8343573e12031f9d81c3e07a2fc3c4b271ea10101f1f2a7f610e48a818d56b0d9957a26604315595213231b8afb51232d8a0ebfb13046ecebcbf3bfcfaf33042fe18eeefe7ee83e10828d2b5de11dc2647fe3aabfc1521f61a32db103e2bfe12e543f189ab7e2cfdcdea44f7961254cdaeb6a8bebc568b56931bacd6f70440600a5c0ce54b8298d5f03f2019c3c4226c8f9b5e9e34f586e3fc3f16a7ef48f0d2ca1110959f3ca2c374ef2b3befef940cf94efa674411b99aeb17d1aa795074c7f865cc042744f277367b8c017e1d9330964b37191b0195b8b81bb29f302e692cf8e32e9dfe14ed7a107e4c7f3d23af44abfcc5f242ae88c3a7cbdb4b967ce3f24f7fa308099638ddc6a77b29b016fe77365decb80f208cb2e94d185332fee86afc3a41fc2823de849683596c0e83452a99040a7f488e61ba7e3ac53be315162ce2f65c0654a5f524c5cf84b570786b9577284c8e7cdc610cdfe86964361010f81c6ff1c8639f448e59523b1a7b6687a24fb355c73e4536be142b4992350ac9710fe42f4716c396bff66db937eb707b3b82543e0a37b93d9c52baa1076612edd2234c2d88867d27c56db568e5d7f5c1cca4bb4e4736a70d34069d154713115d61956391cbeaabfff3f0adc09bc23c05fff1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8505e4ff30078824d1d0fe3c3fc7637702463e8d1db59443967bd0c7873ca9623bd6725ac5544adb9fb8f702d750c7dd505819911eb85d31a360db4bdb362626a15f9874f3a5c92d0f46dbbd488ac0aff7c3496d9ac685caab69e4cb827e2c26208d7234bf2f75c7ae79a8e2fc5b9def9221896060a0f2476b2b803606555db64e1013e12506549e0e883a7f0cafc591053708633a9062ba8aba2803e3c029bf1e4d3b1b91e26cf2f56758d43077819520fe6343a0c820e9294b895f3a4750e4e1cca07736f87422908beaf6a94471094f8a4c05c0e3e5165305b989521fc2bac53a4c1f2bfc28a6b42df221f714283c92943ff274826a94908dcd75411839431b14ff7bb93e9491b7a0e8f16a44bc704b3ad06796bf4863dcfc3784a8807a812e067917441b262690b6fc8645d68b346a618f039916d04c9b0351fad2049cd1332fb0e8da8daa3b72e1ca299a986c9e3c539d087df47187a617fad763e80dcac8e234f9c0014879bc7b23380e092a2a0061e7ccf715ca6f3c0ab14cb2f1597a101cf079ee8242f24ddeb3d7ea9b467cdeec7f3b2291df9b57b2c311e84567240630232a51d8f28e6bc4b6fdf554c45ef63f8419f7b7a4b1497e32470605b02d4cbb5ee1c9edf44eb1daf4681c93241ee8771d7318f9d64b8d751ed3fcbe6168358426bd14a8010870e2e0d27a21f3be0dc597f4c4e80bccd608006054f078fe2c7b91ff9320a5bc7fea29b39077444a0ee367fe9001e95c33fda05aaa42b9c005889e6ad70f37bdb4f6bdfdb5c05073747f3f4f4df4d63f33f1f8c54fe8803f9f8b6e914d593d2ed5786a9242eccf2b54165edbda465b9a9e5d947b4fc6813755a6255df6ecc8678f35eac73c4cac180344d155e16ebe6f86334b213a1d442d318bf997ff7b3421f7c861af51fc9040cc67dceaf111f7a46a4094c56acc5f635996ac81b2e561b26b72dfef5ce6ab208325afcc0e4bcf88b84bf99778a39b2477cacbcbfaad802f6bca3dff68f44f24f3a68dbb10c8e2853c78f0211fd7660cb9be8defcd673c56840079d7c2d8e69890dcefaddfc719adb513ae6e0e2ab0487c8b35eef8050d5da07b4573db3b870e8748bfa2e288740bfbd30b0f373236c7e8001bae4c1fc35be365e6e33f45f1a845f3f7843b568d64b666c26ac2941aaf95c6dc7e1944c4ffc5c28f6e03781fa667ae361f8622d563b07196ba09d3313ed0eb738e155a131f9d18c60567b3c5c5baed4af37fe722e5199e278ff6c04d1dba2a4e468fa9cffe92b7e438dc85045a1fac00cff0e19e62a850b690c7a982c7053f3b39b8b7067883dc55ce606684d8185babda73cd7bcc105d2307d018b7667eea2736220a03f4c5b78c4d20dbf244f91b9bf88b34023094027f8a09580416c000d70c218169222398f68e2bac58a30775243db28f58948e38504f3d41977bb1e7e8442ffa253f2688273b896237ad4a169dc0bf9c607f805ccf5d36d74a043fd58563d4d5057562c05b4d52e829c59495917735101e8ac50303b1a5f3fd984bdc5d634d4b2c31868bbb435571b23d209bc16f0a5e787c7882d26ac24fa9c9bca0ad5301dc24c02226ee3aed1d83d9b4d035a70fb01cbfa9dfc4fbf07e94c667f08a804a963e47f59ca229342163cc61d17f33d7418582e41ebc8eaf0df4d941a00e39f7843a6a30fce8d8556827db75385213099e74860911072a57a62eb6f0d4686ef68c8e3522e2ff3c6bd8b49e37b804544756512e8c1b190d341ddaee087a5872bdf3bca72dea4700d030dfc12fffea4c45698f36f23fe7833f55b204184da65370568d019403f56ba7dd8b858a519e93e73567c84d03e6a2f052e9231d87c71d662e0827f0873e2cb98f21f3d1b7a6290cf8aaacbc534d85679634a33351949a5ffd842b2dfdc70364d74ca7400263295b24d87ee77512f03e535e8ab5f6dccd75849e9358aa60a958b42dad641fcb62240dbe09d5fecefa89d47c9a3ed92d236ec7f8842b1d0cf9cd5bd4812eacdcaef6ece76626bcbf0bf884498858a75c3b40d4e5e64a9b2ead35a4732b48a9e9fd9ac4df6bc942e4e72b117f3c71e8b7024f87eabc4a51140ef8d2f13b83bd53e48a90ef52d5da6459c8905298e36894a4096df66f77bf094bf5ec0d80fd46c2aa00ad73d88fd3f22aa8cce2dad4a62baa25d2aaead62f90d7b3c73e6a8575bff4bdd089ccc8dbf05dc2f719819aa9531e24c2ecf63d550088936b8bf588f85505ab0dfbe5527c94cd565e3d68908af2ea6182c9dabae1a5b4a36c231b6e9a4def8b23c2e08d939504192407d7ec391f0576a4404b469d3801cc2e9513c60b50a80b98b4f605b61326799472de4b15887355c5b3ab225a44095ead04bedf15ccac5fd9a83c75586f5219d99b0b6d9f7d0faf52d5650aeaeb2b135b8136b4eb9d7518801f724c9c50e3b5e34078f40282cb97eae38e87860139d21286912fd5e2958052137dfde3c5c6bc3a8b4240b2c3caba5578722439bf2cecac810bca9da586166cbeec45dcab09990f104f595714bc20272f0ae500d52cc917bb41e79e32ae7a77f3a04be2758a3d27f3ba218e71c77437aeac789a4e5f5be246d7f244d2ddec094a0ff3a64eb3c684c98b7fea61a12826c5b2acec892a2d6b3718488b3a971359e726c86f9fae4058bf915f883ed0ee3f3b55ea3ee844a204b6801330da255dffb6e2128faf00c0e309096211476edfd298c6c25b7a08e64c6615a87e232896ff2f9e52fe5ffca678ef7e4cefd213d0f9a14e17ec84845227521f5e3f1855141b02856409155a50cb38c803cc5821812a5ba9373a09fbd470cf77db1df4dec2f5eafe3e7e27b8958aa3e2a4608dd032ecb0bfc7961fef0eb704b32f26a2fbb07698d0b3d3d06ce97a12c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'heb0b1ede89219e180eeb5fa51175ea0c8bc2b632f7fa37814f3086eb1b5923d400a1b5cd8d7387e6dc41fe8a3e578b4ee5a0cac9cc83898c9bd9caa5810370e7e960f5e8629679c6e82b7e658714c54481239eb65a014c593b2b8b2ba40f870e9cbccd44c9ccdcb88bb0b61da77aea8b7f8cc20f7c0b2d77410e28ecee841092d33f23458d07ba57e0384f628241027e8e0bf254159cc01ebf632bbf83a553609f5bf8642811c8ebff2a2bc41509d628362c1823da188dd775d2e3ebefa6afd51744135714dcee2c40f9a32fd46dc6a7f73e0979fada749a57c9950a903d759dc572b95a32f9d11351eff6be574d97294c1160a8b19af81aa2e2410c620ffee9456ece2589f253a54403ee66be3fb53ed482a2cf2169c60b6af9406b8a42548961fd3eb1f8f23035fecee2ff66ae29625979d90dac68a5c13e92deca13ae1132c0ad28760ff9490dce6c77ae178741f7746cc8f3dbf11ae848bc626a610f7836beabb817e2d66258fbb657ffd0335e7e3362d8585b213257988d1fed4dfc48a306dfd818d5baa3940b6516a9e829fe4d647f151c80b441fbd22838827edad983e42712085ba7deb71550cda379ff71efd8fbed8419f5dde742863d2a79f31d6ba172284bcb47a29bdada9c838482129714159b765c0dab87e4b66a9256c2c5c9bbb2508290664c99a9f41e427a099d6c81cee6f9d1d6c51b9f4b7229747bf55cc45dfbc27ae0746f4e5032938667f61dc3d41cc951b2a9a2827cbff9316bde2b3970576cfe2b05b46427ff5980dbf09dcad716af63ace3bd0361630840b8602bb91f5de851d2e829b28dc6fcfcf7db36505fbd05faaa77223cc357a8516087e62609da53381e4f00fb9b1e5ae8542d97214e74d384e7a88c2bea78778fc70ed5a7880343d09e1dc49eb899ebcaf00ddd4bc403bdf14819b7e07a31e9bca956c81fe9eb56ff2569f97c14b66052c0b8989c62b271ea8637ff32054b78b09b03527c7c491cdc991f0e6b1b654d2699920a3a2112f87630e18c22b730c7e9cf57bdff3b88f2af491c13a6dbc1471dafd0f91cab333315e99368f2fae1cb2f663d086c5b3eef97d07a39890e37549c626b9c1f88217fde8882542f1031c43bbc2175b83ca6c496ee11a5f66e7f88b8aafdb77aabf01a261fc8bee97c8ee7ebed288e4957848712c2f0ebeda725aee9697861c638a90e60302c4068e9e5863b6ce545f61c198c1584eb24bd43e80acc2c794c3ac6ef1e405a53154b0e01b7fee0115e845ca2b859d3a9fa920d58eb3add0c78527d95c23cf6ea5959e6ff78b8d78e6839ac83ae4d805c0ef573dcda08c356919ccc95b81b9e7fbc13fa3966e5c397bdc51ee0730a12157186854d59554d844a15ba30b44697e34fd2ca415352ac2943ab6feff45f8862618c3401b79a33549013e8a0fa389c462fb803d237cb015b83c1dd51d4c516a95808d94916e4feb93ea14ca61a0e436b515176c7aeaa3b20d27d1480fcabb0397336fe24c454150c5c3122fc8a8f6fd0695ed1db37211b8a94cfba384bb9adec063173e88c059de7250747cc8281f8db12d1a0d0c0fe4a90b3082314649e566fd182215c0e67d7cb046f41da247675f45a5a1f3c24c8dfbc83b2cc7e73d6d257d1396884e97f21124b2a54d6e37596b02c8ce6e1fee7213b96dd4dc7a864b8b86b6f35e0c43232160c2628842f1df6b3c49a3f32aaca4dc1480054e9632be493607ba7c8c275152998a72d46ae2dc1e7826b58e7dd18fed4cb9452db28ee505721cbcf0d8e5e753d86ce45a6c9cd24769d44fad8c1f967862146bc94b7034ea98c964a59b4afb303f53ca15730584b06ee68ec6089be4d79087833da4032ad14ece70e5be2a21b9f0c80d1545cbeebfd73ac57d5a0a5e5ee30ffac185922ed3c30534c0e3916d3aae31f818f4b8ff3665180caa4e01e42e35cce449bce9dd355994cec6d3f25ebd92b1fda2ed90de0164e76a2cf7d29de1bc946871f44140f8d6d4326314e65e835226a7aa7eb746a6304fae6d77f7c08252ad5bc096a1a47cd8ce32231cba44d36b87265798cf811c178a9c60349766776106519670fc81af91aa7aef9a6c3bc94bb0267c9a8eb47faae293159ed8f6d23377b8a8a059a86a126f9ce7179cb29faad9498ec6edcc543e5da19efb113e5219cfc688abe774c2e4277b8306509c3110b421e896a3b9200b8bbbbb48512d284d075616417223d66160a97b865f610439d1aaec723b8f3f40f28e1d844672e1daf5da77fe6fd8232d5bdfbdb30cc0f96bc7d2daf6244572ba463912b02e54e3a2cb45266c699e7a631f454a29cc6e536f0b6b6d47929b4bd421e57165551e46d9cbcf766ccfda9f8c84ff0a376b234d4f1bef72826b5006b5dec202a27f600e2fae5871af7c08264afa8f299264e91ba5b2ad7576064d203d0640a9c1d688ff1acad265b9def6f365f4286a7eb3b78a7aa15c553c1570ea385308140be3fa5c7f2cc04271df955207b49a16cddd75e8d3039fe0bb3fa7b112203abe9fd3c0cc5319b0ef330e15d5707b5facfee83e70583a5f9661c02cac1252373c9181d38b38323fb7f2f6c9f6ffdd9a587288a7f53940aef08138bda4c50dd01eff033593b21c101f705562e759ca130756d965fcabac5aca961bf4565a820f1223b66c1d0260cade71cd3ada22ec9c5f9899a310abc041253bcb93cf86fecf6f8e06231e049f95ba2cdf6481b73e58aa312cfc38a00863d623d7f7b0409108e473e4095b66e74f34332821bde417dfe15345d056acab76d472670b5fa9ae99fa5a1f226c3d50329a5d428738a48146543bbc9045ed1e07d9b4b4d427df018b059bf4951a8490e7d78c832ef251d1da849c205737c696e5f3aa957ad990008872a028897dd2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd17d7b80688da5e948cf28741887dcf24064937aa5ad3feba8442fa119e52e95731ea4c8763a4340b37d76cc6965d4940f705377d16f056e6dede3f425284913bb37b159c844811ff30a70d62eaad097f9cf2a4d845b439a6ed40dba67d096318e6a46c3344f7df2e4e5bcf1c94e538a7d5e8ec69c3d28d53dd085d9ccf282c2d33ae0ba17a4e049f4252b5e2ac0efed906125fc233a8fb8da410d6335be7330b2d66ba6b4eca489f983e640c16dd57d3f4a7d9a8aed156bac82da14921bb69f8174e13ed377b2f3fd514e3c711d440198e2da380fb45a151d66e3fdff07fbba32016594417ed704101b511f12cd523a741898345c7334605ce2d0aff6664ff3f73d56df2bfebec578e5afe55641cc3502161f6b063059fadaac897e6045c4d90849ec2f7b6aef23c85107c9dfa7ef5ae05156511f34e142a083c21601e15cfe9047e663ff031885fbab3f652e6f8d1223138f0ac763c33cce7a00b1e9a334b4fdaeeed076ac9e0dbed7d91c51ce329576b9604af6979441d599ad9eb8967e4546ad90055023af30c449b4c8ca10248310d8c79092f53ea12bb3750b2732184c41156a147ac4427b890b1441bbe30dfa7603bb684496279c3fa7acdbd18877ace660c4a6d3241ac3836db76306711da5995d78c51547339819d37a461692b21205684f0b1d49f621d3b2c8281d380b53691b314687cb699501d8057948bd8a0630f0ad6a7901c463456b0946837ac966d6a5fde995e035725ba0c90727c1d88d39fded7fc385cbce9c79f6c1fc2b8d4320a6c95ea89133f87250e7a0fbccd0db9d8c06d59d8217353ce637a5c77ad73d17f26aaadc2cafdebf9dd1149d53f9738c98dc23e03aa40b4580b7256ae327263683d8f5806d72e47adcb8bff6fd33ea4e8594957dbcb816fc9f7281e1cb4fafd60ef1acd357a1c32c2d0ebca5dacb580ba17e75b070e45aa3c2bf4255b7280e8d37273882ab163f748f2d29e1ec6cd1e79cfa241f7f574a86b8b0b46d697541b4f928c804d501e7c69c5ab0d5b269faafb086f132d0b0e8e5a328701c7a3d509bb104aed0ee75b86b807f02ea36e9961af77990534ee51dcb593385f6812a0fb56635a40643fa2afa6fdec05840a93cb2e8f70433cecb1c7b63d35a7951edd782d9c873245fe318862009c8212edbbc12db6e337f063c352799a065f9dba803e94a72120570779a38ffee0b9e90324298b23233c6be3255d0c2af99fdc9e3b0455743cc3dc8824a7614723115f7c3059c4f60410fcec409e38e89c4f743f14322a9532b4aa30d249953f16b0c212d78990164db6c38ed476ff8cc5023b8d4fe12ff0e0d40e0b9d543631f1c45d776016ba546e27fcaa4b8d7ad81ccb7f1911c31835bcf0933be7244adeabda6be4cd2b4e9c5749231299dbdd28fd6353f7e25a4568c8c9f4bc2828403050f5cf16185f51707437ce0d65171cc50ef60a609b5556e3cf0c25bd6d67819657c9c40e61b51a141db0a80a95a2a493009c68e2bb53f01a22d009365ac543c642327a513b61db75bfc5a182cbbf4ef26b8b7a701c5ea1f633b89209b795727d4f7128d96c1e141d311b81a464d5d1d4dc729d33a5b7c481c38397b51583e43fe01e82192c86b3967a62b6bffb9127df093c603a52c6aabb163c3938af9ca90a25c65fe2cdd236ff47b7225e42dbef0583de647865046f9f2699a6185db12b4c2f7a0aaae578cb09fa35fd596c667e65fbf3a0a0a439383d9c454bd0f559fb4dfc23ede327be66619765c9b32078c2ddfe59fbb3e1c1604f56a071c7682fee3d39848426a3d8d5fa63d234a4b7223aa011fba07d9733cc80070ed3e417c4695494f027f88d3a50dbe82d9bd25c854230faeb7f91038e0aaa1e606cad03de10a5d22bdc1ebfcfccb1d68628a57ce536516562a6aa31ed5b8e0de9b956c033adc79807dde3298b8d75d1248d8dbea51c75d3c7fa69031539f00fa4ff82dd1bb3c89ac2f63b19b298d355df961b79b76bccdeb6d24159a8b6b3edf16593810bcde903590c9660ecd728f9ad81e52ccbaddeb7658b742d499e1bba3ad2f71c3ff9ff7af805f09f43c15aad79b135ab90a071de41a6af4f70948f6669bef333fe446b6bc768c9f6539ebf6efce966f7b8fc059f7a560362dc73fe8ad329b7c360a567304a4b5414cc7799bcd5a1a2d26cc86a82d34b76c980f7a8407d076e0609fab5d08dc3b354942e1660f3ff74d6a031dc65f16e6f639c87010c32e5a0e12920f2cc243448b67544b03f63b22a338ee85ca2828ee812007186e4006fe89c5c089564baf0b67adf0b82fb459c90edecec349c20a8d0a540a052a7221ce289f3288c2475309ab449e4d4b503708b2fb14d6557beae6338f3aa387022f0c23ab467d0ebce6ca37d32ce47fad19fa28d72171a8c011b914dc263c9a1afff58061d346fc482c36d47f2eac852063b97b4bd60664d50e715026941bc6ce60ebb735f7145f96e9bc45bc1c3fc185c82eaf7abf008f580e3dd300357b7460316264d7accc4a1295cfbbf32b8ae9d64df30bb5e98dd07650f3a174b114785b5db30c5b54c2966f7aeaa587cca25b86fa4ef07086f6311291b0101e7290a98ba5324a44867f88f0789a2a96d8b143a90acaa568cffdc6d9986106394bd8cce310d2fb684e82a7bee9f93cd2afc195e2feb0328956544a6787c619951ca8ca669b1fb92761243ea4f415fcdd6e0739c4563ce64aac592a581c7a65847e6923779742e6288a8bc6f96487bca566a0b8c2a7130f2f250615b52501bd63050f13cf0d456a79fa0c26962034c2e53c6cb760dad5a67418ea930f05dcdcbda0fbf9f1e4c211619db283811136debd721550c9373c0c0ebf5c7ad2b666332d954dc1637f795d70cb6c64b12f91e5ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hba551f6595a5b44544f65e53ddaa130229fd9f7a476830f9e54b3b51dec595251e09682e9d7c9a2452568a8b55aeddef813d8a5eb7f3cbdd2a5be2112eaca79d7c489b711222aeb5cbfbccb3a4c90c32bda025f1fc5f8092ef31757822fc0bc83a45cbdffd73449cb8dddb534a617c84842275bec359147a265b67ce913459fd66181b7493b247722a72aec21c4728eb592f30ebd7abee8775436607a42be64f672ae481689dd5cad36fb92e9b6d5171805cf33c221064f80c2efa42201e1e466e7f122b0b790aba96cfaf1277e39d46b74a16a389d9b7d5001ec07700a667afd00e7e2c4b5f5cb66731ecc4ee2e71e8c83a1cb02f3bb795685ee874c266ba114683c980d87709f7dafcf082729520d82799a874991c9f6431c3d582f954229b6c2f7e6dd00db19a5f11e54ee8884ca1f9c29c35dc3c8096e807f483e429a916fd64fb91d29694147550ee523437c5a2432e4b1edffcd381bf508e11fa69022d3d446d829b3121f6e27085c14066c4950bd9c5492940a584f66565924b8300d466304823e74b87c31b01c566d5cddf0fe118f41f0b10aca4c8afb4b8d112aa695a1026d4fb43fc592fcc4f0a88ac4b293b4c4bcb4b33fc692cb7c06ffa5a56517a16d00834bc570594ae8c066ea2173123d6964bc582cdccebd57bf7dfc4f3fde13d623290025d979aec3410f3c3575969ea662b21eaaffdc86231a4cf56d931e6c71e0a6409c3091eaf85041e0f2f6a53c804ac41e30a10086ddc66c54150cf1b0c114e34348b94ecffe85b41bf7cb9c6aea1b5d0fb67f99d3309dfed910c6d3127da69f8e7bb1251d55505e2a6531df9994d36d3d1bc51141eaf0e6e0ce8edaae77c6373ca99499a87a0556756cae7ed9d9bfd0b85f6ed17a89f1c469377c030f48b8f8fe8150d7423d843cf59c6b997fadd98608d681071e5e31536750f9e262bb4b23cbad7eb6b22cb881ce8d3beb21c826a54067b2a8c09cd0dbd11693f79f2b3835510c1be3231e19d8fcab8272850c0fff5180f08c3629b19f8b57442b7f37be6621eff90b0f22ea1f03264249b65850f096e81a46a6355b2410a4dee3a324e75df942a68407cd824bad8d86a6cddf68204b896fc330df51bb32cac64e14216b1efaa17f8480344e7bf0b4ea8eb00e223e17149961bcb599da786dc3c7467a010c296a228b1b1b3746a855daaafbda5f9501d00fb7ba3b88eb175b676eb1278c7f7b39da1fec3e448ea07ac4009630de730d1490bcb56d8727ebbad39ea990777c9f19a1f0a8536b3776d5b815e6e856377eafd07ec49a84eb5e9e4952665862385ee101bc0144380b54055e51d5a7d61e62344dab3ad7c9aee878c27d7d730b01d4428e96fb380696dab26329cdea81f9b6272dd1438e748f2718be276a547904fc49ad832a08018a113f0e2e302f9ed7c9ca3a6452c91f3e2dfc5cd9e26a7aa87cabeff7e9283d06693f9d3313cf5957b460e9c155c6bd1c12fc56d850f9cca612c4f8394b500db73ddae7b3d58ace913f22f0890f3a555b1816bd87e0e7922bc4efa66a4ac4a935afd1eecdbeb7e8258ea4d42fa8b6eef0ea0ba6cb916c10f5e6ba8a1f20b84e9107776f72071ee579c6ca2819b172ae46c1b40b33774cece3659aaa5129b7dda29b828edb0b07e38572cfedf14cb92f449696bebc4fabc9028f91ee43062371005cc04935af7283e2cd3ecc941c7f3d1a49d92686ad08c531c4c090d39dc061dc012b997cd40cc50384ae8ca7e3e73ca0f0ab73a2e0b5fc4f35813ed010abd5391ec084bd50adbcf7d478dceb3dfcfab247320eec034f9e98778cd96044bc42b1b05e97a9eb21de01aa1530665e0ef57d00a4cee8052b0298257d841556e56ed1ef93508182ab478ced95a03c1f56a20bbdfae4e9173cb15a25e3a1021643918e989e9db5d7e411db4c4921cfb79db968e7a4828e05c9155c604c7bd4493d200dbe197eb1184a853ece627f3f9ec992d675fc9a61e9907e70ce1330487751a9147b5bda7c7b107294e35bdaf51d02b13bbce3598cfbdd4aad04bea74af261c6d929130b61f5ff2e9ba85e9d6e03fe26833725f9ffba4ef0bc27468fcffdb9b32e8e6fea33addd7f7a2c3a7e4e0aa0b9d8ee8071fb7469aba342f6febcadffccd781cdc2682d3a199b065fdedd0f4eab89cc29934746c76ef6cb4d5a98bb9d130e8c39ab83f794477e51a047af82ddf4d5e6061171dc3028ed92dbb29ff182a593cef58137975ff4e63b058ce443b4ccb511042acb7cdf073d9d3d3dd50dc749f72a70c41c8d52ab4ac9595b42b8676e816be65069351b3f123dd061bb744ce5f79dd237e35dcef24d0906dd4f23977fa8aebcfe194009bd79ccd029c2263d3908e2e684fc8132e0fa42620e98e511f60688efa470dc23b28b80adc49fba351aea12f417663e52d320aba25d7bbe15d7b660e963daf09bfaea16a2f5e343a899743a7e817b5e29454ef16ee2da470210b4e17b9871f4df69e29541ba89fdff67c0000a2239e4139fa9745ca1514477cb230465ee57a21706e832f5955c00410a613feef07dafdb195828b1c505d64f1305d15b416201985701279679042179c223dc45de07cfc6dac66409d69a98178c50f9c5bdd724c87ef7d3778abed21cc193bde8885643db0c15fd5d5b2aacaae0264af5f66fcfe1afb70de8489a4a6b51a394a71d60a7bc1085b8e691fdf0ddb5cac693d47ed270ed53bd01c717f0d24a86eb4bf8a43cfb586cca204024e039eb4a12119c45fec3a0a40190f1b4e33e00a87a0bc2a84933b07dcfb7f7aca694d8b53ec76a98cb9fa4708659bbd66728440f4bb7fc40167c0510c302727ca74773f51a5c123b0d5d615d80f46ff665ef814456a43f836fa4aeb33b1e224109dfa5c4a9c06a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he8b03270f5fea625457cca23644ef9e975f9eb29d678d3546528f67f3dacfedb7fff9aa4987b00352580cd0a8d6eaae98cacc6d8d3eac7d10f13f910efbb04f8ee7f19ec4fa1eeaf7534dfd82054b47bb2bdccf8ee8658b2ea1335f7798d51df8de8e54dd6f263cfe6e366895ecfe77b138ba53e47abd47869aff66c2c6b145e4d7981309c10dbb75eb753d05c8f0ce18789f6710b9ab55ae909912a2a95f2919535fab09d482363352a9dfff4ea05c42a83e89f745c992b23dd0654cc71d5f6795f0c39ffe2e3c9f93c23d13922ac7f648749f810316f80caae36090b26744d97d943281dcba549aef2bbf440d21de639048f5c2bb2242bb407542b8d4ff20ab6e1b581a85e7af49d87ebf7271269dc8b910316747585ed1c3b8a2bc36930be9582addeaea14f9f7175e122d1bf36e7f40f1681217b2abd9522f30788957e28b32472075e9cb3419bed4d523ee0fefc881db8a3083ccf3667e6a54d14d2b38e0aab3246d91122e1892789178f91f9ba2714625d1d38676d1ed2a3e9c6520c6752b15b34498c0096fd295a7db6b28d770f60554d17026abb673d796f257f31a5193820767ad1aa2d0f276d987de2b556b53f32358e958635d43b6bd5341477d8d8d1064b1eed02d37cbdbbfdfa92136f97e257e902dedc2f3eec40845b39ce75c05fe0e503ae5565bbd4222892f681a497ffe9e2cb9a65d3a36f24e01bc888bec0b4d705bfedc3a2d7b25030b469438ecc4b3fa3262c8abc85041f796f3cd12a87764271cc60cc3517ec9f3062d3a1aa92b0acbb3c5c1f0445a9bb342f4cf1c8f4b7bd0df715db480aa92d1fe6df0f115ad9c4ea037afbe26a80eacea5339d2dc101b6d01e44a183f69b5a3e83825a33431521c49a5b13f7c88ee1e98fbfc6f1e6675f962ee579186a87f320d70627264e79b61e362966827d657442ebf7fb49c75dc36aaa94294d99e1bd0264b2e75f56996c1d9155cf70217338a8779c7d81e91c167399f8df0026e7b18adce86e02cf58acc05bd4ba380d040b1d8aa1e534be4459b3001a8ddea330f3c927e00135988623f6b64df89c60886932635ac61e2108950d2e46bbb909168675abcd29524d610750e574e428a78380542a33e23a86d6d7a5013f1520b92633f1a1d573308b143d8134e439dc8001cd3539109534cff9e4281fa5e15ebf61c9d6f22cadaf4bc47662bba18f9a38c958ddb44488ad365ca4877e0a23eb57ae0df688df2e8d2498965d9a7c9b86493e9bc2c65318bc9e279fe8666f379895d25e00b88e46171b28b833c77359efd7d525d31215cf04891013cb8d837bc3d7ee931d15d2b567893fb22b88197612560f3073bd251e6690b92a91c6ff144aab10d298abf36451041e657b542cddca42326127692b328a4abc28c12625ce1cc1f6eaf53e66ce99b5b05b591b44136696d19270b0dae811e3937e9d881d838fc27002b2e291ec0abf57fdeb579cb28a1204b5163ce0f15a9666caffa7d96f36447e24391480af999c37030bf8bd3177d054d7bfc4c2f83cde9443c9f3d813d1538a090e6bd47860ce3a458d401a22c1442c60ced9e1218dd0f4dcc602a061b99cb31038ca10f2ecd7a13612afdefc6aa98b8fdb722da53675c778f4c29dd2f2b886e0adea8e745dd10d2e1445b1d6c53c49ecbea9a799539817a65f1249f40278ac16e895b9a87009b0faac15cf82c823c2c97a1144fe94376fde65ffc54dd51878936520c7b9ea98bac51ecb40654558967dae15da02468255a3c26b9f1dc95645490bb42b950ad0ce6901fa249ae7cb152f5bcfe4ead2776595cf1c9f0282c582c4f6cb087e647ad223ef42371e370578e98309090a12e89f43504a1b65e4ebdb603b6608f509c98eb66690f19ee57d1d81460a4f595c241e77b7306598dd0d31b6ce67a95506fb7de73c80409b23378719929becca638ba39c9459472c120dce63bff3c9a5e7e509d1fb772f6f02991e16a75ccca3ac4a0d74ac1a92cf0d6790a8c8baf188a54de0902b81c0b64ead6aeb5bb68678dbcce0afeabac11f1c600cd9a41f1304cbfca29373bfb0347b089c42a4dafed4f06d1ece873d1e798633977db77ea2269d278c4d53b8d5bc182f16c6ecd0a860055a49f51c1150fc5742019d876f535ecec522244973013095a1abdc14c6ad3a98afa4e6ce83f03a6099667ef415a6db922d9663519c30f59d608c1d3ec89c1f32399e00cf1e06d4a66b14aacd990698d39ad708bf0e0f6a9509ee9a1c69668717498e78b3b42bde1bddf6715622058ae534d5c1989e399af4fdb0d90dc81599e41168b916c549150463973aba5cf0db7d1d987a269b0907d9fce089187e3547de599bb9998311ce557e39bab1fe633b07dd732b134ea81060f0a43d0748c51a8ccc243b3c2e119db0279aa63cab42dba229b9ac34b6f28ba75cb8e27fa02f0d87e61417789e8869d8bde9adccc83c943e16f5de3a3178f7a2f3aacbea6a4df0dc21e2c75e4b8c9d63e6ea8a1849c5e9b610a43d36443a6c4da7ec39627dc2cc50dd753e9f85cfed47de00e7328d45d617879b16b0075e280e92df91493c8ad93bd2abf9054e2ded458bdb0ae82d0b4d208fcef64295aa87adace5ed3499cf1e851f95e7b8283ca02f7e33c50f27bdd432f8f4cfb094d3b841c8113cfe70a7b4f38c03f82db7cbd67bbac40ca9ad90a230be8f480aab96a7c699b011df6505c8ef52488fac0b14d757ea62b58dcd6fa1d1bf6cd732e87dcd09f13e29d8c62b00d63523ece8a75824e1522e78439ade9dcad213bc1faf2d3d9831a0fae832a6d3122b0c9982628452dd63f5440be0f52253661268a12104881e198522b6163c2aaafde3fdfbabaab6bbfd7cae7d1b934f3c487e9cc03bafc680b473a60c1b484a27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf426b7ed59c53347c118c6edb10c15c495e00c79f12d2b659bd3c674aeab793ac481e75b2401fe13ba2bd42e3283a732b884bb3001df5e16902982ab89fd77b0edab687fdc3b9c665dea34f6c6935e154a31fc8418123f7b7896159ce248bc64da7ea7d2565b45b474d1eb50572f70d9aecc3252897614c272f5c83dac9fcdbb629ae8ae7ac8c693c70f2f477d0db9faf3f05fa65b126ec6f191e1b5b9e7eb77a0275ca67b4e134850a004c0e084cdc07e695efc9648fea8df408bee7b160bc012c574b4b48ad13e6ffbada97d525c6d21e8fd966fde08f29aed5a7163fad53af1a2f45fde9e7fbfd0363ebc2df43819c6271fac8050182bd2bbee27c9868cc59e522ca56384d5b2e391df359e0d6cf1be847b6e3d8d35acb13af70e18d2ab47688e7f8d1e58df635a9b4c41d3ad9f9d735dcc5632285d6070ae6f876d6f2f3d14d73cef9755ca9dc33912d336012444b166901e76a11757f0a51ab2578c5bd678d8a464126a122bd1e9700f8c1850fb73b8f54c3c26997e19a8b0cc7affc020d930f4debc91ac66e299f4e82a9b87c3e732cf84aa70803bf831f49c243d491a9e0ae3800c47033db9c8743361cd5526007dbb012f7fb090e3de5d64144f9b673dea5f2384d668939bc3ca6ea1a3e21552bc96823b07d5a554a914885efda16c0dd3b78e3eaa97c638fb3dd1c3a92ada9e6c5d2859c16469daa3f3303af09063f0fa1726d23ba57d61932931133b7a4c1ec8b951ce49db06eaa8f7f15c3619300aededc94bf4a097576f5ccbf0dc3fe7a4433baaad45e228e8fe5c76850629a87b14a21e07730138e06f2d51468e20f6fa2384b10ccbf1f968c03c165cface80771bdefc2f65ce51e9d5dc029a2defb7ccb0cd237db77806757ad8526286a478d3a2afb174e51ead731593be56071c380dcf60bac4c039899fad3d9f956d064ad7d183ae9b38aebe2a57c81934eaee6bfc0438162b1257aa043a3fcbef6c92ad9381821c2e9981d8ab5caa9025f6c298bba196e21a9068d7d45a892532409f538f9032d1180f6811e5eb29143bc870d06be6c60092c7cc7b3945d9263d59d761a459d095de1b1dc25b8f43765de11646cf492ec7cb786ff3228d067fd7997a494cbec51ef0db1410d4db0dbd4a96ea9c4dad78f08b14bf6f3dd5f8e6031ecbf4c468c9d90a24a2fd30adeb27afa558dfa16f2a528702dd7d555bcd835e4e1badcf8f69c99c51da40c80f8ddc426446f2a1fde7ad96ce9189795ab65ee50fbbc6a382903bdd063d4fbab331506a5afe96786fc64a7a2d4ddf7ced2941807d3abe8219a4c4dca6cae1c6ddfc22822769e47754df1207c02fadad221ed42a418caff610552964e6a99f622aded6915508d44ff4eeb3878039f862d46021bcd2539be19646191d1d86e66cb466c9e9656d41d341cd8989c38cc2a7ab8f6768705e5844f8beae78daab7da1e5e22c7eb6fa435c9f43827af4c829ce9e6718b71c414e6784d3306d57efe350ede1ab8416341dd3f80e5c18ab24c30e5574b4521f576468e03de2af4dba64c0a3c7dd20d5b41c8ba869f910092092498f3503c6aea58e99bc25d9d3c1fafa386be3131ac9ca815ee0d27a551a3ea0781981dfb4b19234e1ef43bdab1ed51ad598c259c8569c5e091be6a667873063328666ec4996633a33e756aa25f1d837b433c7591b9ca72e069a8ad4f27e80a0ef3ea25551e6c83a6df35fb08708054592209ba95a8753f3c4e5545cbfc6328bc7159d5cb049de4d78f0081abf8a5634f586b5e7d68636298abcedc5a1a1c65cd8c963f1189d8d593c5090c80cbe3e62db333e28a017714d35a04adb3b285cefac1c58f9cb64e35ff04f97267838375e9d81eb4c2780aa1c3a78316c5ec05d7998524d35e83da85fd271f0471de451979cd856c79461a58e9975b36f906a2cf4f6d995433fcaed65c34007e7b3a4bb3ece1dc8c48defc35b6d2df3ee83124a2cba054569b44a3d528fdc2d27d19d20cd68e12bedd2d6241cde678274c13f5ecced765f2ce1e03afc8d0365c27e3afdebc6ad9eff460c8ee4a8d33c3ecfe5ab1704d3a46eada5a1de695926e612bca1f5d156aeeed66d23a2dbff7dc8f6bd62d08207745978c561d6025de4c20b0115306d9a3d670754dfe4b0678e20c41df943d3e16ea4ebd942a39166cf67f6a06b274d41a96c81c8a27e723f3a9dc8469e5c682fb8a85ab902915480fcda9eeff347e58912d014fedac7677a925d137baeef35296f9a5ad0cf299522001268010cf130895e93f8c806529417ebac96918328ab02f0062661f7d464386d82768b197ab78815b52cbd82cca230d3836304dc02ece89950b34531c042e3ae343a9f95b0afeda998c070c9da04a2474ef4fdecf5d58551047e0134e88148241b9464165dbc9bdb4a73906a99362dbf7cea8cb6435b9824c8897e1640a234bc6e316499d3b865ae9d109517a9322b7de2197820d95043acb491fcec7467e5ea97667b7e6faeab8c495d2c2c4f2f44b3e4cc874d8595b990344ca360dc510703b764b3072fed7970f7593641d621d2fe5da41225a03979113c3e30b8d5c5dafd54bb09ac8905bcffdeac91ccd636c9777f7b34c42fc6c100756712da65f78c6f3d2b27120015662a42d3b0a978fe5a05f625f280be4011c558151de99fc5ccde277e50526911c8eb0b718b225efc82c8bc7d05cd05d93c90810616d1cf9d04bcfd9b04e2a1b858f71043c69fe0d74cc07f047504e12181c6ae3080b4acae328cc220e387967f47930ec7adf5eee8dd181f468074777d4b83c25783880172410d3db0c3e498e880daa9edc8fb172a4d727d651ae1e0df8d76cdd6a05badab9ba882b944e5628caada077370aded9b989b267116de181ebc1e86e54aa494;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1935a83277804a779770ca31b58cfae05f4131f4c186faa43b7cd11a997015e722a52a466b78f7a6211c904e57c3576d918a188ecd24f18a0a60a7a36eef30def3e63dd9acd13e5a3cffbeb1749a0e1092f5ee547b990e4af028c61ce451e59eb8b02cf48c8c819bdb38a2e9c03574ad471743a0c7c154b6cbd23a9da14bb0cdd4ad1ab8ea157e118e9a294931caf6383c69ce4faa1a30953eca6c5c77d4782670d5247bd46ff6bc6f840a79104c6fd35285ba01292df1c31cf7c93677c03dff18a0c4e7179e4c8b1f7d5fde2fd963c7d7d886c21cb3684eafffcec9585a179a2d2c7d0a6ed01b5f3107ac6d9c7c258b70f3d55ddbe6959b4fb3b0e72f78c68c362856f7c2727c3fe38755769033c5dc4618b0790c0999f7caa57ed1652049afd4fdafebc5457273c23c9cab6c9632b7774a80e5d6d7bd54bbd50cf97d7acbf5d06533569344c20be4dad9eb54efefae1e1f204ad6a785a01e9e44cb4c58aa0c42a309b2ca293e6271a1bbd24d6fba7bb11b16929b6778961250b9a6cb7a2560f8d106331bdb333cca6da6bbca9deb86e163408fe70afd2ad3a0f1c160f48a72d86c2efa043d3d9fc996de778ed05c08773d28e7ab390141911e30ed21155d4fbc5ac7d6b9657f05900d1b2e3d3445e038ca9b8636c27779e149fcb2a73b95d0f8967042a4f0d0f4ce7905ab98d48fc641252b61a6d70f791370c3d45ed87df8d898ef03fa9dad3c0bb96c083f831ead33444322c72e42829cac61160cd52c5b22edeeeca669b3143e718bda420a6a4f649f49bf2958a5205ceb1bfebb539cdd6847b8d88b4ccf204fbb4ddba4eaaadb5c2ffb676e6f5737e7bd9446ad3f8e8013a1ce1e83efa6bf77d47100a2af71bfaade501647baac2d1e562991dc595cb5f42e5d61819663c009f47c77aea4ef47b3c5dfb4d590a52f230c129db7be2dc2ac6b87f54559d708d2ff270168ae8317946fae178312b71ed37206ea29a865e3075a50309951701e6bf785ba61bf1f8feb05af50cfc1f156708003f318184965520ad49021d7ee1e58e2bef2d39c7a8a7e8f6003984806b647016b58261a1eb1eae35798a295e1350ee9faebd2498fd4997ab34633e033c12d7838051f878db86bc79a16920299df79c8d7d0b8d113e02bac1f6b388dfce42a01066aa2e563712102d01d4eb7df2d591b6a68466a4027fcdfe8c43e142388ceb8cd7688582d51ee51aa3eff31dddb9091b074f432c702e4ba097379c3f2ebc55e014f4bed8fe3050dc49de25f68da567f7e256bb917d1a100aded4609e2033f93407df2f01c1e8df031c7ac8c49f9c6d763f5861e3e70bdd5d8ed642167fc38a2ccca14892cb0d761a34add20a3ea4b03a4e9c7ac634e7de650b8fc0cdf01254b8e5d3c36fd47ffe6b094b80693a624edd1b2f5822dd523088024b8301112cb38e292083eb0e2d69b25085a0fbb376458cc3ca25a0461c9a3bf8158c1833bb8ca6d0a8e01edb9d45797a5096d90e95af64f82a46bde8e30421ba123fdb47a33f6e5f96302789bed9bbc3924cc99ff854c1f603f3b3bce4dccc57a5a127769b69ea15c872c2982bc815d97e13fe9943e1c06179462162a1d7af27db514978de051b7f1b55924712537afc7ec732b15b8b541011b0986d483ab657281cd76d3778ff1c54ccfc32f6469bf5da3886d56792e455559b12b28c8b2bd665d760bea86d86ee4e0e1e1f1c4698e6a55b8455edf4cf2d4e7aaa8deb210decccba46e3542f6bb431465cd5ef78d95bc70b261c3717037d9cad299c0ff090874bccd1a986cc12f83139ca2b6e1823673a767b0afbfaa1e01a1f07a3b6cb227bfb903d6c18aa2b6b3c30cfa92cf850312158f610e937d10c7a956cb9e78d5293a07149d0ba1c7fc671e626dd6824318ea873173464809c4dc1a5dba539c6bb6442f95a92cace3b05b1b24618373c8c172ad47e290e53079f8a833369fe6e445618515c5d1d10593569654bd371c4ffc298f1c412535b89007cd2b40e83ec072f4c01db6be442171965be42f2403a6e5a0182d6f11358cff48b53f071b64fbb42763ba6bdf7d8ced3e72e60bd34761846b2bf25b9d08f39ea5641369cb09f209e47a4ea627e97f93db7c65f656cd62a1ca0a4b0c294548fad73413e06d6dcc7e7a3097c4b10fc18d3f7dacfb02213dfb000647cf0d01ace2fcda04853b85699bce9af03fdb66d88d0a350958bda6579ac3d79e6ef09d19446aa92c4d149b20568d97c38f5c013c7ef6586fde9a338f84a9c442114736de0e4d7bcf01f091b83ce19174a230ad30d34b463b47094487612b8e12236e1321bfea9ac2e2c4cf4e4d9ef740d9baee0ced8b7739a204238628e1d13582a5bc4d9eb2eaa27fc57e135dbca5b943594facbb2ebd508d9ca17fe14f2803f2a9ffa2e78ce9dcbdd5494b63e2af6635a104fb758145b4612ed9e17032a8b2ccba159561fe4f89e4d75701943691b3b7e5a5a617324ef5793c2f120e2434149cc43d5ad50ae2a53835a9c2c1242c96f2e617b76a0206d60bb7e1892d4e438b96cabcbf871318394b49996dab3e9e8c6ffd392a118225c73d2dce6c25d17ada027f48a1da34f59be6e7d523f650592a32516281197c6eb9615715f156d138b0e49557a2310e29415136e51a608dfa4c6e9bc38d15da572c42e92f503e8bd46ee4ebe8c4aab3c8d9b3234ccf8ed6dc1bb907a4a9a4a41ee6d8bc3545043c720692119c08b5511d8144aa6205a8e7635daaec8b68080022c6c4c523eb3aad8d657d730c101f42a367c14c457c65dedefda9ea6148cd77f688cc1ad8e61cadb371388425a8495a88741d6ce8b0f6c3e0003e2c83123e43b5432b477348e870064d1ae18c23996e5156bf73f7a19ea530120de9c790d5a850c0184a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hadc9615115a021631413d57a4b52b0c584515f41d80671679606a60d9428607f1ca3ade55b16280816ff3f5db0c115155f6c4041dea522a5bdcc938cfbc7c541b3abeafd6d3dd4d0c055c0fbff557bfe8f32e2b3a754eb46783b273bdc5f0ada76d6d3b47fa4a19b7296f34063847833489357bd2bb768b832b0472a5539a77b63d44f2ba4331db19fac1e7531cf3896ef100257b75e3acb3df2bb96be72ccf8b1b350cfe7c85e861a568f06d657961d276eded77cab49c3a72cec1feb1891292f3c2492c1c530d809e4021b9f62590fdc22c8e975cb7a8862590b0c27eaa805da2d705bcf4aff1942165e802d755aef85efbbac4f28cea572bdabaab131e1a0b89900da0a9602d0579e4d273de29bb58c6cdf3f5f17fcb630a96abc58b05a9650f3b523a1439242ec55de8a3d5e1ead38aa1514af04ef3deeb1502f4eabf011d2228b55b2d620688ef58f18256926565bd27136483d9a601e0bf9836e674fe1c42d187d975a7ca83048b3266152c8709119aaf62c4d5d8960b68046ba41618ac16b173ea8bbffe01a8c798d7e4e89af27ff2102149e8f851628b93a97321393697db21b8905374e3c40ff4df094dfc2ddf4595113bfce5eb327b95ea622aba7ba6a43a91240677dbf59bb1f1e98823a2818e21f82a3143f830c73a63e06b18c2dc180f3f44b928fb1b3492303b82ebb8fc0e0be961aefc43f2805a372790ac48ad698ad7a205c03b33f67d2b442a930d04aac601796a246361130a7b4c1afe9e0300652040c226b57f48f2302d65212fd9fd2f9e8b978ae8f777f308bf1a2c8039bae89b6ef86419744ec7925506a2748381c671c3e5faaf47fa4f8e92b063019e94775f6a2812cc3e96b96fc220d9f202686f67450142c225082f1e4c57be7ac6991150fb23b7949e055a0828febda5353c4c2f27e9147a46abb29de6939d56a4f6fd1a0ff190ba360d55ac66710db31f5645f6896c67eed4f791251733abb09619a511f19f16eb833c70b43457eb8f45b4e88dd4f06fad3535ee2798dfe1a7ccf119199c6933eec0b67fdb779df2108abd7760e0f35b75dbb1f5f1d08654457d30c17a6e68bdd9e83fbb06c45f78fad1390c483d7c056fb48b1ee731328c9c6e55a1fb74f5465012c64d6dc31d1b2e793d425a9b4b724b7f6474e76ebf58d4001677855099bd3ed1c13031e7f834ecfe145ed25a994b418ceff0685cf04d5a56a9c8a7bb7238ca70023e701ad1c8ec14114caf84a94691d506a628b9110cdbc721cd7d28ba41cc1595e2d4929aff5f77af3d06723589f41629aaea744a152bb3090f52ef6afebd9fb5e2fb0075cbcf8fb0e35f07f180e6a2cfa03e045d9d1b68130954ec3af92ac1d72d165b429b7400afb3a1f32f2f03457c4334f855c6dad93c5585def557775dfbc17d01221124e8563e4a68500afce746ac135554e267096871f78c40cb236fab5b038853bd4a222e57191980995463f0f53dd4a8c9bb73cf62a78c990a76271a1e741f027020796e5b65ec146d87296b84688bbde1825f46357a8f1daf8c3904063789c2778969bd81ee323101fbc1039415382d4845647fcd51c9a9c5ebccd23603a7385aaae931b7090e8a588fc334d584c6d6d93e44730a90f21304bb3f30b34f572d2720ee7a101eeda32054085ea0039fb9970a8e7eff3342fe51569119e2d6f4234af500df160d1acb57d2f55d1da6e9eb1355fc1cd7a3b54b2868abef846798c38f23b99b12950164630922d8b4f45172b26547a1152db8d1327b71edf2ae1cd7c68d32f9cd970f5aff308acf96026285e22ef8d53dafac71953275eae6eca19ab17fe7ceafc16a223e8999776192b3e40ec7c892557ef0ce503052b00530827e1214ce5a51caa307a846ffef99a1d98b76289c2410f3c7062ac801d50a5f8d69a430098e9472f05dd2ea33e3435c25ed49a1128db82a08570d2f51a3acb6a21a7ce034b979e4ab0a737eb05c43019aca94c576558e99dc6b2d4034e94f3a2d81e160d12b186d8db92e2f0150fbdc6e48fd677799a6f70505697d1bfc637056c9d42cce779f4e9234b291c8997dfbaf32f26c4dd76adc7a810f401310f3e7d32cc0da071c3d0d167896f72c0c41967fbe0cb0ef450a314b3d736763b8bb11c8ffef9a18c5fbb6056be21b9c8f93c10051ee898e0b1caa64a31267d308298192189c5d368ddeb2c472fef58f8a421733c2a4921633f8002acd9dc54d972cf1051fea2287b0f4e735d55ce1c2c9a64dac53e5b26f455b6891272545ceb54b9564a13290e71cd2e48efddb0a2e4ee942d85532094a6d10bcdb54adeae4b48bba16c0c2343839de8cc468d0dfa0756edbd744747ff4b130def97f1b8b15c4dca7de975b0a88c34e309995dce128dcc2525dcb1b414a7e0103570eb449fe6089ab8deb8a78b895bfe7b959b97fa0c6a437208a5c17d7a8aad8e906a053c7ae0754292240ca36c146b9a032d0db32b3920e3d40ed5fb18bbfbcde6058cac4327ff9b50288082174c8c53a69a77657c5b852c6464c6e2ae67bc5f6b80ab5740581ed3f33df51d61b34192beca69334eede062a4dd0154816e5c8e2de11b648e5084ae24f5885734d2be2b82b9381a3ec292f0d1d42c0b177914b2ef1316135de7144be96ccd7f2c12710fc4eb3a59c5fa13b4e4f0f569d8eb52c82c948fbd87aff1ba79802451321fee7e3b69435fc527a3b4bcd9f602027ced3e2831538693e24626e20ba503e094078d99c83801fc657aa2d52f40a068ac4e1aeface2d66d2a411387bf8f5907c8fa801cf4b5c2338c6f9a21f659766ac206ae78ddb9d67f08e3ae5f971af89051ddddf01ad592a70af11b188ff5cae2fa7b8f24188fd9365613a03ea6152b6b669de09c6d16e37bfba3590ede01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7de527b0922f2c6a7b01ccd8f51ac7594989e65c9930e444887caea8ba7b5900e2d164bcefc9b82307f9ebeaa7cafef6850a68d6b79458a9913bbbd439e28233eebe8f037df07ab1ca0e0153e70c3964f6aafee11a46a24a1f8bd08c1d8eaefec46e8b6143b3a9d31abd666cceff67fcd85d82542af8389e092bbd99f09d2b09a294593036eaa089e1c853bcb3759f4e6bb2a5a6c92a9b2a061baea6667bd2a0154d9605548057b953cf3e330086730e935f4b78d5fb33cf2c2fd7d0e14c7549ae8f478bb47116d7154efa08b926ece36640bdfe17b65e95c8c332061c088aa2445ad1e8af2a30bb17a95025ac826231e7f2c37a991ad427457d6663435befe2b13cd6415b462fa62a63ac344e59a1d66d4917d95d9b3defb9c9577832572c4388e8aafd171479db47e84ba7364db32e92dcd7d0242cb06c5551de5cfaf2ea76a67b933bb2e285c9085dbb4780ef4c21bd2a69adaa69063a9c33b6bf605f3bc3cf27f947bd81b0d1a94cfe34ff4f40d8b83eb385ccd7ce1485754a30f81efa00aeb6bcf1b3bf4eab6b08f90753b1991faeef8d6b3a88a36cebdfc16c6fcb8d06bd3d6e46d0f0950c499685482efc5456ab1a6473c35c672311f3ae498ff62ae3853d8a567d42eaf9c7583dc80fa68be398a3f2b49211308ebdfec7d7d0e49b3ba05448c94d765883a3afd91beef94d90c7b09c1da6055658ea11e680366d7b162842b2f835e29f66f2cbd440a69034778f9a243adef4c537c69c062768c4d24a1244ca755f988ba2d3b7d6959bb0812fbda2d46a4600abce77f700f68ac6424bf5bd12cbbafb41fecfb9978c359a7a2e18e077a770d03778209a3c0462a28b0bb6bbf57f104ebff823e4f7662dc2d8caeab709c7f9eac1dad5facccaec3de98823489a126fad4237903ef0c389edfda862666a819313eb93f9a5670bbdbe6100627fa46f3e19c68c82d491fc0af7f9d155328290899fa24b2b115693accc1670e5c24b325932612faeaf86852fa7726a073c02edf336c6fea9f2c7d702080b81a941bdf53f2170530f76eba6316ae3c3a579639e21148dcfeff7deb82482ade20d2c20bf88366899c15213460dfbc69b623666ac2674f0540c3aa70526732e9dea4f3ed4cbe363f195a8d5ab3a5ec94a6f6c952c1ac87fbd7b5a9158c0795f9f05ad52eb726c41e224da64ee1b6dc1000307e37af9a7110d02f8682f1dfe39c0c92703e8827cda7166ff4296137e71196174ee1dced7503d0cc22897f3eaf52f8121b5452a44695fca6629a011bbb3acf8588b69376d50d3719c5b87a1b2d33fddf607f2845efdece3c7d0e466c9c001bb71d34b305b6303356048d2d28d6b19335f5bf105357bb9d38218437d389696a517066c96cb4f6e5f6436fb1eb20429e8500196ee40bc47e98d88eff23c70a4ac40924a947d9a3aa8f137cb446708fc00f5c7c79e2b0b1638764d3afc94f986dda8820aa0f6ad04314bc3f529856cb6bbc6cae8aa1dbad390401f7541b116099e4432fcfc7ad499604c147ed8b0ad35b70f37f95b6445f4ef623e5e5e03d2935d76b87d619eceb2ddcf399af994cde76957d8d1df080f363e367588c6939483a4da51e93dc165d73fe7463b77972c6b317eeb5657d5de582ef6ae640c1b6868b01c9bc3c67eae3ef442894d4cb38ae485a451ddfc019a450ccf26386c9e2b7bc76154f3c7e2113d8857b7cfd2b1a13dd45abd87aeb95f08f4707fcc0f301131663f807d4a5e7ff6beaadecb99425ff67d9b354075283139c0fb3e3244a4d1393106fdff4ecacecfe29843bfb09586a15115e2f2a9b132e847f6eb1eedbb95abbdba41b8f81c3a7e16a49e1be0f54e8646acbf04442274d903402d4b276a8c407fee459839bfb7aaf3b585f4fbc15c96233e1d40ba2f3273dfb28246a6caf9b00f0d92778016b0770da1bbf4c4debb1f745d4f4b80b8ae01e72796e973a5d1879a9e29f8b401afac14f8e1f2d454cdc5b4b3e7eb4fb4772c53c6d43469cb279730c01ece0a94098d1813cd4633f3d24b06cd0a9de2b8e3fb18e0f9dd6a94795299797cdca35ee5f84941c0dccc7295e7cac4c7f4b9236f680a506220bf9879ecc91d807eea8b4a94f00797819b760ac51bbfea19638ac33523970436ce13513b9e6191d7acf6355910a115989366628714c069e6ff4255c490dad34c89c3fa0148986d28c996db3c0f9c155609d749ee4c02b5385e66dc27e15722d8c8f161e7c96982624d4407ba568b2a3b6d95eb1961411067567a31eac2ec21a18f4efdbb1cb13a42c7ada150925f8415bf7dcf192774cdf9e6152972128347ba912166bd6caa3bff23c572ef881de958a0564de898f51c818c0e997ea9398b87a77213a6e3af03b682671b07beb855eb9264fac5839ece265b22e9ade362ceca1142a6f52db2ff94da83000e5e3ee6f9b27ac25fee62c45aa0bca2615a5ad170709142c1f8cff5d7c81ac78285fe0dd544bb3840953257e916ae7f4bd22f0914db79b241c321c7f7dda4cc3a6cfa31983ce2c8fd747cc7033789d41771eafdab3377d1a2e8a900e6ef426c964c3a2b5d0da1f38f6474dee744fa5a2e3e69067e119f0615abd0a5494351e72582629cdb3655b2845cbf2250b7fb279bce997211fa5c5fc021904cc39c26e13228cd5530cd878b11cd976ae931aa91e0b64ac97d10f11f2be6de0dde0aa2eaf59b664f73162351febb6a2efad3399d1f7ae912e697bc372ba0a6e0f8aa7caef5b60dbe2f8ee198a8de507e046be784f1fbd1cb3816b485a08ad8f6710df0815f9e14cc6d1e3b217555fb76946c318dc48fa933a07c0dea57f0d32f64094e30ac320e3d835af98274e39abdfce1cafb0a2f4257ad9a5e98dc8570f6220b339725ffaa8bb6c31572ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2a35b75f0ed9b2d0543dc9c0f26425bc4228f490b8febc528752cdfedca90dd769cfeaa58b0eacee0072e5dcc85550017bda78a0b1478e129aa609344156a84d359416b505dea1c8506b748a014fb7fc7faa1678a5785d1b4d35627f2a09296ac022c91097e0f31ad71d507cb0e952dd012fbffa84b54fe3a4bb74d011535dae1b28f00e3d47caa937dcd09430c93378dc2faaeca766f3478817e4ca1e8497359ad1dd00df90d621354fdbb98b4c7efdfce9d0cd31e2e06ba01291b6fc690e304b0e24f01c1fd4a9d7701b5917068525f440adf351419df036055a0dca28ff364009009bf089ec102eb1c4a2c6e31629bcacbb357e6abf49e1c6d003b4f708bf5621f89f3704efd33e79c8eb5db3e69fe9de01c30d1ffff653e1df51c8e36663b879848da3c43461addb5a58b85117bd989b106b3d208ec683b0607090a8825fa856c4fe87a951b0e2a63e340c643d6d282e060f76da17a4c7d76e5911457c499902f516bac0ba7d603ac4a335e1c4e16ced611c8ffe362103e4ced6cc86ed79140af8b94ef5a126794630ceded1cbb8c75f9091023f1c2e2c89ad68a98ff58c2a32d4e11f098cae90d023c71171b094af34bf402e7040d6e6766e190ee05785cc694bf91348c1944d2e0d7873722e0575a4bf51060f81b25f17722553fdc52ffcf7b1171ae9bb8b813c2990d296350aa67c93160bf938f566529b26b27ea2df92ad86959f332c5b117a729d6334dbef1911e8ea01f83f43031793b03e44f56eea72c254fec30ac8e048fac446f23d1096c21f2e691498b06dbecb160c796952f00509704f1d08eb98f24075a0d20ee3118c2adb8ded7e9747c381f75f73e3b1e9fcab60fa393ed80a9b2ef007e5399ffb0914b6e55d421a973f9bd46f65185965f6a1c1e7b0302c3fa7d79e8f58187ec436d8adcc6a0f8983dfcb5ee5b777167b19520edcb192cc6ecbeda094825454205ef3bde3f299da5029775ae26737c007d23b21175157eaeb536f037917ae2c297a9cb41a46fd33940c4968ca99a35240ea0a16b691a1e9a1922d1a98e46ece2a4040826b1081f411075e5ec6f119dd37adb3b5a2c4a5d332896bba292272ceee659866a0a76fdfa36d925abd5f7324f3bb5e9e3833c6f3dfb69ead4b9fe8a9c899179d86f8d29623f7407641bf375268ee7105c8cf0162ec1533a5d3b70e8c62f12bf0b3ec8b55d08176e2729fe991c916e335b3755b942525bfcb26d01b1e27d6ee48143462b02089f1f9da70c0fb41c00e8d88df04be8af9cf465af47224313d000e35bb0d6daa4aa4538e40eb48edfc12e5aff91ba9a60187909bef3cc3f778b40cd52aae963016c16963ab5433bafc9d0ae55f2a76f28db8570347f9c632e37df5ebedc9d4bf66e687176e93e67fb33e4b87d1725d6e3fad396410c0d95f229188390cf022e713e81eb62f08a488a0dd7f84e740d3ad4a026ca050d2b9c7636109c2e0760bd81aec36b39de18e28b831baa10b62e353ae47af237e9ef2c37d6f3e7cf8306c6397b5c759d35ba0e9f1b613e3c09caa81e7459e7210e77f9a08701a302cfc6ed8cee94d7bd7ea4052d5cce646c51a8f71042099fec83f515400b9a3d9daecdc5ba0edba4ba54de331c364902215729ae155e817f93352d16e8bbb1e15ae27cceaaace9ba9829e166f0233f8e5500a3ba914bffe8eb9216d41a316f2607ce7f9df088e1f57350abbc54486130281741dc6dbed17755a167d84c1b0572fb2a259ae1d6b1af2bbac8850bb476cb81665e3f48fe904142271c421533079f5ebd6209631a38ac92852b88de511de327d207b9e0b6305cdd80223341416d316a2c4dcd1c37f1765f2131d7c4fc869b93e98d1f8f580d1e5aaaa2c6c0839dbb85f507d971a59944c030d0a46d667979fcc9c11b8a4a3b5bf6dede1240c10b85f4a76481eb4ef5c7397aecbaee3c2280747cbdded9625505e10f0a32da3765562cc13e038a7fc273511a860a25544fec80c48acf7982e96a087752ada78ff51ec038c0952ec82c8016cca269d401ba371c43486f52ab23bd4318e76a2e65bc9e547fe7eccb53139fa585c92055274bf849f3adc217cc6720b0e4a940858582a3d34da4d37295508b3b9cd4232f8d34874dcfcadc205e9e565c318bd0d47935d47342c752f0696d0c1dced0b0b7bfcc0ada2cbecc35a9b998b4404b2b997171c653685d33c774eee7ecef498e4e156d50aa320b7b2a1b89ecca00df78647a429b7740aca89f0b2b927fff36d69046ebe98acc71dc277c334d289c60cc78f5babb94c89611ea41e55163b5294775de9a595bdfe0d16ea591f77f2ec6524233bb18a2cf1c0371fee097f2337a4306298024a7814a415c9ea9d888e084e4f0dbcb1ecdd49400a913c3e0e8c9626df7c959104aed96ba832f775b1e69e33c436dc34a344a0959cc26e88a861f6f01f295a775139f852fbd91e6bba1990b97f92eddc27087658991f612358f912fe10dc7fec70f9f8631591e675c02df68110750f5e1d613fa7ca0f3ea5979a2bb54e022e32daa2db0a89d5baf2a29fd7a269b7e1f13bfec59e51b85ef05893f960244d794e6e7087ebbdd7b7831e77cacc6e5487188866bd307690ca8a9e180d897b5f8ad77848734f7b4486fc34e2ba05d9fdf5f9223fe0ca04f35a202ab3da0b8efa850a7be3b32ce59b96b80655be09d834d9fb8cb7433978da8981c91c919c7695d2d029ea788d9de2d8829d598e153ab0f3b3f1c2872dd9d7814e96d0b090481b8e2bc937fc01e6aecba604e4d9d92298146ea4cff5b5ae7305a00b27917c1826f8e4fa729be426fd50b90664d84679f0a61b2b829a80553f3057ce6d8c22c4575262e67f738f2823ec485bb7556ec802f39351009569d3a458f0c7b8588;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7870812c035c0d5fd729dfb028e90973295c323f0c8437caf459e637343ab768c37afaad1c429f39be10b764ebf74838b7a1eccfb5d86150d7ff67a0a1961da1fad6cb30c35fd37a0aac9602271c0b28533e21eb4ba4fb41516c08be496ce3df359bac3e1ae7ec387c5cdd620bc57a35f025ed71ebb1314598b17cf8283b48380e62850cc1a32a38d3ac3df2063ee8f4069879a0e072d9f847f56bad79f41315b0bb1a2a0a5371865cea487f10902b449dacc9afcf8b83fa5159992225ae5b7db589186dedcea113fa30a5ce85832929a965d426f6d6efb13c30ed4d65b199f7ce87ceca2d90bc01e4c0ea6e616a148c9909e49543746adc7bcf69a871fa61d1060f107f2a14f460c32b4ce63d43465e14c4988d06015f9926bf8308e9478843d19593f945e6faaae7eb93e67a25a103a8ea4a402b2a8c133efb355e63df2897dc4e1636e7e68cd63a14199317c9a07ab5dbd13333fe44d4dd6f758f3e05fede0c7e73e5765ece407d6da685b3d868fd46b5cefa80378ccd461bc7b18ab1a10fd2ca2e7f4b8e5632ab7e6637f260c4a88ecfa6d6350a0c8d7dd52842983e47d319a7f3dc2ddef39494e5d61da50f64891372d0554611af987828d3822baa027d853618b4171e444882df50a32e8f8e02988a8855fb2ebe026c0a872a5bc635728da2f679ebd89a702df22d028563b8e653cf399be412435bf707148075c4a8bda6f10db61d8fd5f7aec4e4d08d3528a8c6c40c947d7a1b5c7b02a1d57e309f4d07ec02c7584bd054113dfe192f5cf4d2f00e81334f9d187d8bdba47dc4c240388a69aeeb333248a0279611dd0884277a98233a575afba358f2915c9b538c969c4c000e7735f77aad5f526da39480be81407c9101b773bbfceeaedf49f3377094595dda9f2305780a22a0193b909ae3e19faa17b9e3fd1bf795cdecbf81790c87d6d5f02a4d33a3631b95bb7171454c432edc1e85a7f77ff03d9a082cc60a55084b2ea081a547a30766728c179e8fecef9a4ef38c3b856696daf69a9bc32d170e325f91b7b381cae958a961ab156b3f8233f10a95e83d4b4fe71688274e2ee76164273dadf4dddee44f4af841a81bddb70df57fbe4cde262c0b8f74931c1e47085c773703dd6ad93ef1126e61925f3238f6caeee74c2f552db1ec1892de2d29b5b65bb5965404c3a801a7d30346fb6a95f95593203836de87a3da2e53bea15c67e1b9dc153bde73e4ac88c61deb382c86b2b83d8936cd6d47ab6d7a01471ae342af5163017187a631231d434ca8dd57bbfcfb52d7999bec5b1ccb90184572dc4c53111db0a2a9211349f7239391dd44ab477a0839181f0416eeec5e579fa0c088ea10c22ff84cf598255b914276218b91cdd2c4e2904e3e22bcd6668f9e895b79c5fcbd07c04b504b513ab9bae951991eec66bf8f8729dc3019661af63c14a12b0d76a1110ab0d4a5f8ad38839c7be3808dcc0238bd6b7e28760a70a0ec430a6df1f2aaa769b4cac1accbfa7c8b129309bbfe4887a303f54d2b6719b201f1369afa5dc6cc4b55147b58141b80e337693b30be6f1a46e56dfecf039cc7ff63a6a4576da3cb1ffd6a73dfc5798783d71c43034608070b0326f8f8d563053cd2275a7b8512ab3583e96626bc2ac0db31556a0d2719dfd5a3449b04a1a877ee815df2e7909dfe1480cff922f3e9f3eae11c8ee9cd68ef0936940045a01f80972c27130e8967b5ad14d2fcc4e3cd4112fe5f0a25bdddca66322028b4b0934f65719461960d0a6c66d147bf59c7ecd16572a73bddef5b8fa89ebc6393f8e37284ed68260b6022ca71bcf0fc5a6804206c779794aa65a7b1c870d024599425c6f55ae1bf49e91caff14fd7fe78c8d31af62ac129b6b98f6d25ea2b157109ad321cc9ae0f6665799045524b216acf9dd9c8a2d416819178911725efa39ef9592b781876de907b3bb37b9586e639c9e9f179ebbc1d8d14578c8c96251edbad0d975bd53cad4f15598b54ae2e2d31e2b82ae98b44ca8b1ba974bb60bbad7c69b4e650aeada06a546b1f9c8d1ff5dd064bd03ea0379e4518d5717a0e75584e2c3c938f02d4cc2a9ad0b21ea19e11624167eb644c6aac497d279a44eb8ef1717c198bcf077c1742835213ca333b7563dc673464808c4632b179dea80614a3d5dac802dbc95b3f339828f7137a734340579c76f32761e876733930f9149235fa021e6caaedf50e2b08ffd5c92fdf73e80124dac94ec0f7d9a7532383afa7b455056dca0df0ada1c8f7e2fe41dff5911e030e162ec33e29d6bcfd01628fb1efbfa7073572553208ee79038433670a73317a4e0efcf89d7fba0b6fa1e4b3532c919b17eca3623d9580e38c6e3e1c5158cf7f8c0304d8371c7b9b160ecaea62da9c55adc1b606306ec7bd23645bee338014100fcf9a2fded1ee175de0133ad171ca6576a0b38902df2190d1add301242115055b656b6016e88ebe83c1518f6355b6a39264bb8fdfb2256d771b0e4deea8fec979b66ed5055cf09d23ae159a246b58539fa8d694f2f542476bffd53415c1769b7b51937721e331d7ded59d7993e4a46e52c8871fab4b4c1540a09c204366d1b49e31891f9db4cef8025fe8b3d387ff5a8c13acf915a1c3a1a940906708dc71a39c12ead860c42537802611b7d3d3ec2bba4696136749c06c68c2ce0f583ea2ef17d83f888ce9f00cf6808eb3d27fcf3b634aa79d3d83cdfacdd650be5adbfd68a1cd0c06e8548e422c89dbc8f27596084a03280dedb91abff596a700c6f3e1a13af435daaa6b5c58c97ec3997e973f0db80b7a892991aeb73467a7175c2ea4a325aae21baa75db9b562abdcfb3467cd059c684bba24159ee408f0b2f808ea2f04d643ddef5e13d472504dc1f5f8e598dc4cc6a94b55b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h979904099c67428f9df28a067d68e9c97cc6c75883416283c369b00f79df8b7e479828051320bf3708430fe6926a45fbc1d46f2415b8dc9949c7e09fe3ab83d5bc7533d8b97f0e0407ceda864a11639282e2673901ecc663e4d489a45f1b24e1ab01b5418f82e5e0125c71440ea9e727c29bb91036ff3054ec98538a1ec1c68c8401e77d1aa3dc1c18ff1c6dfb0dc3cc311dece2a8fac10c61911cafa5e785c82a750ebbb41b3c69580b38cec6557f9e1d9ffe8a145737d18dab10b2280f7ce9b4e81ede9f800b2dfdec48959798bd26b8bcff0fdcdc6eac4ca2ae5a96d4b801d19f816e56806a957f55d910f58464ea6534cc298b2fd8bdb0a3fe1f391a9180acafc7961ed5fa531517fd43a5237e475e57001f781f46667238f30a535ec4865d03af206bfe6a632657dba1d7f3db6c566f6dff7392d8644fdcd18a81ae3e44998ed515b09bd8d839e2573ba549441ed5e60b887a6f4e55473245d71b202078e4c9fbde921d6a3102243f9d3b79b9437b7cf68b43c3c06b00254fc67113273c7193bacdf335621013cdcf83d9172ae227623de48600d03f366e05e92f4cd7bbb28f0cf46a9a08be06c1df268bc482331e2e223b7085e0d054679ee221d69f477530b7aa501bd5f7aecf00540516211fe21b497293d3940cbbb128c84058fa0dd92731a32fa2cb5c013c2763202991da0e02754e3a5b2a3fe906bcf3f20a75eb4dc681bcae6a563056b837d96388260e106d75d43eec0e0426b91849b5c481364c17251f946c5227d82ca85bfd2c2aca5b692426d8e8294b3ee05ec910e9f81f1c5652d34b629159e6245d53afb1739e218d13637c3cc3d7c7b35f96c12f8ef9929938671edd4579a24317193890f7c2f04f8fd4887f19fc7c133f51ebeb3a35ef12294b7eff2cbab128858bee8730ecfba762d21600e96fed71923bf986a6383cd22240df622d025b1899923ddf4122ab81b09999cbd063df517ca80708a06e3623423edb24e414d7641f19d17283ce43e36220d73f76f14645830581c4f537bfc5314e7b09d6dbb1ee51141be5c88f1d6f69935a607370070a7a1c00debaf4af9632440dec56c7a10a540cee91e8701ced4f0d62e8d59d37a31dff75045a75f01217e78abf8584a8715eceaa1d034487848be04652e929b5a9df2d3d2a9638717ea9c910d06763b1893bffa61b7a82590e8868b862f4ff1dc9bb71e81b438943f6cb98986236c0f63dc6cb8fe4868f1773133ca74253f273e2dd93dd832ecd71fa67f6759f0a2176480a7b4d87344aa6c298e496501d1bd01ea39348a3a2026186d0a20cdbe9181ec8c29fc9a898d4a9bc15d880a1f65fa9d73ad7f87fbab8cf499e3391a21832c16d838be76cc1fea18423dcf761a161fdcc5766013d8d7703cacf11853a33448df1c793bf3f8a846c928d04dd30db4816eac6dda2e59ced73e5ea9942aebfd68879026fb8b3fe9d6dcd6c0af8620b7bf90df87adbc70301f073640ae15f8773ae432452f0e770892d3fb396555448e2ad02aaa34b6e3e84918ac67fa367cb471d8967d1f8e092647d9da1c6f4d749f64462217d19889b4b3a48652abb346a1fa3b5b1949ae5d31fd612c89d5cf5a3be247b740b94e94b940c4e80a56c1e5a602c681e9a9daa98f20ca739433460bcbba96fadff7039d4c8327c35111dfae7b55ad34f1e2e93ec57bd499d6cc9da66d2698cf2fe9203a7640106b8e40d3c7a4680a0d6a7214a0e1cafd348b66adf2def50ec0917cf953c1d02fee7e9d7bacf54039b581b349268f0344c972bc8454dc3d077edb2e9e30737f692bae191e5775c82d5b15e11da75a2a3fb21f519420120730d63709f49a2db3128fde9c46447d80f0042245d5ce85b52bbee911beec3d9c2721f5e720d226c4811f5d195fd1a9e2995102dbeea19b105884d98e250a25947e42dc2ae706a244001aa77f57ed5cf5e3a35cb5a3d47396aa5f895bf2c041439cc8a764e008439a69088632558dad7c50e082b8a91fb9fd78263fa157586f66cfc00d65167ac9cfe57042ff89d318bd3ea6cac190dad4d27c1012821fccc135c8586ccc063291e27b742f0cb06047b37337394910e7612a494217a4aa9e31f075ec7a8337469c0a3c433e6f30d32dc89d1bdb6eed98c2f5f61b0e86de9ae1776dc704e714cc3fa3e7f3dda5defcd5b626662998671c2663a7e9f69b1ff981a4954b3cf5919d8b676e9f167303c2cfbe628fb7936a0969f5e749cf99515a050779d513d083422cf68488a91ea92957acb0d0d73ec5f9639d386eb8b5d737e70134a40c3ce7bfc782a5944b214293f554de922051be2b9281a1d6937cd4218b2a524435ae9f7d5d209c22c4ae5c1cee0706309f4577c330a64d1acad80941ee96d9a2d67c6a56eaa9f208a756664ea9cfba60c0f2b3846dc36afd417a88b458e25a07a27897a88465b8f5de4b76e81afa0c4eb618f8b94b24d36649d90e2f265a80cdec7f54686a7cfdb2f157fd92d613f88de38165c8fe3b85548f99bee4f95cad82b568f251bbda912f3bebefe2f75daaf07f12d52f4643f5b7407897aa5f3da36d49595dada5e2ffc4defa57edab86ed49363b5c55fb874f1f77ef45e3eac72185af9f197659aeca505ad696d20dd44776f2e3907b6576b4ea7a5052bd3741f6f76b41306949ccd0e38aecf97f2a9e2b8826c6576ab09ee38e0c846bbad0423060461f438446f37b0253adc946ed004830110c36a407f3e969a5eb014b137bb7aabbac4345040cca6a71c020dd85195788f8be1f81782e83357438bf680a653c755b468a3cdd00b754c598206475b479f0a691ed8c61138b00a14f6c6be0334770a86fdd3aa6d7dcead6034ea86091bb304b46a6f8d1c5a55f0ddf2cb6fc97b5384a77a64586d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2dca659f4d70621232d5bb2d2dc76356832a1706deea078ee44d546de89544d31b0ddf858df9edb5449643f1c31c5c696999cc70ea55c5d42a0c97a8dfab4c7e300b2d7061144909066ec1a7bf9e921b3ddf17e22494abfdd401d686445a5b5fe46b927fc3e2ef607e3038dfd64c2b06008cafafd4354384c41d554e379b5514a1499ba33539aa6e73a76a9a3c5f2c123e5ec881ce056fbee5a505505c306625d1e0590eaaef9741cf4d1ede77d583239606d19f403a957a095a6eb8ba9b29fc40f9e4b14a8d1681aa009b73a13518b7eba0dacf9d6a36ce7c02401e00933fdb760d5852ec3a6fe5b438d59a96f04a2a8e9d40ce7c7337b342138982010c15d8d7936104b69f8edf117dd474f0b80cbf0747af6866e6fc0d6a75a84c37a06e2b38bb83c75c74eb08de6fe49fc54c02604ca97b660d0443df1f95ec3694877782b93bf387d0e055078864540cf5b0a2e008c3ca7c9eea09f06f937dcaffc6f816cc93fe3eb82524b4f4a536592082ac00daad56859c4065f0b1b9605ee6e04b45964e08cb60407ba92840068b6aed17c0071cc79f112d837b770e936c359226ff21be26b3f91d198f3758266edaf524294f3cda0d2ce1e19364b416a06eacad847dd3386f4b5e0ac07c0b87ddb10bcf345b4c2018ae347d1eee4cd80ef47194afd265146b1aabf000baeb83c8f741e09977173eecbee5fe801f84c17ab82fb9fe29529663e61975ef74ee76d44409f476a99a903bd6501daa43d6c496175c43bd6adc74649abd60f850fceaf27e03f51201975882071763356ac65705fce5c02292a9365f537b5e63eac21d2644e4e5b50abe2fe4e394be99cbcaf7722419c64feeebc991c8e33e1337b102b2ff91413e3fa73dbf91a886fbfc9f4b9a45ed85cf23403bd27e42ce7978f98d9e27f396c25c1be71bf7387835bd3ffbb5aac0f595e8033d73a83aac340d1c49c776775fdbadfdb7770e61bb0cbe5d8fc049f7173286e8d66af788af75b66850c0165d0a1b4aadc9c5d4cccf931522a6f539ac372e77c264e472de806e6a6d4c10e868535631a1af773b012a3c083fccfc61de6875af1051b3ca9ca4bba7342adf43e2cc2f075dbb066b54bad9266c36adfd0bd410d7dc05a642673ab88390425bf29e02a66e136a78141b1770117c0d11b6640bb121c9671c414a49615f98c6528ec691c4337b777e47f36b8cf691aa2200e3e4d66c596d50ffa7042113e462c223e39db34f69d5e1464946e8b1c539dcac412a852a31c05d069e51700888a613e0456254577bb1de180c782379770145b40ba53a775657b02a9a4d983c32192a627f5f93a376bb0693b18a76fb8610d5d92e0a3082da8840aa10dcfe7ee9d040e443f9cb446f0712232276df23d7d76026b6eb6652c018e0032bc0dd54f438c1e65d5bede1e0578a20dfcef89c33d07a8fc8f059a9b66d79a0f25155253cee47403275884442f532405049ab972960a2d97e5d11d3e0638a11c71d05344630dcf959ae1fb1121cd00ed34704bbc7eac74b598066fc09566703e3fae47393f5f96365a97151e23640359add02ac990641853c7cdb66eaba221137f55e561e39e09ba0f2c595fd534d7f8685549188afebed395ca7af3c86a657a8e88b48a23a0fc4e30ed1f25c45cea314aa299bbdcbabffe0231d3d1f6dd489911c7b1b3cd33f58c0f2bd21fc8fae4a5146297c0998d47ef48569332a290a24fc7754a046e9db44fb947346cdb34674578ac153216b46945d5d63c3ba1619290a2b085e9e2de3d685ff652ea56b3331ced36facd9d23bb9be10454765e50cd805c25cef92810a6b144492e2cf252b60a41bb59d44d1522a35a914d749bfb58c917ed2967b6e5f71f93f982637216fdfe6d4d3344b56ed03df714910eb1f6ead785e698b80365edf4ad66c5da1282959609f465b8ca505bf68c6f9aabc1e57ed47e584ec21426bf8d58730c8cb849982950d359491c0728741e77d9a4ad3b94f6272ce58cfaecb6b74908e99795ebfa2dcb6ebcf014cda13da7e97137e5c2ecffa02d72ae5594170a5b80be4b6a398ec2796a153a2bf324000c6083f3e170c69e776aae51068bd353a37ffdf8d1bdc5473fa537b5596cc7e057e58fc381b60823cfc86780f05cf9e8b6050a5f5ff4092cea90a8b289eb559b89ac0b7fcb3bc88efbe6d4c9a229def8a74d7050c95bb87b2e86c707bbd3a9c80e0aa698a1f8d38a02a99194d2d1f12056201824981fad0d62c3933c5fb2586728494b1ce9229b404c00671f15238e85d57125ad23098184c552f0ab18a2ad16043174ca07add39e9446fb734a2fbf7e255b1f1761b4fc37ff12b98337b733e1a0b5b5d1b2be954f8ef04f02f57a4d1baaa3bdb208c4c143150aa0397c95a43866557578b1abedd63cc1c453d98366f1b75ba9a88fd28a1f2a75f58a65f8a4dd3c1f548b218d5ff2682247fe904f14f081e910883012612493b34e2514e5502731050a6176f3c69e183325d870c3bee2f572f5c7eb612376090c3b3b004967fd1b1aced24829536b058989ed98ab03e2370a5f7dfc94674d36910cb7ce93b1b66540ab8074cc2bec62467b1d9806b42aa8a8f939276e3ea1fe81594511e74d3310ce31b4d39604c8d93f6e977b7920915aff6819ee85cdb30221c6bb74e8d43d65042d56be28c01f08d9c27c2db7902a37bac6158900545ccec3ec19e21daa177887ff3271b5b6fa404feb9bee01b562886e6c315e331e212c9783e2335945a66f62f7374887647a28f94126710183b5dc07837c2193fed549ca93fc1cac56f1ba17ca06d57271946d59d2f5c0233864d773522278aa2e20896d973fc76abdea458edb49127d92422e3d0b1338211d8fa607923fd8b53c4af5936d8d102f06d7b34e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h74ea080093e85dc0c17ff43e79163db8d0b7d785f8654268150fc113c9b2d7dee89290834b5c9dbfc0d4a11b3575d8af1158d3b1712ee26023716506ef7ef06b629d35d31bfa97a8e470b6ee8637ae7445bf755aa6a9bd06451d978c701cc024afbf3adafd93c82ee3276d91e0361bed6d1b6dadecb2818993563c8bd6a9c26719fed8db3496b4c3c57b5aea1508f2005b2c6c24aaae5c885dd0b4f2e85832df514427f4e90367230cfc70c1ee737f1ae2c38c6b72aa1801fc289c16ab637756f8124f4ece876cef3a1b1f850b41220a9edb37c21ee466771abb61cd3f594aab66076916ef99ffae7eae90d274a861a7763c6487924f780baa154b6b7c934f46b6d8ef2a0d842b5a395f7dc2befb752ca2373dbc4617951d2c574ca2da92dc58fe2d8957d7ab1a71cc31e03f3f02f6de20f7ba47629f6e42f004f7d5010c203ff2c0c10578da3926a7f71925358b944ba3d2a47f5895368ba35d7d786a4536b5724e94a3f85996c350ec1fd68979f4f3e01059a3f24cccf81c8a08d93efe9067cd7fe8b86f39d1a62255e5e28a9c1ac207794fad8214179b21d52f5c25def34d7d2e7910a77082a109c5e59358163ea8da62d2632708dfa0e82b06019ccacc8fb67b4d4f8297f87b4390ddaca25b73bd94babc8f55a4656d37aa8dd53be52e683e4549909e6385cce85d82e5d49cd252e41b806dc76e138f169b48847509932f5276eb50da4c319809d69254a9ee88f228ea533a21464881fd625ffd9487c9cd790d1feef6f80b85e6b450ed0191688f9c68223dd7eb7e85ff7d33bb041acca4f18bde5819473b501cbdb6f476ef00af7c98f6a8ef83fb5c463a47adcb97a4087925216acad945e8972e1bd10ab530a1cb7f303eb61956a3ff1d2b62edf081e2c18e956713bcc7a32ed26f0e4184fa2f4f09c629d71b8e80b4c9441833b8f9698f69676e9a2380a194f1bc3c03d4c6381f52a17e3034a9af55644ee4d2e3a77b203e1a2752c9e565bb5a9d39d68d1c1f9a46fa5923a0effb521f4c8b7918a09709871559ad79ef5eb41839b5268a1d818dc3a7137939263b0e8b6fd32b5bd36745aadf6ee65393d3707f004adb4aea7f3453ea04087e950418e475362a1a499d4c45acedf3f23ffe8848f9a18c347090cbb57afc98613b298053d302b92b2d994f34a525ea4b71695b7b8797077f54090c699ff2355ffbd8f50171d0a7ed0b7f86bb563d382fb2dc5d0236e145a04e7343176b7cc1566cc4caf6a282034ea701d84a4f03db1eb480226e8d468904a4b4d450ebb0c042033c70f9c3414eeafcf4961df5cdc6562b299bd4ecce1d364c2d1c2a107b689227f3497fc131bbc3732eda33830a88f5637a16284ae22b034039ba6829769db11e0cad313ac14e3b1b8cb69816b05767fb7c477bd46203b4432940f2098ac23f467ecaba52ec10761cd09c754c7121f970da6e19b47aa2a5689e1915f1a7d402ca8eee0a64de00b80c8ad2d519d0ff5dfa3411bf5298c22901ef012dcacc3069ae31664f2689edcb88cf49049d076236373abfb3276a4ee8d5eead6c934f2b6c9790f36ff9fc80bf918b3bfaed2f95844a052bb131ac8ec35093a5453e829ce4827063592bc6729060ecda3a0ffc69c1b59a88235e69fc831857d1aeef3708277e74d37222c5db5d49cb109db3308ced05f210696effc931980e2f6e49a21e4fad2a89e3814abb26e27ff4b02e6fb936849f772647824296c3e03f7ac506e33808edd2e0e39f530cdd4120b3532966f5853ab951863f993ffc64cdbdefdaac160c800c4fbda7a8ad77130399cfcd36b112e07836156e7e8291609494211056ea16faf168912ff227a26912ca57d6b95509e541b94b6c0ea81afb30c86cb8c127a8411077c1549bd4ddd38d094f458cf3d0ea2c2dc2c270276a078c0deb1e6309f1eb2ae16c38e0550aa5151a3c697828997c5366d61137708051b85f9116e7ea4833b604a4eb7acba54a6a570f0ed173b11a62876501ddad07f5b305093775fb31edab9aefd2d34723e576247cbd8bcde912d8d1c0131c79ac39e57b6ec0d4d24e5c6a7e62f62dbab0fe9c0e1488807cb24b743bf742496f565a1764cc84bffbf8af3c8b838bd43eef05ddac715cd474cce61dc8f0804fa1d67f85bd32166a1586ef7cd1fc8236ff40f8d78db6a201befcc97a352a4b270f9615b2040a95a5dd803f8cc231708c6f673e4eb9183cbf238eb777c49944bc7e84d8be92c247ca109e48083c8dc2748e947a525a272b6c512279c13836dee067fafc816d3a38cdf6ae66ce7b1cd2b1cccd68217328fb32a0c901881431eb4cfd76ec1ba2d5da2763a8e22a1da46b13ce4321b6dfb38d49e6bce963d9b310f964937f2fa90c8e61cdb38fb4e12329d8b8c15b91b2009186104bf8f9a4c398cbb653567dc3bd48bb70fbd47f710c649eeeb6c1bf28e699a7f29b6e467338c14becec9c43c199d71743aefac5c77e80ef7bc3c1d892da40dd4f44469f15b4c607792d8c93310d9795422d4b28878641339882ff1dd3b3968f171f0bfcd274babe98a688261c5e9f15945812f3f5ed53bc7a032c14222b7bb93b1ed19435cb4c761d38f7ce17e02160292104f3028d8a1b78d5de545c404bdc45e2a384bf8e39e2062a2ca6db57aef0ed61065cf0fd87ad06199888e2bff8b6b79810c07a623253d901a4a39f167b167af01a1fd934e6efacf7a1310da02354f9e02f19ffa066c77a7bdf96c13610d3fb52eac0a0d2b640a19376a9ae11b40e93e72734fd52b586d639d5266b28d56ee246f8d61d4aa6449927476b57b2ce3698f4e20722b8e9cce7df801eb147cc46a0b386d47028e376cdf1ba6b2ecd5ad36a52c8e2e48ddd85f18e76801b996ea69d49d00ebf6e945ae8c5cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hea8686c8a6f378388db6a74c24627c5b923b204e0fad22847c7d0f6ea860efbfd95a4c6bc0c754998c1aa5932da3631f0ec657ff458eda12083251be99197b74a379e21bf36299c618a530fe630d0f19ff2c35d348e2eb26525fb12028419d474b10473249ddd0e2cf299f64f47fa950f7ce8e37c826473c91e983afd482e903da7050123d1f129b579c2eced0f532232f00fb046561497937b67803d8cfdb99dac55228d2cc316aea4947a64a565fd42b70960cea13ededeb6b3fd05368086f9f86c29d21858d38cb4ca63ee3799267c93181b673efe6597880d757954338c3de0f45d48c7c6f6324c2babfa42ae7672b942a156821618dfe436e41739a78cbdcd5b792e140694c12ea7dae8016202a05a1ed1cc3b05872b32eaa937f449c672608910db1207784a7d99ba45475b6085a54b3177ce446e432eebfab23ec5e59794e08155aaae7a110a1c4afc13ae1e77f6211298b651c565d5dbba49c8e4987e13316e0a98a9b2038866f422eb9a0fb7b51da9bfd7893ed54e38ada80e5cad2567bf66e86cb94f9e075300bd6ec4da17a94d4e0897b281d150cd91cb88cab8c114ab490819e8e9577541269640e070989c13c379df115f2b6e140d88a60d883a86f9dbbe728c4c9be95a70eeb84fdc8a418291b95dc1c9ae2702fdacfb187ff140b9d4cb364244b111552ae511b71615a18be5be7c7ea6c96c14bf045ce52058a949f0bbc9b0bfd4034eb245f77157f37eb1d10d24cf9e9e512fe74eb8be22d75b29aaa5a9937f9d1575d6369b94b858b96a8a8b3f0ae50c0a2304ad7f4571abb38be43cf57661b8a314c9be86912afaa74cdbc84e189c6a4b86e90f53c9864d73d0cd468381c728e516fa1dd5347b3bfc95ca7ad7f40110948b351e991fb5e6fa518e0dbbdb3f006fb194001b090a019b738c6df3d51fa71cc20dd9de6004e43b994a13c24b404bdcaf7951786224109048e45fa9c38f45a3b866eb6ead98cedb541b818d67c5fe5f7608db44ec88716269e6f27340373474ed3993f45ef0f78abe3fa76f4efcc576c4745c728aec65d468bd091ab86fb168987e5909af023a708d95a1ed2388677602d86c84b805aa6f2bed6397256592ed2d5dea3820073b9cab05574448c9b451a5a687731b7c1bbb34f39568f58f41bce5f24609073b59b1e070091cd02b9f2d17d072ac5ceb81b12dc3d05f5ba87094311e3e482d8ff25c0e781c05855bb55f622dff89e1617fb0486538fa5d5d30ecde8345bee84bea0c138baefdb9d26d6e800bc107971bc9499f7f7c9182fca4570b1d6f4a7c70663ed4da1617824693efb7dfb20b9ebee9ba190af3fd1f002c63539adc492242dd30253cf0d13cb96374a2a4d64b6f686aa05c293a77a9cc4239e25e65ddbb8a6842677864d951a0132370b49539b757f2f62ada824ac27072748916f6b6fccf484c8ceb0082afb04b0f1436a75f299305df88142335e0c4ede77926e31adcb21e9a3f555edb2351294f0ad1ddd83bc330ed98caffd787b900b676070b799656ea3f21316425e95346b8ddf1739661fb7a257524a883664df3bc4ea203de5c4cb43516ea8934f9828713e9ad6360d2d38dd0b3684521ae6d031da351a48c2f718211a2188210d06cfca1bea77c94cc8f5764a924cc2f68399d15523adcdfa198f9cd829c3cce25f21e386faa7ad6e75d1b3552c1eb2ca5c2abfdc13327239bad22598253a2ecbb49063fe7325ad487a6f6bb227ced80fd1ab47a0e676c2c7a4e5e61e0028a5c0646caed7bf57fa36933f93d612311183f9120e5bf26c8fdad2fcc9b5ac55f59c2ce8a2663382491f9cb27dfd8bee861b5334e76403294ecdbcef7c9605b49c76bf233ca137112b30b4b2f37b0796f141e349c64e9f1a2e21a61daba0b7dfbaae5406e37811183ddc2209d800e67076b88a61ec95c5f1bfce511ba8bc934d67769ebb302eb4e4c68edc054f873982ce1fd8e4a35efb3b603a53dd66ca2d5984cebd7acb143ba6173faf637ebf93964bdf8fd88697d982cff95e2e62d95f039ede05f7baf613e2b7295d27c4ea1c392d03788577f175a6fdae3e27d117151371ac2fe6497b7b9e5c6bbb10aa4e56423b8521cb42c80e5cca30763dc605f7eb2bcddeaad7fae52379efcb074a9ccba93e218b8527aec7494e4087b3f198e7c8ff14d7c8ad9ae611f0dc01de041a094ecdf26aa0d30c2ca2efdc798f7ca699a45311333bf06ac242d8ea809a31c95d34902e7c5d64b0587e9cf4649ad03b2908f0d1f0ab9655a76d2a4d6d0085ba4167a105e5c15e3c7e5c1d8abfb7dd840b44cfaad792f6d3fe88922f168812029d617cdd75f023c8c6e72e5defff3c48faeab4596844a251052b5d407d65003942564f095b37061d94915bd1329c91608828832236ad06d3571d641956373fd8ffbd991864338bf2ed3b7f752efb90ba25fa1d048fdc01c1bb6149a0bc4245c547fb28e3e8464b4591b6940d0217d2fae496ccdc4d9ca603581bab1957f1a7509ffbab996089f0913bb9df45f981f102a27c341fdb797a0c1f78206d5de65cdfc3c5696ffa1cb64eeb1cb33c731cd259efd3b4fa055b9d96237eda903668a877fa3796301a18083cf301b0e11a235414322cc29e1292ea3f45378d7852967863615d0517b33ea22383e37a6167b06fdeb23bddfeea6fb3aa244322d05666f7140122a5d9e1da5a63f01d9820b2eb67a17577577f47a6699bb30b8eb26ad1664c52da41b64cd5346b706e0141ba73ee0783ecd5c1362e129a2b79065f0db45a27ba961bd4bb206c7200dabca06a2d660461536f71189d52e4006a7e028c6ac45fd678dad603f5a40ae6525d5f5bc2ecb82f4f551fabeb40af6acfd483adddcf286b957650ce773bdb13d5b769fc56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h657a61da095d0e8050f1757f47d8e4282c3c77354909c5e4b93117c51892f47109adb1487772527be2658f0b74bb6580c932c77fed0cd3c25c8306c1843e8fee9f70f0a7bb544087388ce1f7b7def4b41f1d93ce45311b3996c568b7abb27cf522582d8abfbbe44d44a651c1c3ca3e6c5d93418c337b4bb1dae5bcaf3e3491cc0ccf1f545c6c31a01f4495c48afab7c59b9b44b0e2451dbcb49c28682905da05663a0a082ae4fed9df533a950bf3cd5a93264ed285b3d2f44d8b310167084515c415efbd9fffbeed81c5169d78443fe91f8352a7c1ac366e6de7378501e0aadf915394f1d9faa087dc0ea92685d12ab86dc10825f4822225a8cc22f6009f92404df2d5d79b13568ca2a7bf12862f12d27c600526fb17171d4bee9e8349a42d0e716cc33c93d5c425bd6063ec90b4aea5ab9186f410cef1059cf7fc32fb042a29fe40b42c8943a36cb003ee01d6b01ecb711b3fc3a70edf12c05476bee3333c7008df61edf752d7b3f9de621185ea0f442bcd0896a4db38e3756eabc083d6f3fc9d678abf33cd92ef9871c0a4c00555c3e774229dd64d4ad21b355a1d0da6f67bf6258a46a0ce49550474176b04458302fadc33ff38fe88ec068e142936372ad1096a186119b178fb287189eea6b2572177b3d95a594e73f83c28d9c490378965a888e7ccb75274e7034b701f153edccc4aee9bcb97b401f8ab8eb804bea9604283443c564f075127fe4feab8e91293732d299ccc44d895e2fea3505156a573f3ba3e872603387a1e3b8691b614fccb88a02a6f695df4be54a783fe68ab6ceb005fb985b022f545890271614b7922ba3bedb3aae4e41ae91d0ee187aeb4c47b3f7b7bb36cce5542db36419360c6dd0259ebdfc1d91e86f08e44f19b1e9e5d7c2548aede1599deea3e4e5eff2f418e5bb858b5721e1ca1787e0c05bfcb6089bdd2ffdc8c1a3147fbc6fe8fbbce9b5c6745cb928a5b7032aa7e7051fcfd33bf7e95be64e0af80fbc6dded93181548c6a6f4263f99b3d45e88d1eee074551cc5311f91031ccb5ff15d989db10cbe6b26cd3dbf7fc51b56dad3c1bb98211a6cb1f61e4ba25e161b3e05dce291c25883f8052690c2e173f32cb2f5dfeaa6f19f74bef486b4bab40f7e2cbc3837400dfa9ed882f1e3afdc72ef56ba716afaabdbcda26f35a2487dda29dfe942e81273bd40860f4384e7abc0859b044ac6b17658fca2dca93771879cf56f8368a143aa00352661b9d40299d2e8b032a16313adc548cd959886321d03c7a8f9419e2adcf104ceabaeaedf25017b07a171b25827b292e58b6c9f254b6f7d698073e760792b017a09cbd9bceb4d8abffd560f048b3834580701e1d16bad803a5aa15b0f2195c90fdddc4f45ef75d1ada0dfed37ee41eecdb4145cecf75e6e6477e2769678983762d61c13cbe5097d54e51e745372c6eaee4b494e72d469deb3511a540f48c25c58d059651676372ae9c1470d4d1b3c9e2b7cdf62c4485ed814344ac0b4492167a68d25eac4fb173aaa1028244010f1b6bec7d2852342912cbe35c90cf47202a30b08a6831ad919be330d8e2690ccb1cbc889d25eec2b51a1a86eb2ea775604a0708a2fc97705fbd2116017bae375c28ff6c44ddea36571ea42136250ada9529543a111e14b861442661ba2afab6ccb85518368ae4db8d954d9945e9aeed511ab1b28748adc0f78c43be822fcb21c9a9389a7d8fbaf8d9c124690cf029ff68bcfcdd94e459b3d1486ec3181b64983cae57dc0447b68637d75fa206bd2e7660f669c94709b83b104882441d9899dabf8333f1bd89517c3b0995cd668052844f0c590e3bd2b9a5d6d4809a6acebfec3fcab1d60dc101c93a908fb06bb18135f8a58544eca037fe003a57fc59b726a3163319144af2574ae916abb82b302c5db256e7b99efdc61a46a9f28ae48200b5038044d5f1711de8a89e5c6949b570726d87762135c16a2289bf7bf39fdd6f2fed28d7028237f39592c1c45672c5603b96bf8f6b29766fd805815bae8a75d43eed99b1530325cd2f71610c3e305dc94c4ed26a4bc928128caa2e3a35bc8e8934f26a7d7b8037b0e4abc51d3e8289c8780c8cdb31b3a3407f63daf9896206d18fd87ccd94a82cddfd8cee77fe86c1f1874da35a87ffb80e7433fc6c5fe5d511ee5461e42f6bd9cfb12c8d8a227f113184ccbcc7f085373e71a2cb34ab78934a0becbf6f7875056a125c938051a1ef6806f4b982c38451b8f33d05e0e5cb0c9af9cf85dd0e26fe5dab1d67c4656ccd3288b3b59d6350fb39cf7b895482ad0c36f374b6672047bfa88bd6e7a76f18dcffced6a09740137542e888e17af96874d51cee94d42030c8081a02f6f958a14944d1ce3b3d343b94dd2c715dd8d1f6a7be67fb73350d389950bfd8d2b01bc3ff0b781c9c18466de5f518fd2eac44e06381990e980136d4d122f6da6dfac6b1fa2f6698a1c0e73ee5d8fab4da2cc6e50acd2d4bb7acb10a7dc636ef53692d50ccc7acbb73c88467f7ed5d3806bb651b7268d71dcd76ff28e96a028c57b487e7b4b084344b658e9d319bcfa7a7ed047935b3eda304679cbd8db79c49aecaaf43a12046184de3166e047a9b7a5141ef2f4eb6375cf5856d90c291a01edb41670adb5685a5375de93f93d716eeae9ce15538660c7f6274ef834bf06654d1b15fa97255cf48f813c653301a70332e49f0b4a50d403d3b34711699afe86c77da86b8eeabc38384151bd0b7273e40cf9edef2e8985a25c6af972fc15fc67bacab1ac8d2590ecf4578f4184b41835c3f98cd68a94d4af6e93412b69dbba24b94cb658967e62a04eb5b0bde7cdc40add6972187579f3683bb64dbc6bd19b0389371f8e0c3f460d67a986946091a44b8e601ed4a770032bfea13e8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h15e88c00e7c80ecc2ba4904b68ab6c0ad3414b8ba63c1dce565f0165f63f92c302ae32a7fb7906b2879d73ff2b58623eb00eb44a0ffd91d42846a70ca32d3225641ee9c6ace3709af441a418627fade045df0f4eec146bd18a7e25549e54065d0e027f1d2c2fb67588e307bbc8d5710fe6ca811e972415e528c7bd73fa3596d1fac286455b4d191be171717f4d416ea1254ec1a6d7dc48ab530d320cafbf796571e2876c93306e84dc69de157271d1a3e4142e51acef113db180beadcd1889f79499e4600e603f68dfaff3ca0c1de51e009d833a47b9b5876da749b1a611cf4a0db0e499572c56ed3dbd51a9cfba908bf5c0dd1ff1de155ba544ff697336e554766f610fab6828efdb485efe513bf657d0e073e83817b722b220f91e1f2d9cdaebb5605e28211d3cfe5899e2b37bcd6510aafddcc66c7393060d22dd03ebae055a252f22e71528344c68e667f49090d552da67b69b804ab52f772e32c7842cfe1447fc9e65e141fb632e58af82b066cad715d67bf2f0d55b391c460c279d87f74deaf1ec4a3c6d2afc55f62f52b7fc72d2da2b548fa1c9c06cc546c1593c583f19b59956b0df7846b2d25c2c39a40816f6e6bcdd900b9aca9a38ef80e41176a1c0b28276d7f242bb13f01ee3a8823fb2e34951d1a6739cfe388756fbce533560941366095f404eed4b480647e6d5fc5496511488d8d7ed7cf4d64b1b46e67a8f1e6ec1e71f95f6a76f420823653c4544fbd2eee5c0cc7caa7e4cc9fbe9a678c108589cedbbd17e4b95c6d8c0fea7fe9f8ea67e3befabe1467b18387108a16af8372c150118f2635493c822342b49a9eed533f4f85dd858abd7395d30fcd5d5133d431aaf3cb9299ec21265ffd3f3f40903f6766263c63a9c4270952462b3231e2c2e207fca30a966ffce887abd8d76459c3f6af8e0d58d27e73217e6a6439778361fb1f017f66596db7463c4adf9e4a2051e2df184f456b3b27a62d593c7a907851cc2654dbe585f29fffd87106752caa35fdac12a6fe594e7ca4263a94ee458e812ead3223ec898f9fc578e8167a671168b8bb4e92ebd5d05e36e981247ad800758bcd8d24b1eb808c309480c6ba12c1f91c856a692c06e672293c41dd7d944a1cbc8dd4c0194bae3f8fc87333ba15c6f78dda3dbe7350951b8bca978ce33b38dd568db3eb14c056d6fad291d794d8b7f7d44581fd6f22060b13047a1a5e66090fc6f839278667e25c9466b2e7db46de6ad13779dd6a971f646ffc76e6d3a8f420b223caa32bc39e3060e0091b487251ff3ea40c0accf177a3cf4e98adfc048acc01e8aef41906fef5f875d7342a28b2db7c9817a91507f8a67b445f33cd377cc78e43713921e9d3c2dd6f4eace50f7680ff4bfe7b34d2de7f51f7c2c8423d558424411b86280a924a6b539acc6694f385603297ef8574871873820afeb5c9bd09c54537455bff5df4ba5b9d522d7ed295ee06f02a656d4a9fcf4c36c0e6886fbd7e92764ba5e980cde9fbfc6291ef9a0bb1d438bc066a42a83b140d625218cf66b7fad93d9e2458487cb1fb29e84eee3ccd4ed283eedae3e51cf0d3d33480df2e151d3f0082515b1aea77bdd0a68741d00a723d3b3de227fb9b23d1dec65031006426796780a61092c48ba2aea557c5d21c714a46fe2857e572bdbf917ac3e76abfed426b1dcb5eeb4dc5575eb355a30ba79cef6d76b1242131ffdf661b3bd14af9fca634ee053b558fb1dbe53083d2a948f981cdf1db0f4e64f04afb6c8ba94c8c694e0b24ca83c9d25b517f6059033bc49690562c3012e879f98864d9e1efcf3a4aaa375f9554da46845818eef80a745e8cb875cc0bd0030e8e4add2d5562b0b39dabd104ac771a9fd901219d94513772c1639af50ad139abac3e857e02f0920d2df425a7b5367dfe6c135cc11158601eac96b6dd8338e18541d6082721e19f289972d4ced68d50aa791748692b332a3ada3877281aaed8cc83538fedc581f5df22244e3b779ab37b57c59d485d993bddbd69aa87604ed4d95efdd93c642c79d5d969e5badd44a60b070a2a7e1fa63ab7ab797375003b4e6ecc6dcb74c79526a24e9841ec82d1a0ebc9715d2e42419e3c04f837967b5444f760620394532da802c45f79132b3f459a822f61944f54c33c263f6f155a9da89c9693c86f39e8a795b104cf479790f5bb5ddcb16d29422f8d571914db2b51f892c20260aab4601eddc1ea7bc2bcbd63915c8e748240806e2b5b4087457e88c77231071aa1d422df65a14020289e76bfbd62256f45b2904d659b19922f03ad33f41a70e8c289e6e6db1f1f1dedead4949e62bed072b6849c42b7b06ddce439deb203f384673ee8bf2c43c5a9592bfcd1581496b21ee0547c22c1e62275b75e810d84780672ae29e4c4973dab24a8d7e172fd7adb86ec72748952a3d77f901ac69b820df71fefa7e95c332af74344a571d3246acf6d7020b4b20db0aca52205b70a117b3e15dfecec11fc44f38f482595b3d09d68322b4409a9dd3ea0431e7aeb7b736740ea2ddc438ca20d339d8f391ec1686a650ebf52fd6b1fb322aa9f7f23b30620d70c109c87c3129adaea25a3a70e28150b61e27e296ae74730454d30079d4d5cd5dd3005640981751560fd65c6a5b2c9fcb6a6e7fb8227e1fc19545b8e1a4ba2d6777513105500bcef5d240fca75774184484c263bb81913143335a1ca2240a762b0ec198e954d5ac101e6dfa9ef3de6a9de239f8da77a42d50a4576656c89c403adc21e5da3eaa49849a4cf2ea36aa538803f79cf115ed308a1e7deb5020eb8bdc4a79fe8157d015e10ddcb6bcc41f03f6af52dddd80894f068f68cd924162a41c3d00b028b98d1b409b8726b35a2037db96e42f03b050d47584727ea7380fadbc3058;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h329b73f2a1d27d1334bc47f3322036d59b5be6c2fb57b5b51cafbf90dbf4c32c57a7599db89815633e7350144fcbc210cb85becc26a9015d38ea245e3d0d1481958d4b75dd861cb0ac08ec5a5c4da617b57a874e9786a1dc77d26d8c35698ecc6d2f6ced1f64ad58953727f440a94376a4c62fb5d5eaced4c64343ecca8a7d8c95639cf1a8d3eeba000b161c0882270025e9ea23eeae6184adc24d013adb739a913d35cdc431196bfd9de6f7cc3d8e98810924bf275167a31eb7bcf0753890ae1c0da96141afe810fcbaa184b388a1719c897514cff4dcf49db1579af4ecc524dd3a790945a59ca29f745334c59d9b93dcbc3dfe22ea5d4fdcf386175f24fa0bac29b7c9aaffc52de7eaacad56b36d1a1b7cc387a9b8852826826589da713d99ee4d538ba20733bb021ae99bbc0525b04e0e6f8467a69382ea7ac13378ec08b777f34fa985b5c12e1d031d691de42bbcd7535c92fe873654939ea6fb85e926a4abf52c4d659eb7c5596a8937fcc6a007e18839ae735a3f74e7d0b775191188ede944973cf3660b3248094a3308843a55cb8149cce6c4a84a647934751b0e04c3057422a5fe3390490adafb2a7de1522b8ea7f070200db02d8017fecd2b8e5b17d150b62fb5d9ba5f2447caccbd0d44e06688b057aad2115ce2fb9ffabadc32af72f58645dd71d6c0b781d387c9e57a8c6a9f849a78d125c46a35aacf13aaf86e8e448a5b266c15dfbc1a8721cfb6a91a4572cd0894b64b8c65a21a06a159f1147bcc57aa1c995c220a9c2bbe170560218d15c035107ea62f3afce17a90946c6d38f57797d537e20457224fca3b997fe4c791476bd878f9a6604dcba6846ebe3189322f9699dd6d58760198e3a5b3513344f75b86a39af1580408ff6f53fc1cf2b170d1c3d7b23a5b27d61e07f38bbb15c33255e474fdbb4b59e5ac1e793c48d9f01e678149144ead6d4de0abb0a195e126bea71e42db4e176b5dbae7fcb9130dc6a6f213fa42cab1b666b250b05fc01a6471e5af8314c8fd5de0060839c4d9496321f820d9ac3e73cbbb1dca83247627ca6bfcd1e04c4de783f14fc53259e40050cea9afa2d7c64db7fe5434947a05f71397a35601bd45366d85f067b9bc0680fc77ae186b0eccd24027381190260956ba88131db8ac8da0a680624bdbbbb893d19d6f463c449bcf10e13a3c496b66fc1b6618f990cbde44864adcfe81963ee94b444ca6128f592006f9777803e0e4d7e5d88b4885489074848d24ed93595ca05acbc17487f0b2bb2282c7b5e6c0a1a1e4471b5f5406a5f761bd6fcdc252979437e475643a3be32df72ee859e3c199019730bc352c3a89016f052e87c89604c5eec8a654f133111daf0f95b3d22b0bf3445dd1542dfad902b6ef6f5ea2eed50ab94c16647f072fb88fab99daf1d98429e6f756e8e52b7d618582b250f5d908d42f2c3dca53f80b185d821e03f9a10769730aac6a4f68c3e43725ce58ebd70090964435c823e996b45262082423b07d317769f2074d5b2a95d3a29496f1ba84279b7b011badd8472c2081ee2392926978d6073182e74dec5859566e97d267f0b81c4ad998fd51d3161b28552ad22ae3f0657e91afeaeee20c3e5e913eeae1baa17232b91c2c63f2426dc257104ca202dad092b78fc91faafb0fe49aee52d162f93d2d8522905b51d14e226c7df44c4a932030d5584cc8a624df936c5495ab319e3fe8f465e473af4cad1e49466d5a6b0be873dc810acf5159833a0ffef7b0d72bf1089ed9ba463ee4e86df31ed808abc4443342f234a3f1c77278e22e922afb5f7b73c7ad8a8af0af74c28ab50655047041b106e89975d55e38b5dd05e4e8c22be17d6af4abaf506d0f3b5af9db01d8b5f537be2c6f485a674bea3af0dfe7c9e76af6e4e9774b8cef1e163ca6bee3f671f79b6fdb0ea5130f34df86e84db3a08a5fe5b80fc4e2441b2795190e0533ccadc37ba819a6c4627da53e436ef9a1fd5a19ab5faeb9b027b3926ade718dabf70af350f5d430a8db12cc7df2f3660eb5504fa5b8125f8d2ee5be35a0c930132c5f7921d6364629cef183ed628551cbeae694c2f6f39588e7f4b4fc7b31126477466cd9c866a07f86c43b92f9fe8096cb04ad5dcc78ec0185533976c752fcd95a007415819b03e3bfc40c4ad1e3f7cde922528867f14723241e2d923c97467db7c77eb87ef9e808ee4070042568e55752b8b56131a6ac12c3092e2a4612ea0a573380a544c743dda1b26f7d7707797761dbfa9e39939da935b5d8d65113007bf837baf01472fa52c5affc80343e5698624b71b5bc4c639415bf1ce288ae62a5f9cb3b82a11b42f09b87c0e9e34f98efbf8ece6a5c0dfd0bc8c2d868e0fc1d8edd9d0cd696cc948e919dee13e04d2042f54f110beb3ec7f8645ece0612d0f9f995a3fc01a3357fcad2f6eb6aae4f5b824a1c414de8af877dfa48805b7f0fe84b4b9a5154465500694f653bf9ffe0426158631a0dc7d728e1a97ab7f95c7c6829c555d4ebcbb98db9e390bbee472ed00651888048602d75e046ca987748b62002955c966459d2a7dc8719885541bf163da620b5c4cfdc711636b967890cbdeacd965eb6ab8dc8ad30b74f6224f6760629c9adadc781cd8b2e12521b9151ee62322cfd8eb3a8470765b900cf2f63cb47e06512c1b744cb6f36d227d2523f27da3fa2450e7b8914cd487f1cb40bf7423cf678ac7b198f1bb6ddb6d68407266cb43cea6471578c8019ddc02244dee8d1e1d3b62309ed47b14f3cab17c68e08e7bb1a8918bc62399aed16aba97e3522c850f0b000d5d3c2afeb089b94a8a49920ee3709bac02662db4b28439f49daffc2dbfe8775ce4303c28780b3b66c3b1b956dd95d1778d78da8e01cbe63280bbc42c5d44576;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd7ab451b8f66c4f3592f6afa0b8f17411faf4df9812f1a2fcdfa697f069f517a5628a46ad2428281c6ed3a16cb15389b6f27b79bc4d07d295158389b61afd32f7d12f8c9d99b1d943c6b5f041bc1df0fbf12d97015c67f6f182f7507af053d1f03ea62b83f73a8fa82e25a69ca5ad24ac80d0f28b2c2b49fd186b1fa7c8b6140dafea1c84211c685c6df61e9bbfcadca616811f876d04e6a7cd84cbe93179cf17fe74c411431b2291731fbe8dd1a537f3fe6ed1199766b2b043be47d3db77bd6aa514d1c776e611640fe293e5dd67258914fa9b34e4537127ca3355367cf019690a558781b33bc8268e43514239f3f794c3abb3e7c7e5b0b39a1b16e374e244d3efb1120d6849c9152f4386503b2e766a171c8a931f0c4bd2ad04b7920d3045568d914546f9a3455b32882045152717304d6dd2b133d90d325fd3b4deab3a54dec7dff3eff5b19df0f0e3e2d852d8b2d5d6c73694739a6e7beff3ddca62e535db410f5300b6919f95ffb71bcf0e8fcc8e18f9e2a2260e7aa3458bd1e48c9f459d8ea6c62169c872de99a5a5e566f87bf43a6a9ba8bdf00f2ec42392af8a06fc49c483abb6e5b56cc6e39cbb33c886589a1bc5241df6b930da62d574a19b29ddfbe5d72a082834e78a3718447525cb91f0b693665b9f73ec02eb76ca021911f582af7712ed9eb6bbeed84209bbdc4105b19d15c27824353c00fc5736151e449b8624860fbd37645c8f1cb267c764edf1f490dd724b9968c84a7dbf153f874a5f707aefa8e4f5493f90ddadec44b03012c1daed4de702f12ed2bd79b524818b97245217d9c550f4ab1791139af585cbbfee54e3deae09b8bb131c511f8c34853ad7b54f093816447081ce846d9381a560df6fa587d61e5c0040ce513b4ed6cf6321f11deab5ce3babaccdc474ec0aef9de298a2b8c4cc177d16c8219bebabcdbda2f7636f0c97da24a71124c4cccfb0e23d1dd7dd5e40b06c25611c9d78a708b1ad85a621a1a8d0ba8f7f1f4498c2e5b3664d3a08018de2402851c57be541d959ebdf38ac5b9ee3b3677acd173243dac8eff081cd0f9e2593cfaecd15e8d8c68e4db0e0fc6cfea7002c06f2f2b71f64a17bb6babdc88c4e606276adec7357ae7f09828402fe85ad76d5e2fa5df12a19aaf10553a823b85ad14062962c28d46586c0266ea2a9594f9a870a797a55b9aec6186c0e354ad143ee08118f07c449fcc6060dc53cfeb27ec5ed0703ec17023629250f16de3bc174c8d093bd3fd9e23fd0db973044943765bfa3ebc6f6dd82a999f899345fd68fb1b72e6538fe2898e0996494c006f77269b3b89dbc216ab6bccd1d8228a15ce161c1d5aa8893aa58443c03c15fa2221a0c6fb8066dfeccb601df499c552c12484a813d0f4f2e0ece4b05e124dfb7ff32134ee517be8d95af22cc906ad1aaca895d551cf9aeaf1645d54f020ff8fa9a23000af158ff3503193bdb1edde0c1b195857145550d8cca3b4d987d74c9e0c9061cd17b3b24a4d0443237b61e4a849695e961e8a205fafd401b8d09b60e241f7be710188bd57cbbe7e0e61f71cb10520190a08fd7fc5202958f0cf4d4da9eba2a27847f0033f16d2b37947de57565934006e6eca371367f50dc1c6e8b327d50eef32ecc599bfe82aee1d74618a0f83affcdf33f633885615c8fa2358ebdcf4c3be83bb06f8a08a82b2af3f2bdbd790bb279d3a821590e7b217fb4060594bb434bd3db1efb8e3f57f1cd57341af32e07261cff1fb578a86736114cf363b67da4af89fc4a063516bc03689737843ddcd5679da1eac5471e6b08dcf2f8da4af346be42ca76ed7ecdb9b4fd4f775f66589f35e993f0018edcd14d52264358bbcb435730876f53a8c19f9d6046abd234c543f43185f6fa24a0b76a1ed6551f2eb7cb333d3db1be859133cf57424ce70fcfff6d50b4d2fdd9e1c698f2c16a53684f1b6c21f53a6d08e3a4bd66f7ebaf5b5b0ef491926f79c69953f158e96ad3001ed00c4b554fa9fd6e8f6838eea181a812a976bddee69413a3460bbcb3830154d18ca9d3ae359a32cf53bf798e3a6b59b1933b435cd8c8b41fbad4afcb620233a4880bca62bd1dac09ea54c401f85938cc7dd00fea2244c07c0205570ddb3596381e94f82c75b16c56c87da6a38da8b20c88bd65f7af18dbacf27eb9a2ed1008393834692f22e230ac0f725a919e08cf9c55d5f74c5561cfedf5b3d31a92f2f3cc438c67b2703d58acc2ba8ee6f23e652bcd56affde3721d674c8f6ff2674e215c550a7654b2fd8c3eb40f70325b8c1c7778eeb098e7ae1cea819a881ee3eec8cbe5a956949210d698430e95581138f9bc8200039ec66768276053995af3ee4333d6d541a532f128a01d361cc05a71d080ce1cc1f4ce5fc65748cf36233fde4f6207659e9cc4af52966c8acdadf684646803fe7e820d0179f783cdf612b2ed29722f14a5e2ced5b7295dccb5b900d89304cd827f83475e17af0e4bf2400bf8834bc0d66ac68234d4cd508b6e8410cea192c48296c0bad1fc91ee6a3812c04b8a8dc268fb4a961257a1f864c1f036172a9f40f700934163a0fc5ee4a295a0910bfacf68cdac2253a56217eec9da8dfb9c426bce1b06aa5d29d2e538038481d8a4303f2d67e86755af658b200c4f7690479cba1180a51d3489f988222318d7ce14c3a0c66e1440184ac9a88724406ee7fa4593d70afafe7e00bc70f035b2cc9dfbca7d5e2c0997f27c153d1cbda12efcd1cd35fa10db3018d20340d6ecbf9de80df84f79f989eb64d1f543379980c6e80ef7f8975deabb33de54de22b58b4c3f096e7a575bfb5af57349bbb4e4a3b29db6df9e92ad78e578d0e3fd331ff37e9942a0e4cf979638124a0715055ca59e7b285b51e5b62369c113fa96dec387b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h74ae1764612a8f200d488b40cffb1705fcfb8feb2ec786630e9dad7d60a02d5a18d869375f9e2a54d33ad884a0b893625326761bec2d737a676a04a3311a430cb2d0a76c1e974a4aaf9c6c0dc464dd90f79052e0f64af6e7936e3d5beffd38017a19deab9138d50efabb435fc394ef5505dff8fe9ae6fe774d21e79589145a6c9f3b509160f98fe1f75665be5a3654a5f5fe22c3382f1fbb5b37882ce1233be3f585374eab0c3f4a9bb233bc6c4372ca105e0ed10e95df652ca646edec136d057a99acb317f9e9af1c3b72f19676cf092bd7a11f0e6115faae42dfc51448436742586667101e1c2a5034a58c01cf54e3e7d667d042c5c2595496ce9b2eceb77f2ac20a0cf65213987bdca8a07fa81865405f9786dea6141bec2ea24d549aa5ec8a038f579ca52ecb8447419d374136eefcede23a8b84f54a549d4be1f23b97daa5d7e993e90de9a717be87ddfe55c00e217112bd457556fc382979db6641aec5001dad02a97bef767058e415163767c6bd53479a054017332841a1a0a58612fb07334a40263c2bb143e29acd29242389e445e0acce68b7b055f7ce61975909ca4c1cd47df2f73067651758348ba5a3612c67f8ba08b5b0c46d1b6a06e8719b08ea36f15ba9719dc729f1991b746bc8850e8f84780226dd82727fe5e909cb885957d49caa5d0863c09370b9dc1668ed190b580db6713b78b7d4ee97abd51e69475715fb15dce1aaabb1482fd2e7b50543fb78d255b755d8a8df8b7816994fda1cdb5b45c338704ae05f7339468d42d481aa5e6aed27d2f5f66d0ac8111360313837e544624aff34227adb2d1bde2bddb60553a10a48b38966a2fbe62bb5088e3863b55bef3522c09f11c81cdf703b69f72d9fa44f83b76d6129eea491aca0469bed2ebd6915346bb8d19cdcbafbf71bed24a5552a8302656c620568bff4fc222a4640f5d6ac2960dbef847a61d59233882fca7bf1bef1f8043abfe60817e2e7a684ce33515a9d089246801107c35a8e409afbadfe29840345deaf5ee53c57e5c17fc279f7a5cfeba0cec17552fd17dbf7b2417a004f67936501a679e401aebd5491fa21ecb3b3da0a110869551082db082df59294c1ba1f9173de6feb7757fbdffb91d9f1781fae22e2326b87c57abb19cbbd5a6f2ed33937ff5c82aeace6c6570efc1505521a7a4e09659cc74ebd7c9f5bb1832fc4fd5150fcbcbc6f5c33afadfa5d288e50d04ea22323354b2e3983ffa1bde2f13b07c88c4b4687442cd30b64271307ece5fa123b9170897c9915566364a25a120cbe9d2f481cb590a3054a99966c4bc478d3f238c061553d899d4ae96c5be03bfebf2aeccb7983391a92150b0f851c85d85b67cfae305c2728161d95885f1158e625af5e4452a057dbbed56c1fec8cc830165bbf20b642e3ba6f0ba47ec70ecd4fc76af20c8840cd8c6b0d83b849d3636663c9df6df0dda69186076459455c7d92e1ffb9585f87463a16da0cf5032244d1a371dcafabb44a0e45c73ae9ed638d66636a6bcbf51ccf98c5818f8652f1911fbcfd43e9596860405dfe4d36f22a506bd8fa7e6b42934cc9b59ffbbe36d51c31e944115a872fad9d73a02b02f2ca22808b333cf644844b4ccf651224b8f541f285fe07297959725ca4cd7c60aed62d68f7522515b4e4a74ab83ca5853e13a30f4ffe0607688d4a4cb199c7e2a7f54709a52930d72f7513863dbec222924d8f83552b1ad0c4288e28b2e478b32f4e6592a2db58e6049be631c8d50bcfc992afade20ae36746e15f300dafc8159249d29ada11aefa6383e715e1a19c8f63db786c0c2a38cd498472b33786e5f58f9aca1a07f52dd262b737ad85561ad0e119d80896814bb0fa43b01deca49c685b89af90c0e9f4bbeb41f9ce78d0137c423634b51cb528a44d8c8a4a7f7d509f6ca90b9040d2740d844fe46c2e49782d2311805d0a19b8f8a0b0ec8c87b98cd1f7dd0c9d446b064ab0509f71922e7def668ce53040d5ce09ab2da60957c74d3a867b6b2cbc4eb58aa4a8c74dd4dd4468e6b1d2084ddbbfe269d8cc57a3c59a0ee6ae7f5bc16bd50d06ac4a1f30b83523a301d90a073d918f8261f3a3cf682304a2d886cf79a6384461c7f5acef89f564ff0fdf9c0a7e682f6305ca018494e69080c9c25f290f486aff2f48fef6ab85164ee1eafcaf10907d2ad1d45575c42cc422ed1531af57f389c31897f94574e93ec8276107d1072b23b9977cc387c111e6930b793aab6b3f09323517350eb94b83c5dc35e53d100efeb3b5c52db22432929f10d9b2e82be877f04e01aa64471eaa85aceb90ca1eccfba09f5a4f980ec5f29220d602e847f63f65e7c131879222076757253fb0c1526ff923f81190c147c5217d0c5744b9972e36bc23cc47e235fc3b58ab89e1c0e1a3475f2f53ce1d0fe867febed62713e19a68b6e082d55d05d3b8d21b467fcd010a4fbd7406a026abf46de3554480fcd0119db0b1f6b4df10bc7c6a2b6e7f4cecc50ca316a69cccd2a9a69717f1a479c8b9dfb95a0342326ce4ac12e06a427b8baa0c359d3c327115d9bbf40d963bb72ef963d43557642157855db3d2fad95319da5bf3b2555d3c74731683fa2b6d54202883b656d262fdf260ae736d1fafcf836f03a415291f239a963a15771915b9b71945323366fbef16fa842153adfe90aa5db405f407dad6be72bee71e702646406bb57fb9b42e7130f8465cd4fa505c68c3249f893bb856b38e47e124ff697020d2f955b9262001d02754b772dbcbecfb7fdcd70f2f43077d2c341794e1d7a0f7ceeadb12a0f6505f25f2fba12970b7dbe2dde00e5412fa1ea6dc6ff1759d40785c06888a0c6bf452f3c1f75908d247925afe6e60de9939d2bd36ad15df5621d7925209a12cb1fda7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3b725099f60db12a6ff3fd0b9872027a1ec7d40461c40f92f447e2c2418d0a64f7063b20df514b18c192f43d9e7a2b6f800e6f4f64ed78b3d5cbff3b03b1934e1ce41d673f65c4de08eddf8ec379f50cd4099f71aa58425a164106c2db0e448b4391c639741c047652af2bd8107aae8e68d7f0a6e88b9c7006cd9061a191a2f37c7c6d60202b5d1f0445def10bb51291e8a34821a5f2324c4c710e3a551986e69f3f765eef1675892be9cf1434b3b8a82cd7718199f1611ae86d9fd133a9faf487b18c0feb30f20bebd79ea15acbca2363dc8fde95a69b613833e695fdd2e33130a284ee228296795c4dca2ec9531c3938f0c7b8ea783c6622685d673a8de7ef4681b19c4392aa14626f4811cde87aa142adfe187fa4e55706a6fc39ce4769aa986dbd6ade6ae014c90dfa43b89ba20c16f134c743bae19e9dc040b77d3bf93f25e22a6078273544e640144874b299acb5870dfbdaafb770a221e3754c33d4ce914043565e6154db3d508b1790720857237c9eae17a1f1fcb08b929fd0a5a1167f68ca9b84ed8729e3f9631c124a0a738827f1bcb19f3b2443ab54d410b0af59a4e978f67fc598892e8906e7af40001d28a7e5e92c04e1089b33fe782fa582643c4670b79fddce20dc6bcabc8dc74a4e7d191c2b3790ecb3b216ecfdf7ad85a6018b8033233e35f4f4bb6e393c94710b33ea0f79c38a23a42d1433647e13209c7d47f19ebac6d90cc138f6a0e62be501f3a9b1970a5132407671f77fc4c9b0cc41a5a4726f2eaeeb0742a4d0a9ed8a646932492479fbef4e04de35ba2b0d9f42b75b02c73bf65c0ee1fe271594380d7f389279ed69f7c9b54a1989fa15f747f90b34acd458db1a3cb08cdf3f8a517c6263fa569f16f8461187fad15dbcaf0a410fffc31699579ee2990e77052264eaafa49754e2f0fbd156a44132cb50fb4224d6572065057a615a779f1b49c29a038bf048a6aab09e46cc91a2a4a905e085fd9076c4581fcbf71d5aa4ea1f5d85509be07e4573e4cce313efe2ab3a1c5b8af55327d2787bef83084cbda0d11516894b4685000353a98c8c03cb8f9ab4ef2469204fab0c0122fb13a616a2745340d703dad13ecc29ef0718ea0a510e68020e7f7993350389b20993c86117a754d0f93ffa54047e779f085e2189cf49abc4ca60192831e2938e7fe948385a6e5951c34a6f7162133feaa69894ae7e79e04e70772b1cb2538df672553aac15e4b7c5823a1ab8fdd75a560dc4b631a9bec6dd8857ac73d9d016c7a39a9fffc98cf4c90ed5e157a3e6f3b06552746b6f4df2abd3f8e09265a95ce705c0ced8612b3e85c0fede115c2805dd22d5f3bc87dfa7436fd85bc353ae83d88c0cfdcf121b49ef3fff77fa4bcf1c25c4da1663eb6e4d3b9e3d2c580d2ceda0055398b18d438616f9c6cb6d57c2138b50082af6bc7baba4300828756ace6f3744ca9293d0c1eefbd4e5267cb2b0cdbd288edd64386160b7213fbfd094ffb02f976816745212ffaa3132354cc3cd04c29c11bf49b3f1175ca62a1b4088e0c7ddae9997ded3a12fdffc89b949c4c943a3265fbb02197e6466af77278f8af74b5a84ab90031942e26cc4dee141978280723b4a43fe1ac00514b2177482ba08830042a0ed095e017d1e6db869a75cebb5b804c33d761926eb214a1d47fbfd16415107600ad55143995d373fbdf0b5cbc34c577ba8e7db1fcbc63ad359c16a9b877443682d265ea988eff2d6b4f09d0475f37625fe576bd34df5210521bcde372eafe867cb6188061442b4335147804cdc557ea3d95df412205683c0594670244b631a17e78bff929ac13e1517aba55fbd355612be39337d5f7c89441b71d4924fc005f88b2119f3552a68ee2f9c42ea7c3462b26dccb0b94a6f0804003dd2fd857a7d99ce684cf20caf75e66d5ffd03a56f485b29cc69565ef93f7b78080051b97cbd2a300e9ae030d13925e7185a83ca736451d2fb995f041ce4c5f40a0994b79f32de2cef3da6b57c0d085a0de14ac2f9bf45f0c3070e4880c8fd7ff7fcb259ee9b758f12085132adf8749ff2418ee119be15aeb091ac5da29babfb9cfe53f7504ba7fc494586fc8b8021d19da1c0d7f2aa931c5ca8fead11c7023421b46402f53f1d19aa98f3d767ae7b1c6ead4a19bbfc36bdbbaa5413660a0016d183268f92ff3bc0efef4b613c8c113476e2b74bc9552e1d70ea29cc2e4a33856e85684119150f8a9b9eac5ef0f703f1e285f6081bf63de129ce596c216521a9f53e93dddc51fa83e871e1d9f3f31f1fe33ad536abd870aef39feccb22f9559896f026d99ea151ad12ffd84170391a3f8dc1392fdc505ef72defc5fb99b50df8fbfa7cdce601d91dae64efa83346384feead06c568e4ff42af1a6bdb30c66ee9d459e0cd144ff737ba6e8d85f996f5276c29a0d3a388db1c81f018a0df689eaee7f224d6bab76aa2e27cbf46927bff7e91e39faeb1fa9b80c1ffe9bedc9ae27eac9e1976714b23a6118805bb2f39bcb663b38174b1f84eda66019cd6b4673a79be881a2d97e469d370de7525109c6b9ead289c1d87b01aceaff24532d9906f561e2cd881ef280eee23ca9795cfab59f946ad6df340a4738a7ca77717d79a206dcbf81bedacbaef034fa7cbd33f0dec59895ad19ae9aab8955bd7e69ecfef289dd51be74318b494ec4a3e5e7e513f3949fb95f4f3d1c5032389ca187b8a7d799e45105bacdca59ae446473b04f31fea013ebd4170586e6e174c969b546e2ce5ce9df6a8499c326e612ff6030db905ffe5971ff627a2e565949cedf2376ca687a7c5331e27355298d680ec4fa31d639464c26dc1f679370badbdd7c7e5e52955dd5fe6d06be57d3de5c4164a70a51a77df4c0cbb127e7d5691bf7064db81f762;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbbcf32f8e70b70116e96694c083c4af31ae5ba73a32e18ca6998fd4ca4ccc8266d297d7b54657733425bf2a8d030bccf6649a503cf0a0c3ed51c917abb2c6fd39a1ddaa2c556cd9005f1fb420ee40b3c86a15265daf7715810f30b6cc0bc6f3777200fe3666fc7a2288fba0f25cf9f82b2b32da180528296212be97ac0aee70e7728dbf8378c00cbcd985588e47e7df4e5471ffee964601554c6740b318846a000d444563d33d70bd9a26a4f3f6628cdb55f39492fe264da89afad3ab5cdbd16469c8efa8ec255f694263f7b517a872de5fcd929b502fedb35d81184d0ac35fa90a171b65c7f95bb7e98350190c7eb10cde8377c60713d71e650abe9653a50cbada801dee30bbaa8a1b1e6f5c402de3f7c622aa4a300a466295e481834594143a7fbf71f136f63dffdce095ee5c4decd71d8d9305cd8143c0fd16b8590dcd2937292c6a2668bd6257aefe184584eb7d1e2bf10bc03eea7281d8d969e01ebcc92d256673f12c64a86c09c21eba511b852b9373f76002431e2ecc042ec374dac871f69bf320b2d354d00676a43fb22ad5f5c60150c4ea1e5a914e819e0d0f705f9685cbdd55824d40ed2366dd81483e6d8ec7a0b9bc6a10506862e7e20f726a444c32fe0189f9550c1766331ba50e9540653364630a182b46630d1d5a71f4aabe2d4d648e5e03d7d8c5decc265a085d7f5d19e7406b5a09fc8b29c0cf66fe9e5e42eacdcb2e58b69958918a88304ad688470ddd2c07468a06d7ea34508abafea3268ed811573e784918b1237237854302754feef75f489227c888a2d8df0fd743abd760456f4d43351ddfa763b1f880b1238cb5ceee3e59aa448bb979bbea32dd2390c95b32706dd4a64856ee0e950fba6e783bbfbb079588bcc5da33c9dd93914a5fd8a6227d58c872cf266e7e43a6148f95f158b9f726549e721aa2f389bf6a02dd932cbfebf1cbe90420a7b3c331bf8ec657401b62415220d93eecaf226af3f1864a2aef8522f86dd85a6dc29d7f2ff38bfe18f89a4bc1861033eb89984d03f9b689f0d80a49655c5da0fd9150a6485ac108d588e7b5d16055bb680c12425a32daa040f141c3932a29036f51933c25008bae7c215a06d632e6aef56d47590f55744958abdfc6793122edf31525717774cc0fa49423e016a5707e19f3220caeadd1b22f2867cb5d0dc08c94a19e4c25bab854b7fe70979ace68b5e7364827b85645aa9d5f4ac886bb4d97832e60fff8e30f41c4b5e726af3fb29b749b3e298384f4785f4d8f4c17a98c12ec0445ad9270ad35eb3494dbc95002fe2a466d12c695387ed0d84f05f311d93980d7184c1b532b026152a4bc6f5954689d636d47aaf505b56a56a06f4affa23f29105bae611ae869def9dbf0123978fd8a360c579b3f85964708dbe5a6b73a588d80b7af8ca85f3fe2c0f685f03a909e55b477e142f43660b9b9979a167fc5140fe3f3fff54e3de1677e3d690457bbbe04d8a2b5daca75da2de183c01ba24c7397fa1727d071736c90021b37849b2f47a280d0693cb562f45359e3444dcf6f4d2eee1d3eec4d66cc819333e11ac769ba887121d681ae27e04887d702caf462ca8e04226f291f5d6d919631eff975507aa06e081ccbba09f327cfa2cc73bbc0f0f8f95338f3363a6f2d5bc28cdf2d94f81ef49866eaf4ac20edd2b8a89c8776d9f0b3d1f7398ab8083159acf36e66f92592fabbb1e21381e333c30b51e60fbfb611dce96b0e842f39a7c272fe2b48bcf7630ccaa3e32e0357c8921a5b75b6ef6f86107c85947cfb8ba81a96214d71eda01fdb9fa969840f3562e305198336016ba4f517846f5994965c58a8ea37d150f7571e9e7115c39739441ba4fa0aa2704cc517c4dc1c303476887f5e9b8b822b48750cb600316e8f0475dcf513f4222385434e2964c4d58bebd469316abdc1d697242cbdc2253ebef2eb645628784be6773cd3292fa85d4d157129984cfc205de71c70f9028344f6dc5fdaadb8c0bfafd450a5b5d4369bb1c24f933e6bb25982c0615d50a1909f058b470d47d80fc8785c9336e69c03decbc8c5c69a1dcec342fe4f908776b620b5009da84d216a0a55d7f849cca5601ed9c87a505518816c682bdbccc38298b5224ae4ce0a8f70065da93df18d818946c82c2ef39f3e08b0d80b44e9bd491e045c65c5357d25e47bc6b7d3329fb6d428e66896edfe9d716a454841ac44e5bf63b30748a758c5a0aef81f718909dfcbc3e183850d256574fd826e4ab3a9acd37fead4ccb3942998e116dd0daa37b678cdcc75934322cd6cd56102d5e225e12df6af000d2aaada01cd1239fad4f4ff0f2e8bb6fa63b8c13d0ab00fa1c289f60d039ff52b72abd5197800e8ba0bcca084e9c1d1df23fdd47bfdfc309f28ae2901035c2ada5d1ba878ea5a4264c336b8b797f21487129ee6541e45c3838440adc9af452233d6fc1c49203a9b025a73e33baeff8581eee18b9b91383cb5b1a7dcb02bc2f94a8bfd10f5e84e7eeb3107724785d2a6decf35f133b361c9f3d9f481f7679c8000c30489afd71f25e63b0dddf28718232952ea31cdacecf5246b58befe8143614e8b0ea451379d90a4670e351daa4e9ed483c49b83a962be7775dec7577b66d9110bc3284fff1344c7bac2f098d8a0f5e94bbdc4a51534f331da63bdda37541c40f34adda819c39dc709c72d22359dd0634c9a229bcef0b2b0c2c7ce7f2075687e94f5bb1128d542f7baebcc58351c51eba336c6dce42eb59a754ef83845bac88fdf369a44da98fcc3cfa31e668d3a9f20d701b74d63cd7ab10bb39bffcb353303d1b76a2203b7d3a8e23a0c9321f2286bec96eb7c1bff69ae30ceb9db9063ae630ac2c5c0a84ba75bd44aef1229ac09f33253feca555d6ac2415adc842;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbb5acbd7511b789a99cc9b1d3f5a52ee483743d2b273dcf1d28fba73ade2cc60114f8aca39d75b0dc073b1a4e924a74b9f536ffc3755fc50154c58d0cd31735b11ce6f92cb8390507c2a42b06d4a28f11f4c6160092712293b05bfb607b3670b40ebd57bcdcd4858ea89aa094e71d516963b3aaa2fd84f50bfb7f883bf4300736cb551a5d106f6629c2f811d2bb53a0fe6f0bd32c3704c607bc9586e3987895219f72fbc892481ab9bcd1223c24be71150191ece3cf7c5b7cfa8bdeec3502d0265432896e0d7dc8aa01db4515268cff136a7340e06618e7bebd432dfc93c419575bd2a195583bbd922110c37407d97b71ca0f12a43e194bae4c9b7caaa44b637fe58aeaf3ef826cfe747a13fed83721337584388889be179e8483025c19eeb39e92662522c269860dbd0e7173708a85450c09c3b8b9731dff7e60ea05c6b65f76458c44d34d46d01688da03e518f6061eec56ac44388d841766d248146d2941fe43c2c529dc002667692e03416ceec2260746f754d3ce5875a248d1bebd5bff5cc8031f2033bd3e2ce277ba2584f6067f374e761bb3fb3644277940181c8cd836c8b2b7d3c79ea51e2159c7abc9cae09aca3581a7adaa35f92d2972e703a7cd92cb10e01d58d473e10bd7be38c4ba39c5a2b2e260fc18cb50f6882fd62387e9066d74dd2dcfdecf4547ed2547dd3d53fdae345fb71fc3532a193ee41c84fd39070201b5d4338cd5ec36661d62854e4e13857b08ef93f31330645aa9595d62e331fbb2911022fcdcdc67f64d783f7ead1bb9caa9be006d39a742c685756a49cc14278d4e38467c18b2a60300e085e6bc412a00d69aabad368f0f65cf42bf32914324fd62b12244da9195d02fc81d72cb448bbf92ef8c8f157fe458a703bacded0cfd8a4c3308e031dc1999010c9a91832fbc40c9b69d24e3ffad7d9c48d78aebcbc4af2acb821396d2031fa0ec3466c73973129a1290eaeccedd84be1946a69b45e6c9998343b89b105a6b494cdbdb88a268b7f4fa26b7f0441d843c7d37ee7abea883c0db4fa2b575977f7079059f4d388e0c426d6942db94f15b50c7730883ce72d8e20077dfcf0e72a0c9f62cbdf58bb5a918202cc9a37d1ea8897d3708ea0027b5ee03c750c331edef3adb9d5611760359385b0122f7bff1b8e3ecc2e86e84e4d991d87cc3b230a92e9cd965a41d6f069b7e3c03cf751d182bb97cae405310636870d6efbfc7e3fb1086415279e62a7223a300152a1c03ae19e090cd305d675285b5ebca5c97d7a10ff72e5206e15279cbdf4b7876c26c9819dcaaccce47da385a0db75a1a786845f5cc57c79398ea9dc2517242117113a4a71916d47a93f03107bab1e94971f756ef95573038600720044bfe7cfbecc177283c47e54f84d5c952f1b1d3c4c83b66fbd4e3e104f95d486ba26699c0edb2e281934eb5b76c18bb47dd21432bfc711d724b0668cc875d1e4a65181d1266e0bd42c25a684fccdd78a73267801c4f21a4865cfcf279592dbb108b3bb5d2bff5318a9c08163c1307013caf7010abec27bce6966151dd45475716e524ed63b2d8679b18552204f02d73052c50c5b3e9beaa7b8307a6cb9de4005637bdcdae21bac218c21bccc238d3ddae90771ed710fd6a368d2165a0bf80aa1dacb1ca71515715e396dab97e125f92df498d89da3c04f72bbfa728c3e8d7491e0e2b52bf5827177fff5bcc6b1ade3eb4ae3e6cb4cc5396336b88020533856a1d2a097c3e11f539653bdf69b57bb9ca408846d26fcec5040857ee0806e1b15ea8a988744a8ac6f8c3a4d08ad741e0fef0c42a6fd6f98756bc9e8f3f6d180445bb98bee804118c3003d53f7d55c24ca2210fbc34fb449ef1d6f81fb7ae9294081cd7dee67028e67e29276684957eba5eb839cef7248b4c157c2bc5cf043590ee41b8422af95358750ab39a1e27de514dd1763b35df77afa526b202a19a676f02ffd27dc3e75b28f3f228bb898ea9125313beb9a722cec6a16f1bcb6407d46ce99447283280915bc3b6a24d3e8482db298f8ec13efe55859809f005e5942804f2d0ecc3500ecbb4324722e3bedb9962a0c99125f63d92c4f2ea08fa6da6e074c648d7335196af1b7deebf866750260fbf13bb7f13cbe8fec19b5ff7ad7e6d592754ee7075675f3fee47de2b6869a4f81b5b16506d2163acd63a778bd0843341e42b522d4f4c5dd8b289833584ff2594fbf80fc133428b43a35f51e97289fedc28f4181f14e20d32505c593135d2ccf12a1d52beb15f42d54597e10921c04e7cd27497b9a372a9d58ad8d169ca235caec0d84621323fa2e34f1467d6ebaabdf17da0c78da1a35e3e07ce1cf7e4a0ce4b17b4aa495455f6be5ca11e89914a00b0349765a96fb62b60e17a9407d5d573237a972c107969d2133003ec320fb39a88039b4e5d172964df9fe374de1cbb714e2c91ad7b4b4a1a2567cbefbdaf08fd72675a3f792a0bd01da03b113408ada7e456f22d993c49a44c9e1e5d6d56507409e0ce9d8892018c76529bc746d3bdb371be5a94cbd951e7fd87f829c63ea9119fa6cb1a811fd7630ff681e0532e6ba77fcf3a9c64064924706f1ed3efcb29cd3177e9e63ed31fdf8d75d6d29fe788bd45f578fd520ec1ae2b14877649c534823aa62dbca2f36d819d37ca5487749b5773a0c4ee3f32c6705473ad8f89cc60a80316b61731320c9ae49f90517550a5aac2df3bbd3439df069611d435b3365db9fcb51942920346ccfcc589c0ae6a9c16223785a9dad406b619946671c48fbc2bd35a10ed1dfc6cdc7f19e60602dde783ccadcc507f515682d084509c25fb2d308b5ddad3d3bf717790f0abbc8e8ccc8694f2910850585d9c128dd98cb02f685ba7ecf0e0c1efb7ccd463538753fcba6f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h80f98a71fcfc5ccc6694038dc0393354eebd8024e718f46242b5f17cc230f535eb65d56c2dc49726c6ba1868e7d40b08edacbbd6a9f92a240914c89e2c8320e0fea2e4b929e5ee6d0f047075915bc1dd7b5b2e8ad4bbffb144af8bddee7b82a8e77421c8c4156a88ee4aaad748c6ffc0f7b958b0620bfded77667fd70e35a2bbcd2fb0874e0020608beb2b4f4494b1e036c1eb4a2e58dfb48b0402dedf0587d1c5787c1c3600b8bcc9b626a44a2cd6cbf9e473d1ea07ce135b859707dc74a01cc9f3168c2d11d147fd714ccb24b929d4511e0df2d24604636f6a0908217ed20d895718ca5c93d668c42b66e3cc119b61969e0f349ffd0007f718683045c1b80abf78751582a1ceb7637045f134d9bbea90071425cf31b2984066172b779054cca7f85fb1f74d4dde3c67286f275dac99d912770d4cc066c910ff394e9e0040cbc105b7c7a817943bc6c2d699b0a5181ca78a7c6254e0e0468e2df9a0893470f29205f528c0f5496bfeb04369c17407a6a735bc2631670faec32cefa5f602e8a1ff16b8832c47442696548ba36aeb0c4a31e7a04269a053af6d3ff1f594a91544735cbd7a6bead347322864adfd7cc8a93bc1e2b5090558f45b1507283cb5d87670f8f6195172bb620ad018969cb7ea83c13f7541274ab59b59d4de46f7c4c9140f22f13c075b6105b770cb18f8627d60b5dc73b93b0566add0436192ea0e2cdbe9ae70a31f3ecaf61ac43015a50d6284fc8f6fe93700214db00efd53d14e8787ab217e3f7b6ede250210df6dc0bb57ae63dad30569276f763658995d8eaab080da718ae796f3fbe68b1b276dc2f50baa3e27c4433eda4ed695ea6cf1417b80e2ee458c37a42dba29e21c3f8f7fe8b620009ef3eb5e13691c2252db7a478ff485132ef12be33552b4924a16c676d2fe99d40d55b90e619a22d2f37f8d7a7c266e9cfb03fcb2d5f1fb17e4505dd1d2b5974b8d6488cd702d8dbc925d756abb403e14f72cb363a7053d7c3fedb1feb34b6e7ce06ed191563330ac3899fd4cde5cb4c77ce861bfb757780a4e64aa62ca395d221ddf5dd79464d9e5c31558f7968c8636b0df1f6a88f3e20dea06029fea8699512d579ea36d4664fa903a600cc7b8c725dcf743294f9322010e26318fc1e215d01f186375ab32e85aa20b2f08624201152fcd53c3e5191d319b3c2b9606ebaf2e4a0bbfc37ba48c7f63715634bcf6bc645617a885f3fb0ffdca66b9d5477f897241ff267218ee7ef7feac376f717e6c93a4767da3bcd8d6ac0cf43be208a64cf810472ebb71f1d9ccc575f718d3474ada2772504ca745ac522831f3eb3ec57dfac749bdfc921208fdf20fd33880e018d81eefe1a7c68ad0069f083f084af67a60e05c55711ae3d0276632779f60394a02a942047c49e6619c43255d1f1f3b616ea0d5c1e071ada9f92394460d3dfe94b9047f2c12e1bcb3be202af690a87c75a583def27f5de225588bd7a80bf7c836dc048b674f6d784a96e0c4e6dcc39762386ad02502635c67be17ad4d119bbe739f6be0a0d34612a540a9c32c2acf0bdd52db40789e3266457e9af10f023dd632eefaf3bb0ae1c3ed6a958086aa5ab9774d7490fed44770443c335b6d4fac521abb767c08b3a6d27ba1b6eedca0686f673acfc36a3b2f3156739d677e14c1c24dab145ae35cf1470c11fad589a5c9d6718461d8952f15460fbbac3caf02c3ef8e8f0c7ae92a728d9cae45417f48bfdff04537ab546f196e851ff7dc4641f83a60a9d08d3e41fd0271db24fa0d4b3969f22e6d54f68869c3d75e7d3d88fb4aca79fd78ff9ad8198ddf6fad60dd7c3b5724b921cc6ea6aaa0223c19f570bd037d3b61faeb44eb2ee14523553594cbcb05a1c9fe962816a4a22cf597505f3f3466f6999ca7083dbefe323c9723e568af31e452e0d5f294c9f3bf4020ca3ad78fb3228e06c81f17b1ff8d6487c8621c32809901ba8c61ce6093f89d8fddf72861c545e65089af62df5f8be9da09b7d02feb1df1c1e36682582e4d0e2b57befb779cf8347a29885e9c019609dab72c3f3ceb599f4a3e646552619f3c5005f8a9f7e867d850f0f6f96f3ce1a729547e30879a8d224467a5f1f098e896783a17398f40b7794539b42cdb17640acde9586c5222c89d280b0aab6de04696248e89b700817dd26014798a40dfac15e0c4c006a220defff5476c69d26877d94fa1bc81e7f620cf1af9266c55e2e37dd9c062fb207abd381daaee5f61e3a94bda1df151b5fdd5a6e39e45865ed9bada9e80da923cde2e650b36b681bf8fbabfef9af74689d5789886f25f4d73868ed323f22a8d56d05182050baa0d979c1eeae08bb31c7c46f293b0bf866dd8116a1773764adb4a1456bb48d9f6ac9ede14e9375bc81bddea9439a2a6ae4c02dd5eb45baf75020c64edca5dd0bf7e7a5b25ffc5d55c0e9f7e0922b21f339ffa1700bead442d1f4ea31c5cc1fe9786a9c087e6565fa8c9f6e23390894560bd4c0795eb765115218a0e970de5337d3044897734f9a4915ec85a403bdfcbb07f7f2527cac35b2102f3a4166619ce0684ddd9a65a5ac46f60ef6c09495e4be80a49790e893830a2537b349abc0f891c1ac5d8ab3ff75d52aff6d2dcb5d1d7533b3181d35ddeec451ab20e76cf4d5d64b1071a82a28ba2b1c59ef5e2b12dd1b865c1cad8c3cd609bdf30d25d413bc29930d6f571a60b70498bccc74278b06ce02fb5a787436db846015fd456d838798426f30df8ba40d55e59fc1a8ddb67e10a1de1d4d3ac038388f1e32467747e94710010f8166d44e2062fb4023f1333fdd230ec8399f9163d5b0ae2ced6c7840440cb2ed6c5da188c730463466d225fa3fb9531df8fb47f02e4afd9c179d974764ed38642c9ed2a1fea734b6dcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2ff095ec3d11974a6003ff1525d614f4ad95f23f189b0aa16d4888e650052fe3124cd2df832e67e74c0586e33cb860964e79a21e8ee8e53784b815d83d80a5559700ce4900ea3d9643d3b3d2d99e4342d00fa91d9768757901392068e5ff27dadb896f683c2a06618c35a3bd783456fa92de04167d9e8fa765ba06e3b11bcdd07be33b75602afacff9e877bc22eb1d0b975f22247d1171398a316e81abb7d71d1f85a6b65ad7689d65c84d416fbba368718a4b7a2706409fd2c328f3c3e28d6c565c74ddd23b69f7018daef6ea4f464edef5cd7d471d4e6258c45b787fb90ea75b00c743d77ca0c3ef6263f33f3665d01b61018cbc057b89c0efbb46e426c4d24f7cb5e172df2783a81350376996fdb92ce9ee27893299b684c3996f246760fe521ff1912bb3fe6afd1dd6b0722277dcbc1d4110afd7bbc8e75737542e76d4df9ebf9759bb1763349e7b91b2f043240448c6a63861a3e7256cbb1f5f899d357fb7163a5ec5af27a99e345514d331f0b590f17d6870bfe69d0238419e0386909880a4a2e6d78731dfb5af7209be92efc8680a3f376e953f69ed5dcd03ee9fe87084669a2791fb2b5db3e8332a0ff4ca373632fc125f28dda5410ee2883882b60ad281d4d18b005fce53d30ab3cdb5851b72ff878d5651050e7129dd6f5cef2055bf71e03032457a850ba41fd58251c1d70d18e10f5fe2b9e795206030fdef03d55ebb4d2c4ce92562c072c949a7fdb866bccb7637a1b1f25ae0e6240adb9291f04e2231c2a181beef7b099c71c45bd873e7cc141af5250cec7478f2c2a3b55a4481f4630ba5fcb48e185fa56a016258d1ab96b590da114db1222e8a8fbe6a1658598016f5fb9a2d634472086a8dbecc0428f37c58078a0204bb3cddffc2fdb7e90848f7e6a72099b7027556d0007335417ef97049d0719e3fb349a6fe32562e94cc1cc5a691e81e028c311299cc23f99d2d27103a7a8d14f72905cfce032386802d753f755b1203119af6afbf100410ba2a5eb35aa3aa535162307f985fcc98f12beb78ad3c7271eee1d135b25a3cccd1bb38c0afcc686d91a5b8227f1cd86f3abb4e81b2f742915d6a181b96e163f39de26c63293b0d5650a6c78c0053bd3fb4158f5bd82018ad1e740c0a777d1111d4bfbe319f1142b26386923e7c878799f810881b481ec6485923b15bdc16e2ec3d1287dce94420656a5a2f72daab95ca83df73ee617184cee18d5b9f72ef0a43c74eb6c84baf145ebd42c579e9f5d32cd023e63a7fc2dcf9e1e608829e1eeb916b49afca9d7c166ec147b0b2acc9c176e8b7b0666397f095c0e3cdee251a8efddb741673eaeabc034a70ec6755e2039497197e58b5f4527f31e520e628d34406d4a56ce44eb1f1f8b174a1ecfb6602ca0c587ba8763cdcfaa13cf859fac5ce4ae4c47c6784480254e9ee4681200dd610ba94c587bf87f5d30dde085a165f35834188fab0c5a9dd905e1a8e9972ca597e0c7540749d789137e12db7299f280952b044d7e2c9b31fb52e18300544022c6a34041521e7ab753b96a25e0cb0a3a785adf0bb28360bc5ce541dbfcd0d28bdfe300dc60c3aa3131598940b845e5471506374d7b5c2dd43de32f1b92cdd1e965993cfb79be71686bba80bf69747773fd1ed1f1412c3c5697f8c2144cf141ff42bbe8d1b1c00c5cee170f6e45e0343a3dc8bd740f27500502d4a95a8d476233f2104adae17b43e8d04ff63b4f854ec1b367357b3bb2dbe2276c230acebc3f7f150b44091240eada6a179fe393312e515af63db34b89ed3bb95e56929b248783cf7f0a50ca853f7b1d645df3306ab46ec13258e337d00889344736ecb05b85ce3b8aeea0172f9b9e97f904a05e367991541c3b6c77b008308ea279cbefbf899f3cadbe71d5e3a7b9261800bc6ce53f618453522ce4d8be09d8da1ddf67cd42fb13c784eb8eca6b4ecf384108c287783a8912a36aca50469b71fb34c005c84a2b8f2aba9a5fbd37b9cd1d4abab1e56a6fd42e44c0a702e7c59f5d9a3e9628bae65040096b934098d6e3f95628d572f135a3ea7f9a6930818fad36b44aff8996cf7722d3394faf01aa1dd3f0c659cd9900cb0f08302c71af74df710c15ea5291723c7f0ca43f965cff70c4bb2c7314a8cb2e67f4b4d7e3544f4d86b0d168c58dccc25ba2aea1c96fd6ac0c7f2652df4f46e5c10139f0fe29e1c7b0a6f6c6ff132975e291293087def93efcb0340006f02cd466e01e31557fd6af6cf044df1ebd9c12a12fd2d6336702ae32269f74fc1cfc28b25067dd306cb1df29d283a67bf3d8adf91314a48bdf4b94ac93e2e9f30061180b4ec78cd3643e8cef872012a325c4dc27391dc09258739702e2924f4c99f295fc0182af973da3f9b6ec21502fae178c6b5b53b14d53418d3e00badb00a8be4a76c661ca0d8855ac2c820d7cdc177428ebe6c54596b3c1b55a8edb8c6775fcece5870563ae7dae0579972097f075fb2069e5f8e9b669202afffbb92e07d35fa18ab1127e2d81ba36f0ea831cfde4544dc3383a50ec4470355b41da33e9183c87fa062a6678381be197a4cafa29f0170a841519c83494d1255a98b502286121cadcaa60a541cf45da046c194b6ce58c1e9504b4856812e7d38d531076fd761fb8b723ae77f9c2c305cd580dd0d993c83e2233146add1ed4a7954ec39d0699c6c4a190f40e290a458c404bb72a76d95c6c4b64a24d27f0581439ecf68583450fbb72f4a0f4cbde67e0269a4c57e06be8ff0cfd6ef8d1a2bdff9f44c105b6894e8be818acb79a9c4c6ccbf30c95d2c996f6aa2cad80d036bbe11fbf32d1e2e1b5182070f737e2c62c8009fa023e709e98ea64ccb897268ad043b393501dfbabf2fe1175ca4aea162f947012396181c309edd20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h31a55c1daa18b19c8bf0fb2aefafce0bff920ce55bc9eba811415dfe3310d64860ba28ac970be32f021c993e672ec4f0fba3ca37f4352e587a2225a43ff0f852115a20bfd04f27f981cd204062835e166bd12720345f8e641581990e4474a19e996010c45cee37e9dd3769ce3d04755b5e6eec4c412d2338105f525110d09ac81c235d8546396bd69cb49300717f1eabc50323fe399df9bece8740f07ba2e355b81cee24e38cbe98706291aee7f0d9bc25e926b1686cb3c9877f92b00d8b0935843b2b50d3352256950e663c749538e1ca1b37746ff7fda5c713f1ed3d188c84879f5f2ce7c7381f84bbd657862a5df1c80e560de9302c666c31614505d20e339078694367279e878646140468ddab94034db753135f38795e050126f20ec7a91dc0554496e752d30d94a92327d39290876051df12c668e1eea96606dee9c708f38108325bd65c959f24aa19941028748a28349018df4393a11d9315e9556a706ca196ca3bec312b18dd43b692b23ec24841b220f9b84b1a73fa0a4085eab8a69a08b7c408b6aca0ef1b605f6c041f127a6bddfa8017b13686c8e4600019e7e480fc023ff1b87fdb540383e9940e2f48e50f7e5ba740c927a90f7cdc71aa3e40fe7d3fac447ca871cb096061640f5bf71e8826b371592e8f773e022ef2f3a554d2c55baf1650c9450f276abad8dc4b11e6f3b3c298f7e36ea3ab9378f8e35d374bf6d15c77cc5765326efa0f9a451a07a1a241bb1c24fca2dd871cf7b0585cae7b30d7124e3f4cf2f08d5254a69b73f20210651ebe5ce9283f3b1974f5b73ae26d34fcae176615f89f6f75cceda79e5c6edbeb8cec07b1cc7e7438ef4447bc4801e6ad6bcb61cc33a72fdd096e6c95bbcd0885c2e563dea5fd7dc1f138d338666042f8bb311c9ff7f809938d650c4da900e5c4d61db4cd96c31110d5fdf0747c2f1cfd6c1af9fe47ef34f3a50858c04421ab12d55fc9c2f66020bbcf56a4152c948b0ea1303f5c3913b40938c63e028de93ef23541fa1c1362010c4497078cb068bd73bf62ed43dd33d05232a6b54ac730988be69ae78ef4fe8d865ef7c250b95d853b6190553a68410687d01fa7881108128b996b0ea9102254bc98adcb6ea0dc3aa9f2902037ce78405111f5a04ee503f6a85701acde76cd352506df27c13f0f57a257e7fdcabce9b8d5c7d324f898381c43d843777e0cabfd985690ec6facf25ce335c5ba8ede00ae64d31af99308d9f6fcc92ec7e3a4a25f89fb82789286a2a9bf6a3d581db35ba3df75d1fa0dafc02c2acdcc03f3e7eee36416333f54647a7e257e1cd8df81994c5012569079bdf52aecd95d30c54a4d8ea51ba7e14bf01575966991118b45f4696d32e2d662e09fd45681eb7ab72c2d64178ad4d0d4433f3ad578d0f8b0db79449b00055ac05a5f8221b8bfe670df3e85bf3cb1a61a27f83c55c706931956d76b7ab4e887b70b9bdbedbacf8c2ebccf8723adbf9191a4ef96e038f1f37dd76dad360c2ea28b8923d437a68a8faa1f6e94b367381770f55b59b071a908ee560820a565209137e2b1b17995e5277dccdeefa2c941208fdcde533e224f1039d6f4cd9669ce108159e774097369a59e00dad04bf3763ba40a76293ee3d07cbf2fce0479a5e0a3d672af167faff66b4f5279f9f0773ed4bc348d39197deaa121a931b2531296c5010fcf6b43b1dea41104d09379f0206c5a369e30e63ae2172a592ca7d41e804b7508dba9498cc8ae4542a73a73b81f20555a51fde579dada19f48c3a0eeb2cd9cd05f764e364a97b190b2b9206061b4af058100ed23f5a3cc640d3b7dae825ffe3d506c35771b382f505665a973899af009332fda80e2aaee614b651e8c782f0519df70397c68925153e1553931638019e0a4d46eee4269f4b4b1434419b7c01ff9f1e2c5f3751037e20291e7998b934c29b4e372b351f2ec9d111c60132153d6bf1e59c73fa8e13fbb9729ee1d6085856831a913702e4c4795d0501f2b4d4db92a0493aab13dbac02c3e2e50c7dd49fbe0d6a97d94c1589f877492e4c9c613c7db860289af8ca1a9bc587b064f340456fe9a24c962771e6f0079a0e1a385091a2dfc5fbac315d54b58539516e19acf888ceaf1b9f040d52a4d2f104b10548b071df40bcb9402db49a095d9889adb4b0e31cb0094b26a99b5036e4414ebf4152a15b85ea5f1c13ecd4cccae69e364c13ec38d25bac86f8c8902f2a09ae9003a6debaee55c9ea6e9271e083c1fc454a038d915cbc1d541a8c6cdfdbf79a49b8338116d33c932b83122cdd46c75df70e19eda1540822b78ac27d775243fa43113e7f3d87d2893a6e095e2e01ba2bc5f38ee67e60dc6e8bd9a3704e85a50f0fac6c3a9508bf0d3e7ea156dfd771bfc3b1dcd9f6b294648c2690afc03297e01bdef377fd8bc2d7929148f9c6db4ad11eacdd20d33647111feed15e1663958b1fca3692c786232ebdda1adda7bc798b9209c37b95247c4301ae47177ef8ff260a11f3545bfe83e712ada0d7ec7d655a9a23229646b1bbc371901ff73a3470167f98b61f0fae7ac6e88a1805a5273f83e5e992bb3ac4e6140ee787dd9a80b7168ce3376eb849a2e15c38bd92a319b108ea07fc060f56633a37b10c12e5975865f8565ec061d16ed7187c601e24ad767a51692b0929a7ddb02176f879fb3caf0afb5b578052ece46c500071445e30812782cde7c3e71d42ac4720e49654177e2c7b34a5feb89e7ecfe5e91bfe2b7e1fefefcd6492bc5ec65c57935de6bf5e655c788d4b3af9ebde9640b113b999dd39907dd159d9380cad48b721cefa0bb41262dffe65bbf03dd1172db4435d22e4bb3c66f09a982931d018b431bb7dde758278bb1d22e9226a6d6d869dbdcb5056a7b1ea592efe33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfa8780945fe33c3fc92990afeccb7ea4af80c51a6156c04c40368b6766f2209c4fcb1c02a75a69dff2c506b97a39c754a29f169e896ad00ae4f9df9cf4f9b7e56883f521561e58dbafdb1edfd98895c2313c2ae24394ca43278053ab57805d334843e072c3e347f0846c2d8066e16b0edd252f6f375c71d3949e2b6a578a4baa7c6e11c64abf7efe94fc08544d4c419104f88fbb16937f41bce35bf7f4dcc80adfed357f47aeae4c6318598692eb46a15ecff543b069d790b101012e17d8ed7c9402fc6ba641410d53749291c7de4900b1275d4339da6647a37afa838db55b2829419aba3399650ce8b7873bd98042d7e462fa14abc0b0dc91bd2f91efd84fc13f5e0fd9b4c15b8ff040a0900f60697a5d76751f637b6fc5acbf8533ab7b62a49b09259febe84a87655e8a4173da7c8284e9e7e5266f68c17a8f03fb21c513d47e8962b5ca7366a5ae64b1141403b7634ffee5deac22fbf1aa7c6b8b9265de331f5f05d06ada4146c1ab4c880f5b0309a4b01f7e1779cb938503a39370b53e5326c84a9629470a86702211510804a199d172452a56f33924594cb5c74585bd0d5bcd3ccbad098c35f440648ce7f7c0a236829f4c017ac312f13cea5f497281e2b6dbc6863a69e6cef0c55002d947a6da45ddca46e7029ecd61634def7f70fd3a0d8d1de39530bdc9cac63b75512f0c17a3cc4b9baea3aab29c56c547ba7e2f8b77c950b38e18adb2e7ec84793325e85c64fe83dfc45aeabc95612af760baeb3b356778c2bdd05c02d0469bb2b319c59baeb730cd239d8ca9006bdf897ec98ab9ac461084629401cb852f89027cd74a932b31c5149c5cd9fe0ec87181efcf69962bfbcad14487e046016eb07590b6d3acff3fe19f3a128214bbf83bfa0fcae90249c357d71205e44f3a611cd47c2437260264dd436eedb1952ec151c984f5ff47c5aa937ce1b52215e31f9c03331716f81ec5e42da93003695e72d9ca2e2f62e90733e23797c49f1ce653df42fc9417230cf55bd3b62e20d6c1365b04941ec36ceb3e52fe98503bd992ec915569ce6fcee4796c3e9f83d9e4128e4a72c72e3a5486cfe93f5fe19ea70405e4f105c02712dff4b49d0ab0a2470a5ef22a1e0c72b6472ffec3bc9f9d6863364a19f9617268a41f6e8416af354c79e3429c82247c5bccf381cfd8952ab0e5fd72126fefdc9fa4c50be8fc0a49229c3140037498c9a5be2203c9b9701dd32696327f2e53b82a4f09799747b248d525d537fd6f4c028dc48b405d0de23910c79a4e3f68fd0a85eef609ef654b176e7d965fc44c745c76e263a9b25df12d97a3e549bc74619011082e23bf30f8c4392e0fa071d5cac332cf57b6964b672cc4d366286b428846ea43a68df20327c9394c9e650573866406385eba332a38e5a58e578b1a58771434c2eb53ee93b339183c79af56f724af140519102104658c50246eec8548906e6d80858e77053e0715536f66498c82216e37621dae7ced4a2025cbfd202f049335e8a4f22b59054508e301bd6e360ff0dbd37d8045f502be276a6b89e74b60c82d5473276106122a1450db9c5049ff213b7fa3b06503cefc5034a6d9987c42eefb287b0674b569e3d904ea95b1f65557e4190f3c8f6b1844eeda923c58fb0f3eee8aba5513bb70b21446a2de915414f1a429ac2471b9412db8ed8a99278eaf4eddc0dde8b2792e5d956cff8f78b8f52348836da8b4224cf36247923a6e8a570b75ab87ed75b63bf44af9a1eb3c5af1ef155e677c9c266d9c48d42ec28890445d5004db8caf3729035603adad1ec30d94188690976f31bd2720674c71e3349520adfb862d841a59bb8e9e9a0d5fb32bb761214f76a396aa2058b68022e43aa420cc1100c33c05bb8aeabcbce5a8cae67b60ac5b4f0177d756f66e218c35adca9cbd1ae666a827160b5fb35579253004a3f72c51e4b1dd0e5e1753a80fbff08831bc31c2e529955b69228a145b422a6a6292dbeda5ad4417df5e4697783251aa1e17aa67c0e0e4e4d568d29767f0e74dd66ec72927430301bf9c44460d34afbb44dc33d572f84a1cfdff2dfb6c58692137c0bc165f84ee26eb3641e1e360af01cd5bfc862ce89a1bcb2b2068ed45285f3bf83562a8edad9eedf2235e21ddc2b169a5a2fac3b065ad44a2e520f395edb20a4fd16c05d264dbb212dd1a34e8aadb0bf04ca8709c611b05d07c9d50029bd204914dde573a992d8a8e37d7708da9aecb0df43a0dbcd756ad03254ed7ae15cd67c2df3552c665b9e6ef2a5a4cc9338f7532514a137dc6c8ebd9a684083fc77b906b6e1e203e4e654a65ba8b41ada37f42e3d6ade4af9d26237ebb84b69cf8e8cc6c5c9456fe36fbc39a725d0d1e45210a2ec9d6bb7c95c7189316e14afd7b481fe9d7d6ae5a6e46d856b244cf1933fa060489f448b21c26399727c602e0ed36e635c6a7ce97d5460babe404893902c08cb20cf8446e394f23204ea8ad69d5b5c1f689a05cd4bf7f26b97a552aed374b9a0d5d8c5ed98a7b1215ca4c2ffb7a4de2afeeca325b6d20240af61c17eb2e5d74001282f64d5bae5aa80d8c5ee61d16e795d41eceb473af5d144df8246c9019d903472c68cb9f48f6cb109f3fea391d5d9275094f9a6361466d406c270502b68716a7e1eda65cc02f98006cba2c1db4cbc581975fde4eb44c6114506fe7ce1d2cc15f0aa0b5958c34582d949286921ca831c05842d9e8a632d1b5db9bca4f1b90a769f6818107c0437df1942b93eefb523cbe32ee6b73fe0443e53c5e69eecbaaa24c8d6bc01c09ccf8c57c9be846921b4d19213838622cb0528df4cf979b6418af84fb1c084a7e7b7076acbb3fa1b53d4e5d420587d1fd9aaa016476c65713edce61e7830d0e2d1f32e68e6f4f3513d7a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7a52f52943aa836395a7d53ea35dda9535d5b5d5e3e8a00717624c132ad5687f0cbc64980620b8fbcd441a1dbf5ac75aff25df9c68eb65cd8e825237dcb696ea04224f6c91e836f6a21cc420431b648ef3ebf5af5537e4b389794054a7d4e8981b6ecb15ae50809045b4d3a1baeb3573c68287fdb48358df20c333802594a51fd89b984907887ea0fca00929136bcd504f905b8e217642f74b73770b5272d260ef843b3fcc0de2b0ae7a025a015c81d1f78a5caffcbccecb84564e2cebaa3d29a94ff7cb5d7569044a4a726894011d6b2a0e98ca1d5f6922a6af9cef9ebe223482a5326d7a80d24535e6b7ea67b2023cde8986ec9c0d578632e9b5b3bd46bb7524c1c94b8184949c815189a8985e07869127221729f350b82c10dab36021d10abef99cbd270fa79a41c83aef10e71d1c8ce0b7818febc57ab7a500729fef5e30623cca5a6cfec9ff48b74b8bcc9554ec0af41d3cf6bfec67c654e387811d74c3601c213e39289350d8ace61a09ce15a79ff2b841f6b00e5ecf0165f67a7d76ffda9cf8cd89b91854fafc9df30de8fd5cf22ab5a20f40b7839abcea5c34adce959ad30703deac233147a4946594e4394176b65191b5ac49cc414c1bd0fbb7538f35d095202f0959cfcdf3a10437e2f810bf60ee3600dfa337763820f87806b34381916f67807d2b9d24b9b78730d720472cb2b0bd47aee7093de631e2f3c1861de02d44739c99bc1584b7d42b7fa0515426f76f4d7fd412557e2f1be6785e6664938128cd2676cd8629069cd5a618b8f6d496058fc4d8c397b02dc450325af4a3b24cd17b1a93edc07585af48bf33abd1286eb3ebcac9e30605e9174f5b2b0e0623f5af6e8544c936b000974d2059f487e3839aaa914e00eb15c7df5c4c6e38b1303acbed644d5edefd9a6f7c4a9006bdb14552efd23bbe2b95464f68d6e61f7f1c05dbd4bc850f1c3b53f76963ba15f5cf01ead942d24ec4b87400dbdae6cd7599efab802d25de8be064babbfe4c84f78b002eb2c2ddef413b9b703a117a805d6b6e7d957f507da093ee36fe8228966238ffda8f456bbb09e85db25f6caa12bb9846d9258d4cf33ad55a42241f6408688ca31bb8ec93104787f499dd8bcc29b962f51d173a8a414c9518cb0ed7e0a9c9fcb33568eacd3b632155b0955c72ddbd6727c09c749fd5dc4733ae13e774a1ef76d4a55c58c4ff7752235e1365e4bb722a9fc7daeb1dd52bd625775a4fa24816ae4f8f930fdfcae9b8df98d13c38c6fdb83a700c0df2a62494c8e5b5d5f0b1c940c6a7e7e1747192ff562cbd3f6ef8ebb714a8f4ef3d2695ca72b7d9706749fc6fd1ea745bb090e0985656d2886a62e4b1641fc985ebec10e8031fca3762f35cc7cdb3bc4865fd1739afe57052d836eb83b026188f0be1f18dac321a37bd0e361a37640add64ded1b8c1848bc4639854dd20c359e1850328be3b5053eb783fb84d94c66286244f02f5fd748bcab59ea3aafca34630e5fa028f4e821b60a40d2e346b4cdb3a6eee88e861efa45743f0439f7fedbbdfe876a225356cc6ba256ddab781cf8866cd471367d53530d2a8eb8ca81e79a524447371f0abe526e15c6ea6f78c02bb1bd6e8eda2f17719020887e70211d05f07862c2646c5f8470407b3d11cde8ab2e7143d04d2bf5108f4cbfd87616582574d96826c56a9af466be0ec1f877f113a6ed1297136ec4b3867c7ae3ffd2e7b1c9d1e3d0535025fc0595222e00411468222cc411a27850a0e176541e9d8883912ac1135ef130d18f2433189a271bc03e6ba1e9c7bade701039d5371ca0b1e9b2dfaf68b8aa2cbc1618151ac0584c501e2a0d69b89cf1293a19340a447eb91e14c7465818f1038f4a01315227c64b06737d92f95a7dda2a65e540330514d58c3ae37c78618aae00706169ff7fe23e803d820e48a77a191d8b8848c5e2830d50be8ee18de10982c01577ce2782bb792ac5adeffdc4a5e4dbe5418417c63773398a3bcd3b93cd6491ff585fcf47e4853374e1ee440debd1b0efd37259ca943882666ba0200a01143e4dbee1e043b61d12c95101f14c88b66acfc5e7ef2b27e734469cf52ea6c04340ac205c7e9f47d0ca80927cf9fe0beacc81b82948e1a7c8bc0f2fd5b3e8155781a3f51ae2e31cecccb738be35947bc6b1dc649058bebdcd362f68f704839e0731f1b087cbbe2366b35b2de789949a47fd03c3dcdc533ec94c1bae8e2f47faa597198298b0b045764280f86969bd7b88f55a992c69bb033b4a7e1f08b8c515708098f24cd1b046c9692d6b9500090234541e87ef62bb1c15493bc137b0c9cf847113ffc9953b4da422ef4f0e1e8f9b5b06270f61c5c1c8e7cb7be1c286240c247b82637c8092517befb353300530cfa5c109ed7907831759d0fbd0f25e86a795288fc6218a286efe0c082e83fd5cc1105d310bf7c1e9a3a7a96e743be2aa3d3d95c192e698c3c015d0e015733e1b658f96a6b8b6ca22afbb4216f7ce6f01952e62c3e8deb32727ed5a0056cbb0fcc409ce0e9e6931e4fd09ed34bcd6abb020d766e6cdea8d8621337d1394a2845c6344699acc0d3017ce8cfac92b9a9294a80862795d59266ad876816fba7491205d4e0d43e691a932c5383f1a3988683434958e9922c8a80d8da44cfff00076ca90e8f2ecaf4e69b346e27ccf9d3adc3c55c13a278ede9342d47ba6943ff18a5b32885561f1618951acff8f426d0bfd59b68c44d88dd9bec2d2d2fc6c66f805c3d1abe6656fec782739ef0beba75160d1511bcc2bedba5b87ffcb4dd6887e54ae2f3f64ff01e0e1247e934169a53e7f5427230d2f29d67485abf76cb9ddb3cde89b1ebf3bb56624aee7ffe5535117ba18955da211ba253b5e4ff346ddf58cddc59055e45cd0ff1de18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4d2d8f78b2762bd82558eefb8073ae99eec833421323ffe3643ec95f7b2d3682a2a1bc215ffd2eff08b726b481379bf2e2e9136859421692856db255a986b101252ce3914bc11df5a99d0b3cb1dad53a2ce40b76217b504821bafc1cc05de214b7205ce13b17fffa0c63d3944814214c7dd54ec7ff022de6e6f4c015659e4dcc29ed5e2bb98051e904fcc05bb860a37652b410a44adb5225587bff5ea07b1a260aa6bd9017098c7c00b3e325c8b50586f43b0ea76063e603f157d6a90b08f1d72646f62a8412f180b688203de9f669e8e02ad3b22eb99a13132d64f3e4f38a73fd7c499535d20a07c5978280a87fb6add0715de44ea0d9ffbb4b575eca32c6269cb8833c8e3351f51fc09bb6cb274c2b25b0651ad4493cf06c9e35205354f63f172d283b303eeefc68f4c9e7ef9346b5c00cac6d909f863c041390bb46af384879b6ab871e0f8db959b253cad68b50be063c1d646648c64b5f737e4c4f778ab6068f96751e63e8889213cc5b83ed74dfd3215b10fd47a44c46b44e042b8f364d95fce75c57304b89e32be8ec19c88fabe35eb8f184a947d090f0002f187ab2267d2d045fa167ca813c3cdecb05a31d12c6f7aa04c413365a56a0041b43ec02e25c4e7afc4c3aba9f24da45b7eaea8a0dfd17d2912ff9083ff6e2b464faf519430015628714e9f30fecf4bc29a5c6fdac41baf4db1e22e1c9483821dfb7271cac6047d2f5727a041c233f41d792f0bc440d9486a87f89c41cc3e4ebeb8cc7aaaaacd3120961303b6dcda0e72186f97639df65025ced579d2b13c7f9083b01d965c7c9bfacf096432f7c275b0f25c81d95e182393232ddae0b4836e494fe6a161ec10f9a8776fe9b788be8ba4ac0916d0a91a5c19bfd449ad7df7cba73b1b0d41eae0cb9db2375981ae9a62b9012fcd3267c0500242fa122de2037bd050fe28c78bdf5124ee81a6bcf6e061b14c861c83ac38a3bcfe5a9715ca78880ad39fd047c272cb2c2ab94811825a4dc6f33d11aff808e265bba1bee1c38f075a9f6904f4388c416cd8c6dbab4b7f006e8ba03e97e6c668dfe1738fcb8ae82265b316694d4dfed5fcaed6991fea0c2be13de93c2c7f99ac8fa94ee79709174c47231e2e183737c43ee93af2f889499b3cefe404884f17f098c38cd15ad2e585aa480f94aedf10214ed20ff9568c2e946e4eeb8279754e1078bedb52340698440d78aaa2a931eaaed6b8ac589c8d5d5ed7570f675e0046300aec1cf8b38ac317f03febd987ea622afc1f22778549f90b0e7b69b5786893916945325d93d6566fb433dc2788e56dd3ce7577f1c24b16e513d11771baf4972f0fefa742582f360c78f5d5d25e706205e3690d9d41dd4ac229fb9929c4f1d9506ac1569479d522bfd9242214886cca39087892e617bc08b9a36f9e558d3f6efccd4bf16dfb2d3e5954683104f9f943fc3dbfb31a462176811717cfea2d3f8e38008b6ce40510eac7cf1d960cff0860097854712b40cbf41406ce22e7ce4e7d1dac2a9eac22bdb98d1799ab12af05f0c7a63baee24bdbd5e77e97a667671822ba7771fbe312ddba22e75d9bdf190e1e5aa9fc5636b0f5157f0240f54ffc0bbab69845675eb9daa971c43df8214017e89825c4f807d83b44a06e63facc0bc56ab24685e5b10c90c88e834081244b9e7ed3d5d37fb8dbb2259f8c99b9cffe3d7620cd9ddf39c04c50d8b9e42072499a12110e52e676eff7964d9a1a4a93362a59b211c0ddc087d9ec7fcd101f507c1c09322ea85fafbdc93bbe6f8fbb8d315cba44e81da2ce700c76eece9d00735ac08bb3d7bc9ca58a5d87644aed40ece01f8c31bfc693874210c0a9ef590b4b6b2a6337bed97f29865aa97bb4bee2877f5e674bc809dcdb9e17e73ccf41ecfb6dca53c41f5327495d56726a2b14d69941b193a7a7e09d4f6af7058add1a33195d19903d1cd98f883214e636ec5302beedd68d6c8ecb61776305358c97376b537d352dc651065ea1db32e34a5fde034a1dd4af2fcfe9be6f1ce4bf06154d6eadc5315c985040c1be2d6d74462a11fc63f0464580e52a7fc240ef8fc9521d63ed3153f1cb4200baf4235284708d72f6c07c11618f598fc028ab91451c513963eaaa7ae29f214ac6b4ad7db09a5c73b180cd39bb7dd3ad5070278d24b2012112f17dad2bc95e2815f4e6b681929a755adacafa11b5802206c55fc9287689c8098b19b43ae976ed5c0ef9f5c5e6ff139957070071bfd22ac958716f07b2bd9643844ff1ed396dfe448d3a2b3208dfc21d4ff851410a89f68f88d580d2dc6ee6c0b0606281ce208ae35dde9ab8fa02335d8b4be9631000b2301b3f694f94fe14dca70e0356b82739065d7ef749fe6fdb87b97fd79794ff8b28ec02528982acf02f7529f42c78312860ef40fa6bbe28d83b15a1e9d3d4f83ba4e31b60cba9a2b00a836c2d0d6cc3a2c1d48989e23b67235c0a64a5091dcbef2c1358197b5102e9643b6604591b32bb8de941314ae82d993f04119cb7a6334bba6bcafa197cc2bd3cffc7d065ece709cdcf2248b481d38c2ee94a2dc23a2fc59afa4688216bc4bdb6701c65e1e27453b6b595dd7ad17e6ac2fbf99d77e54fa37514684e27ce2a3778bd231e01872860b10f2781443e93c02b22a80d2f527b3d4fee778bd10a6b9371cb5e5c3fe149ad6a24a7844199771c788cc3ffea00556a64d298879920374b24ccfc2072d13e969e8016ce046c89f2059d70612af3199b6331068e96c84351a2bae8a48278cdfb51d0fe9cb415cc9d1d4e13befbfe77823c9af148b43b22a5f929fbf6a471e2b11f124297cbdf9473ed69f63979e548dcfc657189614c5f7eca8ba325f2676043d52d786c5c1aef894db2b274f68fa4a4114e42837424126d0878ffb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcf9c4af1e16113b19ac0405284dfd28f456ee4107e6bb47fbd359257c38ccee74bddd4d64dc7ef9111a4e78a6b88aa0ab2b5ed07717d35d4e461971843b7cfeac31c24fd24583cecd53c3aaf426453aba2326ee16c43e1af83bd75747d0884e6df31df127faff68c152167ea8a3fe50a4b4889926aaa70ffeccbb42cbee43f26ee158bc04c542382c43e4472285d00bfd4424096549d5b5ce256d04e22fb182bd39ae1fe2474a1ebb2a70aba03a17799eef8c85e06491e61f477b4398dd492e36d760e1929d5b4d149a8dee3668dde68949410a20ba2772f09515406f1e268b74d4d6e4f1eb73b182bd1a3e9949606c0cce4cbaf265114c260905d86c34df484f5296f17e1b8852c66670bec322282b28ad4f7cc21882caca6e597f1cfd25c653e2695f3b1016a9d6bb05f5f3728b104af46310cf9c5f4b36ab631527c0091a08b3471d4e30b08db24c5121278c587506802df2d2c39848efff7f36b3ecbc1f4a4c0bc4eac6475dd040f42c0c15d1c100768ebf50ab845cb70577c26ca2d830af547289d872b08175e48f4e874b70cfb3956c19c4b4b19a63f83dd635edcb4e6d40a9fd07d8837f2bc0ed28432d0dfcf3ef06b9b797691cb8b818ca0f05c91b0387dcf65c43e64a33d066c6fe4c19a67bd45faa2250fa518d06e2d42d5843acbdfa36231891778b9ee0e34011ed7224880e1c4daf313e6ac1dd24627e06cec2bc61365538f9e47ae836e4931b18dcc08b25425161b4abd63f60211ad9e30f57af55cb1611f21c50b2473460fa39ad06b4e08383658f0578ef717dc46f41b30ce5edbc832025773afc968139acbdf97ef868afe9cd6bd6978581a90737eff11b40fb84b0939a0d659e42544c232e507f5ff95c4443a1fe4e2ddf5a71b3945b58b9addd328035e8997cd68a4598f8e5c411f7cceec764479d16c439d58296d0eecba0278396a4ecf925b238223e982dfacab09db14a91126745373f731c93c6f00c2efb8268dce15c87cc731e200b9f409018ba232626400176a5cfdd0fbf1bb540707f4a44d65015de7f225b3fdcf23aebe2897bcdae0711569eb2413bc3aee1f70f1fa6b70100643e2386b1242d561ee73ab7bbf96b7e08953331bb09c9bdd4c8aee3c47795504737c19709d341b226e1f842697b3ed7841199d6e5e1b215174f569a7df04108a3ebf78775ce5d51569824f0fd52b13d52c365e88a64b31ce4f081199d19505033b8aaafff6d6771e86d9ca814112a4fc4c6067c0a814ba2ec0581a59ff546e148dbfc9a91252a829a55283120545141890a5db1f0f04b1d26779443566213136bc80c7dadc20a42aaf94c037afe2599ffd6dd17dc64d750134419493894e29c2906691508a952c7cd920cd09720103069bc43c8bb57cac6c8311b25be6bd7669606a83117b1eb5c67a9e024eea834066e56a287196082f166667304cd3d6c7b464e63d32e6146017e1f1cdae767fbdb83d955b85b23f88d9e7f287b4203853b2e67180f0abbb1584d14a651ae484b3e35dc980c2fbd48573d0ecc5169ca77efbcbda2fb45e1d44e88ad8e43d6d9082b58582e1eb995ee376838e5fac951340b45071e244e573f6fb650643cfac31ea8277092b590b2c4af68e0f1beb01e1ce11079c519f918496561f558bd8a8dccb1883ec7068d1ef7fc5a52b3085c7e8269b7d69846474df69d52a8a3844e02de769b4d2550d4ccbb978b937968c112bdba6f3bc7455cf9a0cfaeeb83b53117baa48d83dfdbf052c93add8490fcafbb2286b1b87e12412261bc52f804b54eba328fd98e458e8206ca3d73a671af560919b5f35cfa3bf6ffca09bb4d221bcfcc2fd1b9a64a066dc61e0ac577c09362aad00a913e91d3c4062a7b2a07e4b1f5e0a5e4f797c1bb0c852209caf36bae396ad45684a9fd6f27ec3b3af18ca6ce09f5d38d24dd36f20a26a623163db47fad3b9194cbb501180549d73d24164130587756ed2715e86ea613e8d8c722fc1f7a8e7a3216a169e6c91645390e1e804eb1026192233b2811c1e57a8affa74ec021680e8dcb3b0629b045a60ff6bd6fd8fb279e3c97c54918031dd7d19a8ba6af4fd2a896a5682eabdc0a1fbbfac71912c33bc6d1df8e214794a70c114d2b1ce821b3bc55b9c6bed8fc8c12fc6c893853d4d9783f7201a6bfa7ba28ddc95a95e0e8c3cf7f60956813b5b5a44d5017a96d182caccfb60003a7b2faeab360fe24a85ef52d30c424dd5e96abdeba58468c5710fa2884cba386ba674c2060f2fd803b43333771507ec34994278c2e11794a75a22bfd4b2593033f7da868e3e40c1dd3a92cf66e9b6ad09588502a3108fc8d10e2e1175b3c13c83e29fa8615fc1598aa904c757a635266d41367be7e5c9999fa22c941c36c4c8a07d09b715556c367e80d671af5ee3a9379522e93f91035992e29cfd3e3d7a5fb3a81cc6acf45656f8be7093cabfb6d6674a207620a5145ab254001cb2b54490cf28848f1fec514371277caf8e4d346feec98f094c5ff4091268b17fac868e71082dd5cec7e0bcbbf7cde7e168c72562950dcbb4040605a9f88a9fa239b6b3b4b80c85f829ec5a9d989d530e47d2b9d017a9a31bbef1b2d896b31b67df599c51ad01a229e10640ba916d647bb1d03b4a56352f9b2382b68eabaf468a19cff216e69b468d6ebc6b0d073d7224b7d43652b2615f89622c06e691532d449d120e42ab80dc2423c2930e04448e9e92c35371ff52aaa2216d98cb8331b13567d74a27c55baee81718e3394dab0c8122fd233e05cf187cc6567328796c3100db65b2640687fab9475ba763b52b9f9e1baa7f2e0d6fe7015887bb5c4d088f2fdf7d8dd2746158d6c8ef760a4f3ed482f542be74ae0b23d29b30faa6099c9c63b442f2c545a27ec0102e82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8b481a8ce7141547efe1f1039eb155a8ecb0cd8236f1187e3ff8b927245ed086da16881316db9fc52181173acb7805c089754fc5f8c46421b02cc420e300289a627092a0f4e7cecc2a6119fed53211fe59b47341e9d3ea0b15059ed163dd668c5f4a7a3f4123c2846cb30b967c0b33e8753e0aa9b308cc16d1a7d5a098618f8b639319a4629a25a5eb738a090df171631a1f72d50f470eabf9ba7b31389b4caa24dd9d2c5d168b469784139f2e2530c65c52b8c09e53833b67b915ff8f25014f15333b558d0ebb33228fe0c530fe0b1e393021422618ee216b76c8cb269aef3d23856233a8cdfd6d42054ae48226ab405d60d808bdc952885571c891781d8c8dd006cf3fac147cd64869ee0aced8e8067524909f8cd84e24ecdbcc8ed6a690bfb7f587ab0c7cefe8f415c023341edefb9342454a2c75f185f11bc043f35d161f3a8835d0d19e1d6b5058f8c190cad7a3e06f11da435df1c851dfa10c29b8d911d1cb05dd3b8b1777e1109e039726822ae32cd70b9861ea60cb994acb2e6009edb313e64122f9006efa439b495f0cc390dfcc07b951ca2af4570526d85e7b805abce838ba6cf708a2b891b5421811618efd4d5ae2213bbdc8b75e5583eedade0e43435239aafcc3ad45586aa7a8ecaf1598680381c9e2bc37895e76886d251766f82cf1fc7fefb12678caacd0ba21d0b2cb6ff35a85250c12834efd3381775af88314bc3051906405a3ea656bf180f561462911fa07f45eb86a475527bc7e11b6a538181c0bfacba5c84de15950e72933aaf2225ced7a40edb5d1792de07b6467d03971f22bae1268658dabab6b73efe016aaba1aa0233751b5ef94c4dba6098978ffa65ddc332c388fc2f7190d5abbfd7fea5609642879c7594bacc88faa212b29cb327e1ee2c131d4af86134d193f50a0b6a6636d6e6b1a685510efa95b3549a9816caef3eb45e36559a4de43ac36decce547542caadf9f94244283c44539473af89ddce6f19c807e67cf061c79dd7f4ef97971a3eac530f77bf26e7bae85f582dd9d343c6f7175cf7956a7526608a28dce6950de87a3d269808df24877ae08849e13d7a4f5a6704cfc185e39c38deb65c936f6e53c88a1416955218647e47db4faf8e5d7a5af4b04a205fadf7e337e675954c05f280dc4103613fd9955e5d7db0ef1278f4f38ab5569a87996e8bb0362f0254af0f9923263cabb6d6f4189bfc185ab2289a7688792bad224e484bf0b4bab3db477c17133a8a9f9d91c118d8a166ff4a1bc3f589f43a52c4d3135267ab7791e4f233cab40e090dcbfcceabd83b2e49d106099cd8f732f27b7f3282ff98f63d6fee7e4d80fc45c96774c8019f9699d5a80221c2a5d7ca42f0e8255fec0bb7a6e7a0595ada8fee2cc27d37ec8cf1beacb39ec4de48203f66f1e2ad0580ffee96cc4007a5b3ffbcbe3b9fe5e3e71d4c97da9c99cab74807dc5d575c8ac33262dc26c0f02e89e9899746d1c9313962c93459b7497af2c672535a738f231144b24fc4627b4d76921db736137a59951fa2a4e834afe7e774681ff545c372dee4e65f7cd2f2389e84ffb007fabfc2eb0cb3d82393831010aa63f387df293501b45899cee98b05b5556a194a1a93937abd6169ed09827a3e61704c81ab0b1aaedb5c125c4a89917387e4c06f70da10d172c7a609668ba28be1e785a0665bab15b529c52847ca8b4b73f3a817900f78b09dd3d56f959ff6ea89383b1f7a67060d3c5b8c9e32e4521ad6799d6944cc1a376c27b1dece2189e5e115a7cbb6e4a25ca1dab2e03174744a17fcf3c838fc1ea741c79d19ba51e1c5167fa9d56e0d36aed72d307f341f479a683fd28f8af85c2237c27b28120e1fd02e37838ee147b3c46b0a2047fbf01f94592d7cc823830855a8f49b250e34f77de190c5380e1ee9a8a9052a171b974fb59a32ec8ae8f94fd0e4ce5e231f6bee3624f179b09bb55465ebc48cde346a00e583d8752239a9f0310b691e575b6dc29918523f098299009486b3adbdb83a680c721e86d76fda507476b0c0dcf0539be18e71b90c2de707713a5136482a276b4928ad911e21fca0b768975ecc5729df18265de4b5467adf9d01bb7785119c72ebf110ab19d88a6606d1ba0d9c41c3856f32bb347ac76cb4ca2ed41bf6f1c9cc287ec32b41779e7e466c91257cadff9e153afc02100405f5496b99457d4cde65fd763848db4502c4e6f949a764abe2075d8d59b2bebb54c3304b1568911d49c0fae80147e70a4a3744babd5e98cd3b2b978b094977cc7ef7f79b4cc468844a6f15c5e19845dcbda853bdf7dad08b37475087e6d5f1db1433c3cca26af5abe9b6d9a03d81177a50b792b633741c6b9c59354f4a2f4520892f878986e39bd103de7dd890283d0950ad6667719fb5ee3b3a6d82b4ee8a600ffc410aeee8a2ee1abfce4a2564bbc0fd1b49732282dd9bf304b49b2b5d106b3c01b46507738a52b2fe83b2deb5caaee7d14a36f2b17c1fd6290b4ccb388d8d4faec87e02601307e23e0df46e7373382e3786c4f288a4d58357498da4a36229eb170f196543fd638d19cc501dbef0cf0ddf0ea397a1f2b7a004750aa89731347c71624714680c5da76eb606899a52b2f4f20dd04f87f061f28fb6213c5213de05c7610c45e86652b7ad0d5e2764a09b475c1eb1a3b33f945533b4a01caf1b1a7488487b2207f58b40cf17fb6b60112a1e2b0c19814551d3311f880da81488d242b3b12a5453af9ec3c5f7fd836df7fdfb6ee37352b597dde9b1d4fbf526f9e71e023e0f91ae5f72e6068c2cd19df984fae5b3d4af337b9192298898c7bbb8f648d8f1ac6c5aae2ec55060528fb81478bd49855f105bba904531cc632c438d774aaf80ce258254b1d32e009ee9233a9549b952c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h811cef09afdf6d10cb1b10613a5f49b907fc040f853a4c10d4873540a1458ae3ef84a1b82d8a786df8066e42bc11102240e1bf159f9b8eb70640bf9a180dee6b90b71a195bab83cba4887410ebc6ec543ae80c0efc7d8d979e23dad29f3a34ef6b6e07bc09ddc2cb26c5ba9f2b0e0669c245a6a7347ae393d7720290bc88bdca1cb4b2f1d99934bf4f27b3f8b10b75f75c09e034d36181584db1cc4d4f512944837d71301b1525331b58c93ef7d3c5988bd9ff64bc630d2ae5effbbcdb54fbe6622ab03091a2a4338df6e70251886855508541957f26be82e0eeb91596b93dbc1f39635c711a144c7a067d2b7131ff7c0ec68cf3a1b01bfe935903d587be2da7345abd12fae13026325f43f68fccaeafcacb08344a4090de448c5d75b1244a56ebe547d2f8d48a9b359bc742d8ded5dc7c8f8e34354874699a129f9305cd8baa49965a816b2e422ce0d80b1bdacf8beb721d36d26d8bba1deb77052e8379c103f41114fe7a0728c4c3c1b9d0d876124f892bea678058164ee8920841cc802f9c55d689bc4acfb5f13197f709c1e61acbdac3d19ab0af86a1ce8464428b42fdc7de51a9c258a64a355b7ea9a48586f353fdf2a3eb3d261f7fa93a762abbea7f1ffd37d9d99ab43c24b70ca1ab8346a82afdd75f08b4db64b5e8504a321297ae08d2fb67217f6fbcdb852175fc41f9f7d79c3756977749ef14b76b4437b9f19dcde0dfdd88c7f1e1c7e3e3f7d7214480d3aa28ba6b2f11e58b09e8c666ed4b7a956c28985b5cb06c495976fc17f11b241d9b31c68690f8f6ebae03b97bc959f682e37c79ce724a46cc8e3bcd70e5e9c14828ffbff789b651ba10e9d2cedc0a7f36f68ae50b8155ce042818d920def325e5624cfad9bc731ebea2624eee13f5893779f3a79125e7c17d8c944bf995218dc540941348eca39c0371e6e9899479e7020db985014a4d8fdaa22ac6931b840cec3a27110039a33e095196f6085741cb101e1350044aec892bff9918d2b015ed19e3f37b20222ce5fbd202f9ed089966aaa0c69b88413f6469b8f5fd248b21e301d798871ec954d29b9c0be79b69d55181d4f3f336edc39a2155b65c26e1c918db685e6671655fbaac671d628f2d40bf7c3688d98e7473d8dcc8efe8e328305f57e93e1a5a60f4a1b303b69b2a2f8a4565dc7b0c9d68433be61319965a2a3e95fbfe9e15846d803c111382f5cc052970d757632b13c631b3c5e43bef8ba11b61afc6b92f860656a9381e0787ee96987ca121d8fa4e87dbcd7516fe01ac182ce06f273e51f40f954d3f835757f2106e60531fb2b4eccf48b0f7e7d838eacb41426f1c4bdbca54d0aa05c661cc90be54e149266a861feaf8f17db9c12475d50dc8ce43a331db8592fa25699119f89ea34794b1979a2d33336daecc5cab9d903526781c40d0b81615fa82bc8ae6ac748ce77967c32978332ed2be73c3ff018f5808661bb54301f28196260ea183d5c448fa0977f2caabfb7ad22773dedd8bf04dfce36cdbaa39b5c5262800daed89eb37402234047ba6a1e492876e71f7897ac69a8f8cd7b24ec198691f31fec605d276f4b5ea7add1787c123302186181398f22e1a2dff3c73dd38134adcddd9826eefff74b1ecf4faf52a993f157e6e0d2cbf3d2742848f942fd480ecff0ef848dfb235acb1c1ae07718bf493ac8c9e10dd4114ea98734ff45cbf430a453a54127c3f40e4713292e3a2a849251fe5ae90779daf03293d7cab8db4e0710b19dc3192eea6576c39ea3508371e75fd212aab3be1f97f07a5ac5a1cff657b63fed97c2f19204b94d0cc357a69cff419c8c3009cee1943732d3ac88f061716bfcfd4fdf19ab854fbd5d763a21cc956e9153354b8ee712b3277a07611ce06698abe6c6a87f833e5cd0c68e016bf4ead9578d21ac53762e040e7ee772e50e6a84c6a91600436d622601ee95fa35f50307940a4fa29ef2f691f9ceffb8eccb2dad6a57094feb85bc3541e57d162b4171abb46901bcd4608174500051e5a5c600b1ea17f8ee3bc4c94188be74ec4fcfc71441542ad501b7e11fbb93f83ab59f6bd752bae996c309477e87b181f02b5b320907170518ce42904e49c1a0af4297379e351e8af9e81100dc36a6bed95339ac2d3eb89a859198243277f941e4039bcfe90971a716c0aa3b6d8885014b03ce9b7c22cf303f84e8afc96b6debc1296a1749d635cf8e6dbf0a1eccdcce06b7edd4cc5483a5ef07ba6b8c1ea9ed46876c4b6d8482f55ae53152df68a6315414155fbad17b7792eec29b6dfc4ae9a762d1a5506cf5b987db0bbd4e67c07cfb74a9cacc80d58c9a5ebcf710bb8cc37eaf56929db571f1d501d397ab436b4995a9a08a711198a75223e5157991f0f8c6ad25beddbc1bff2fbf53899e4bb1afb734dcfd4276d25e980ad9a773ae5d7931a141664b2bfcbd1f32039eb815792f7a9f95d4db3224bbe6a8739d3a43f5872b7ab803d937ce4a048f3524b7aca51a66ba7c2ef12a51519be5161d535b10b44e7ba59afa488039f9f96e09cbaed4eba4589b0e64f01a0c51acbf8188a3b0b6ff5029112f097c9ce86c003aa0271d63775cf51a6d57aafdd2113277f7b473f08510d7892071ada16a65b002894082eb674c65848e23285a8b8e48ad4985a32ce97080aa6a5b50a3a13296c58765b8e411636d69211993dcd74ed0dbc7a353f315dd3c5784b594fc13ef998dd92c32f7907e01f158cdb63e2aa3d03e4c5e71d075ae8e34e0e35b7efaa926e99a5a48a7b48dd001433cfb746c8b2ea54a2b0f47774aa2f891364b1977a0f8c6512a33630630f1aa3fae69bcf60eb4dd02e67bce1598e7c783cbcbc4eec9e466d4c903d14fd9d50cc95f92fc88c1a2e2ccf53d06f145a65d2e063dc5f29066602;
        #1
        $finish();
    end
endmodule
