module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    compressor_CLA486_16 compressor_CLA486_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA486_16(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [0:0] comp_out24;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [0:0] dst24);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [147:0] stage1_0;
   wire [134:0] stage1_1;
   wire [167:0] stage1_2;
   wire [243:0] stage1_3;
   wire [222:0] stage1_4;
   wire [336:0] stage1_5;
   wire [196:0] stage1_6;
   wire [216:0] stage1_7;
   wire [195:0] stage1_8;
   wire [210:0] stage1_9;
   wire [281:0] stage1_10;
   wire [213:0] stage1_11;
   wire [201:0] stage1_12;
   wire [234:0] stage1_13;
   wire [182:0] stage1_14;
   wire [154:0] stage1_15;
   wire [150:0] stage1_16;
   wire [80:0] stage1_17;
   wire [37:0] stage2_0;
   wire [62:0] stage2_1;
   wire [53:0] stage2_2;
   wire [85:0] stage2_3;
   wire [106:0] stage2_4;
   wire [107:0] stage2_5;
   wire [89:0] stage2_6;
   wire [102:0] stage2_7;
   wire [105:0] stage2_8;
   wire [80:0] stage2_9;
   wire [89:0] stage2_10;
   wire [106:0] stage2_11;
   wire [93:0] stage2_12;
   wire [85:0] stage2_13;
   wire [101:0] stage2_14;
   wire [74:0] stage2_15;
   wire [76:0] stage2_16;
   wire [95:0] stage2_17;
   wire [25:0] stage2_18;
   wire [4:0] stage2_19;
   wire [19:0] stage3_0;
   wire [14:0] stage3_1;
   wire [18:0] stage3_2;
   wire [40:0] stage3_3;
   wire [38:0] stage3_4;
   wire [39:0] stage3_5;
   wire [49:0] stage3_6;
   wire [35:0] stage3_7;
   wire [47:0] stage3_8;
   wire [42:0] stage3_9;
   wire [43:0] stage3_10;
   wire [37:0] stage3_11;
   wire [46:0] stage3_12;
   wire [39:0] stage3_13;
   wire [31:0] stage3_14;
   wire [43:0] stage3_15;
   wire [44:0] stage3_16;
   wire [29:0] stage3_17;
   wire [25:0] stage3_18;
   wire [18:0] stage3_19;
   wire [4:0] stage3_20;
   wire [0:0] stage3_21;
   wire [9:0] stage4_0;
   wire [5:0] stage4_1;
   wire [8:0] stage4_2;
   wire [9:0] stage4_3;
   wire [16:0] stage4_4;
   wire [14:0] stage4_5;
   wire [15:0] stage4_6;
   wire [20:0] stage4_7;
   wire [19:0] stage4_8;
   wire [15:0] stage4_9;
   wire [17:0] stage4_10;
   wire [18:0] stage4_11;
   wire [23:0] stage4_12;
   wire [16:0] stage4_13;
   wire [19:0] stage4_14;
   wire [27:0] stage4_15;
   wire [18:0] stage4_16;
   wire [12:0] stage4_17;
   wire [24:0] stage4_18;
   wire [13:0] stage4_19;
   wire [8:0] stage4_20;
   wire [2:0] stage4_21;
   wire [9:0] stage5_0;
   wire [5:0] stage5_1;
   wire [8:0] stage5_2;
   wire [5:0] stage5_3;
   wire [4:0] stage5_4;
   wire [3:0] stage5_5;
   wire [8:0] stage5_6;
   wire [8:0] stage5_7;
   wire [13:0] stage5_8;
   wire [8:0] stage5_9;
   wire [7:0] stage5_10;
   wire [6:0] stage5_11;
   wire [6:0] stage5_12;
   wire [9:0] stage5_13;
   wire [7:0] stage5_14;
   wire [9:0] stage5_15;
   wire [9:0] stage5_16;
   wire [7:0] stage5_17;
   wire [6:0] stage5_18;
   wire [10:0] stage5_19;
   wire [11:0] stage5_20;
   wire [3:0] stage5_21;
   wire [0:0] stage5_22;
   wire [5:0] stage6_0;
   wire [3:0] stage6_1;
   wire [4:0] stage6_2;
   wire [2:0] stage6_3;
   wire [5:0] stage6_4;
   wire [4:0] stage6_5;
   wire [2:0] stage6_6;
   wire [3:0] stage6_7;
   wire [3:0] stage6_8;
   wire [5:0] stage6_9;
   wire [4:0] stage6_10;
   wire [2:0] stage6_11;
   wire [1:0] stage6_12;
   wire [6:0] stage6_13;
   wire [3:0] stage6_14;
   wire [2:0] stage6_15;
   wire [5:0] stage6_16;
   wire [2:0] stage6_17;
   wire [5:0] stage6_18;
   wire [3:0] stage6_19;
   wire [4:0] stage6_20;
   wire [2:0] stage6_21;
   wire [2:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [0:0] stage7_24;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[12]},
      {stage0_3[24]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[13]},
      {stage0_3[25]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[14]},
      {stage0_3[26]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[15]},
      {stage0_3[27]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[16]},
      {stage0_3[28]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[17]},
      {stage0_3[29]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[18]},
      {stage0_3[30]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[19]},
      {stage0_3[31]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[20]},
      {stage0_3[32]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[21]},
      {stage0_3[33]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[22]},
      {stage0_3[34]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[23]},
      {stage0_3[35]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_2[24]},
      {stage0_3[36]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_2[25]},
      {stage0_3[37]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_2[26]},
      {stage0_3[38]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_2[27]},
      {stage0_3[39]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_2[28]},
      {stage0_3[40]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_2[29]},
      {stage0_3[41]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_2[30]},
      {stage0_3[42]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_2[31]},
      {stage0_3[43]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_2[32]},
      {stage0_3[44]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_2[33]},
      {stage0_3[45]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_2[34]},
      {stage0_3[46]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_2[35]},
      {stage0_3[47]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_2[36]},
      {stage0_3[48]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[255], stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[261], stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[267], stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[285], stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[291], stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[297], stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[315], stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[321], stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[327], stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338]},
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344]},
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246]},
      {stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[345], stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350]},
      {stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252]},
      {stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[351], stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356]},
      {stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258]},
      {stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[357], stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362]},
      {stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264]},
      {stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368]},
      {stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270]},
      {stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374]},
      {stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276]},
      {stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[375], stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380]},
      {stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282]},
      {stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[381], stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386]},
      {stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288]},
      {stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[387], stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392]},
      {stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294]},
      {stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398]},
      {stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300]},
      {stage1_4[80],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404]},
      {stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306]},
      {stage1_4[81],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[405], stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410]},
      {stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312]},
      {stage1_4[82],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[411], stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416]},
      {stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318]},
      {stage1_4[83],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[417], stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422]},
      {stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324]},
      {stage1_4[84],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[0],stage1_4[85],stage1_3[85],stage1_2[85],stage1_1[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[1],stage1_4[86],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[2],stage1_4[87],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[3],stage1_4[88],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[4],stage1_4[89],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[5],stage1_4[90],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[6],stage1_4[91],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage1_5[7],stage1_4[92],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102]},
      {stage1_5[8],stage1_4[93],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage1_5[9],stage1_4[94],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251]},
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage1_5[10],stage1_4[95],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257]},
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120]},
      {stage1_5[11],stage1_4[96],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263]},
      {stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126]},
      {stage1_5[12],stage1_4[97],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269]},
      {stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132]},
      {stage1_5[13],stage1_4[98],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275]},
      {stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage1_5[14],stage1_4[99],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281]},
      {stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage1_5[15],stage1_4[100],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287]},
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150]},
      {stage1_5[16],stage1_4[101],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293]},
      {stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage1_5[17],stage1_4[102],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299]},
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162]},
      {stage1_5[18],stage1_4[103],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305]},
      {stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage1_5[19],stage1_4[104],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311]},
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage1_5[20],stage1_4[105],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317]},
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180]},
      {stage1_5[21],stage1_4[106],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323]},
      {stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage1_5[22],stage1_4[107],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329]},
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192]},
      {stage1_5[23],stage1_4[108],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335]},
      {stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198]},
      {stage1_5[24],stage1_4[109],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341]},
      {stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage1_5[25],stage1_4[110],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347]},
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210]},
      {stage1_5[26],stage1_4[111],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353]},
      {stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage1_5[27],stage1_4[112],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359]},
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222]},
      {stage1_5[28],stage1_4[113],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365]},
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228]},
      {stage1_5[29],stage1_4[114],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage1_5[30],stage1_4[115],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377]},
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage1_5[31],stage1_4[116],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383]},
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage1_5[32],stage1_4[117],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389]},
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252]},
      {stage1_5[33],stage1_4[118],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395]},
      {stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258]},
      {stage1_5[34],stage1_4[119],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401]},
      {stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264]},
      {stage1_5[35],stage1_4[120],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407]},
      {stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270]},
      {stage1_5[36],stage1_4[121],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413]},
      {stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage1_5[37],stage1_4[122],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419]},
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282]},
      {stage1_5[38],stage1_4[123],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425]},
      {stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288]},
      {stage1_5[39],stage1_4[124],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431]},
      {stage0_3[289], stage0_3[290], stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294]},
      {stage1_5[40],stage1_4[125],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437]},
      {stage0_3[295], stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage1_5[41],stage1_4[126],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443]},
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage1_5[42],stage1_4[127],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449]},
      {stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312]},
      {stage1_5[43],stage1_4[128],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455]},
      {stage0_3[313], stage0_3[314], stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318]},
      {stage1_5[44],stage1_4[129],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461]},
      {stage0_3[319], stage0_3[320], stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324]},
      {stage1_5[45],stage1_4[130],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467]},
      {stage0_3[325], stage0_3[326], stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330]},
      {stage1_5[46],stage1_4[131],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473]},
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336]},
      {stage1_5[47],stage1_4[132],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479]},
      {stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342]},
      {stage1_5[48],stage1_4[133],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483], stage0_1[484], stage0_1[485]},
      {stage0_3[343], stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage1_5[49],stage1_4[134],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[50],stage1_4[135],stage1_3[135],stage1_2[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[51],stage1_4[136],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[52],stage1_4[137],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[53],stage1_4[138],stage1_3[138],stage1_2[138]}
   );
   gpc615_5 gpc139 (
      {stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_3[349]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[54],stage1_4[139],stage1_3[139],stage1_2[139]}
   );
   gpc615_5 gpc140 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358]},
      {stage0_3[350]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[55],stage1_4[140],stage1_3[140],stage1_2[140]}
   );
   gpc615_5 gpc141 (
      {stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363]},
      {stage0_3[351]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[56],stage1_4[141],stage1_3[141],stage1_2[141]}
   );
   gpc615_5 gpc142 (
      {stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage0_3[352]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[57],stage1_4[142],stage1_3[142],stage1_2[142]}
   );
   gpc615_5 gpc143 (
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373]},
      {stage0_3[353]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[58],stage1_4[143],stage1_3[143],stage1_2[143]}
   );
   gpc615_5 gpc144 (
      {stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378]},
      {stage0_3[354]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[59],stage1_4[144],stage1_3[144],stage1_2[144]}
   );
   gpc615_5 gpc145 (
      {stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_3[355]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[60],stage1_4[145],stage1_3[145],stage1_2[145]}
   );
   gpc615_5 gpc146 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388]},
      {stage0_3[356]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[61],stage1_4[146],stage1_3[146],stage1_2[146]}
   );
   gpc615_5 gpc147 (
      {stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393]},
      {stage0_3[357]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[62],stage1_4[147],stage1_3[147],stage1_2[147]}
   );
   gpc615_5 gpc148 (
      {stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398]},
      {stage0_3[358]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[63],stage1_4[148],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403]},
      {stage0_3[359]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[64],stage1_4[149],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408]},
      {stage0_3[360]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[65],stage1_4[150],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413]},
      {stage0_3[361]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[66],stage1_4[151],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418]},
      {stage0_3[362]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[67],stage1_4[152],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422], stage0_2[423]},
      {stage0_3[363]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[68],stage1_4[153],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427], stage0_2[428]},
      {stage0_3[364]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[69],stage1_4[154],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[429], stage0_2[430], stage0_2[431], stage0_2[432], stage0_2[433]},
      {stage0_3[365]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[70],stage1_4[155],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437], stage0_2[438]},
      {stage0_3[366]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[71],stage1_4[156],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442], stage0_2[443]},
      {stage0_3[367]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[72],stage1_4[157],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447], stage0_2[448]},
      {stage0_3[368]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[73],stage1_4[158],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_2[449], stage0_2[450], stage0_2[451], stage0_2[452], stage0_2[453]},
      {stage0_3[369]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[74],stage1_4[159],stage1_3[159],stage1_2[159]}
   );
   gpc615_5 gpc160 (
      {stage0_2[454], stage0_2[455], stage0_2[456], stage0_2[457], stage0_2[458]},
      {stage0_3[370]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[75],stage1_4[160],stage1_3[160],stage1_2[160]}
   );
   gpc615_5 gpc161 (
      {stage0_2[459], stage0_2[460], stage0_2[461], stage0_2[462], stage0_2[463]},
      {stage0_3[371]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[76],stage1_4[161],stage1_3[161],stage1_2[161]}
   );
   gpc615_5 gpc162 (
      {stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467], stage0_2[468]},
      {stage0_3[372]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[77],stage1_4[162],stage1_3[162],stage1_2[162]}
   );
   gpc615_5 gpc163 (
      {stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472], stage0_2[473]},
      {stage0_3[373]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[78],stage1_4[163],stage1_3[163],stage1_2[163]}
   );
   gpc615_5 gpc164 (
      {stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477], stage0_2[478]},
      {stage0_3[374]},
      {stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179]},
      {stage1_6[29],stage1_5[79],stage1_4[164],stage1_3[164],stage1_2[164]}
   );
   gpc615_5 gpc165 (
      {stage0_2[479], stage0_2[480], stage0_2[481], stage0_2[482], stage0_2[483]},
      {stage0_3[375]},
      {stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185]},
      {stage1_6[30],stage1_5[80],stage1_4[165],stage1_3[165],stage1_2[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[186]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[31],stage1_5[81],stage1_4[166],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[187]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[32],stage1_5[82],stage1_4[167],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[188]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[33],stage1_5[83],stage1_4[168],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[189]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[34],stage1_5[84],stage1_4[169],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[190]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[35],stage1_5[85],stage1_4[170],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[191]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[36],stage1_5[86],stage1_4[171],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[192]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[37],stage1_5[87],stage1_4[172],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[193]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[38],stage1_5[88],stage1_4[173],stage1_3[173]}
   );
   gpc606_5 gpc174 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[8],stage1_6[39],stage1_5[89],stage1_4[174]}
   );
   gpc606_5 gpc175 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[9],stage1_6[40],stage1_5[90],stage1_4[175]}
   );
   gpc606_5 gpc176 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[10],stage1_6[41],stage1_5[91],stage1_4[176]}
   );
   gpc606_5 gpc177 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[11],stage1_6[42],stage1_5[92],stage1_4[177]}
   );
   gpc606_5 gpc178 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[12],stage1_6[43],stage1_5[93],stage1_4[178]}
   );
   gpc606_5 gpc179 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[13],stage1_6[44],stage1_5[94],stage1_4[179]}
   );
   gpc606_5 gpc180 (
      {stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[14],stage1_6[45],stage1_5[95],stage1_4[180]}
   );
   gpc606_5 gpc181 (
      {stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[15],stage1_6[46],stage1_5[96],stage1_4[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[16],stage1_6[47],stage1_5[97],stage1_4[182]}
   );
   gpc606_5 gpc183 (
      {stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[17],stage1_6[48],stage1_5[98],stage1_4[183]}
   );
   gpc606_5 gpc184 (
      {stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[18],stage1_6[49],stage1_5[99],stage1_4[184]}
   );
   gpc606_5 gpc185 (
      {stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[19],stage1_6[50],stage1_5[100],stage1_4[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[20],stage1_6[51],stage1_5[101],stage1_4[186]}
   );
   gpc606_5 gpc187 (
      {stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[21],stage1_6[52],stage1_5[102],stage1_4[187]}
   );
   gpc606_5 gpc188 (
      {stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[22],stage1_6[53],stage1_5[103],stage1_4[188]}
   );
   gpc606_5 gpc189 (
      {stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[23],stage1_6[54],stage1_5[104],stage1_4[189]}
   );
   gpc606_5 gpc190 (
      {stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[24],stage1_6[55],stage1_5[105],stage1_4[190]}
   );
   gpc606_5 gpc191 (
      {stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[25],stage1_6[56],stage1_5[106],stage1_4[191]}
   );
   gpc606_5 gpc192 (
      {stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[26],stage1_6[57],stage1_5[107],stage1_4[192]}
   );
   gpc606_5 gpc193 (
      {stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[27],stage1_6[58],stage1_5[108],stage1_4[193]}
   );
   gpc606_5 gpc194 (
      {stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[28],stage1_6[59],stage1_5[109],stage1_4[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[29],stage1_6[60],stage1_5[110],stage1_4[195]}
   );
   gpc606_5 gpc196 (
      {stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[30],stage1_6[61],stage1_5[111],stage1_4[196]}
   );
   gpc606_5 gpc197 (
      {stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[31],stage1_6[62],stage1_5[112],stage1_4[197]}
   );
   gpc606_5 gpc198 (
      {stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[32],stage1_6[63],stage1_5[113],stage1_4[198]}
   );
   gpc606_5 gpc199 (
      {stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[33],stage1_6[64],stage1_5[114],stage1_4[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[34],stage1_6[65],stage1_5[115],stage1_4[200]}
   );
   gpc606_5 gpc201 (
      {stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[35],stage1_6[66],stage1_5[116],stage1_4[201]}
   );
   gpc606_5 gpc202 (
      {stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[36],stage1_6[67],stage1_5[117],stage1_4[202]}
   );
   gpc606_5 gpc203 (
      {stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[37],stage1_6[68],stage1_5[118],stage1_4[203]}
   );
   gpc606_5 gpc204 (
      {stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[38],stage1_6[69],stage1_5[119],stage1_4[204]}
   );
   gpc606_5 gpc205 (
      {stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[39],stage1_6[70],stage1_5[120],stage1_4[205]}
   );
   gpc606_5 gpc206 (
      {stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[40],stage1_6[71],stage1_5[121],stage1_4[206]}
   );
   gpc606_5 gpc207 (
      {stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[41],stage1_6[72],stage1_5[122],stage1_4[207]}
   );
   gpc606_5 gpc208 (
      {stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[42],stage1_6[73],stage1_5[123],stage1_4[208]}
   );
   gpc606_5 gpc209 (
      {stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[43],stage1_6[74],stage1_5[124],stage1_4[209]}
   );
   gpc606_5 gpc210 (
      {stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[44],stage1_6[75],stage1_5[125],stage1_4[210]}
   );
   gpc606_5 gpc211 (
      {stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[45],stage1_6[76],stage1_5[126],stage1_4[211]}
   );
   gpc606_5 gpc212 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[46],stage1_6[77],stage1_5[127],stage1_4[212]}
   );
   gpc606_5 gpc213 (
      {stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[47],stage1_6[78],stage1_5[128],stage1_4[213]}
   );
   gpc606_5 gpc214 (
      {stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[48],stage1_6[79],stage1_5[129],stage1_4[214]}
   );
   gpc606_5 gpc215 (
      {stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[49],stage1_6[80],stage1_5[130],stage1_4[215]}
   );
   gpc606_5 gpc216 (
      {stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[50],stage1_6[81],stage1_5[131],stage1_4[216]}
   );
   gpc606_5 gpc217 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[51],stage1_6[82],stage1_5[132],stage1_4[217]}
   );
   gpc606_5 gpc218 (
      {stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[52],stage1_6[83],stage1_5[133],stage1_4[218]}
   );
   gpc606_5 gpc219 (
      {stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[53],stage1_6[84],stage1_5[134],stage1_4[219]}
   );
   gpc606_5 gpc220 (
      {stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[54],stage1_6[85],stage1_5[135],stage1_4[220]}
   );
   gpc615_5 gpc221 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_5[48]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[55],stage1_6[86],stage1_5[136],stage1_4[221]}
   );
   gpc615_5 gpc222 (
      {stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485]},
      {stage0_5[49]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[56],stage1_6[87],stage1_5[137],stage1_4[222]}
   );
   gpc606_5 gpc223 (
      {stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[49],stage1_7[57],stage1_6[88],stage1_5[138]}
   );
   gpc606_5 gpc224 (
      {stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[50],stage1_7[58],stage1_6[89],stage1_5[139]}
   );
   gpc606_5 gpc225 (
      {stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[51],stage1_7[59],stage1_6[90],stage1_5[140]}
   );
   gpc606_5 gpc226 (
      {stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72], stage0_5[73]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[52],stage1_7[60],stage1_6[91],stage1_5[141]}
   );
   gpc606_5 gpc227 (
      {stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78], stage0_5[79]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[53],stage1_7[61],stage1_6[92],stage1_5[142]}
   );
   gpc606_5 gpc228 (
      {stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[54],stage1_7[62],stage1_6[93],stage1_5[143]}
   );
   gpc606_5 gpc229 (
      {stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[55],stage1_7[63],stage1_6[94],stage1_5[144]}
   );
   gpc606_5 gpc230 (
      {stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[56],stage1_7[64],stage1_6[95],stage1_5[145]}
   );
   gpc606_5 gpc231 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[57],stage1_7[65],stage1_6[96],stage1_5[146]}
   );
   gpc606_5 gpc232 (
      {stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[58],stage1_7[66],stage1_6[97],stage1_5[147]}
   );
   gpc606_5 gpc233 (
      {stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[59],stage1_7[67],stage1_6[98],stage1_5[148]}
   );
   gpc606_5 gpc234 (
      {stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[60],stage1_7[68],stage1_6[99],stage1_5[149]}
   );
   gpc606_5 gpc235 (
      {stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[61],stage1_7[69],stage1_6[100],stage1_5[150]}
   );
   gpc606_5 gpc236 (
      {stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132], stage0_5[133]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[62],stage1_7[70],stage1_6[101],stage1_5[151]}
   );
   gpc606_5 gpc237 (
      {stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138], stage0_5[139]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[63],stage1_7[71],stage1_6[102],stage1_5[152]}
   );
   gpc606_5 gpc238 (
      {stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[64],stage1_7[72],stage1_6[103],stage1_5[153]}
   );
   gpc606_5 gpc239 (
      {stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[65],stage1_7[73],stage1_6[104],stage1_5[154]}
   );
   gpc606_5 gpc240 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[66],stage1_7[74],stage1_6[105],stage1_5[155]}
   );
   gpc606_5 gpc241 (
      {stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[67],stage1_7[75],stage1_6[106],stage1_5[156]}
   );
   gpc606_5 gpc242 (
      {stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[68],stage1_7[76],stage1_6[107],stage1_5[157]}
   );
   gpc606_5 gpc243 (
      {stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[69],stage1_7[77],stage1_6[108],stage1_5[158]}
   );
   gpc606_5 gpc244 (
      {stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[70],stage1_7[78],stage1_6[109],stage1_5[159]}
   );
   gpc606_5 gpc245 (
      {stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[71],stage1_7[79],stage1_6[110],stage1_5[160]}
   );
   gpc606_5 gpc246 (
      {stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[72],stage1_7[80],stage1_6[111],stage1_5[161]}
   );
   gpc606_5 gpc247 (
      {stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[73],stage1_7[81],stage1_6[112],stage1_5[162]}
   );
   gpc606_5 gpc248 (
      {stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[74],stage1_7[82],stage1_6[113],stage1_5[163]}
   );
   gpc606_5 gpc249 (
      {stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[75],stage1_7[83],stage1_6[114],stage1_5[164]}
   );
   gpc606_5 gpc250 (
      {stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[76],stage1_7[84],stage1_6[115],stage1_5[165]}
   );
   gpc606_5 gpc251 (
      {stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[77],stage1_7[85],stage1_6[116],stage1_5[166]}
   );
   gpc606_5 gpc252 (
      {stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[78],stage1_7[86],stage1_6[117],stage1_5[167]}
   );
   gpc606_5 gpc253 (
      {stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[79],stage1_7[87],stage1_6[118],stage1_5[168]}
   );
   gpc606_5 gpc254 (
      {stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[80],stage1_7[88],stage1_6[119],stage1_5[169]}
   );
   gpc606_5 gpc255 (
      {stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[81],stage1_7[89],stage1_6[120],stage1_5[170]}
   );
   gpc606_5 gpc256 (
      {stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[82],stage1_7[90],stage1_6[121],stage1_5[171]}
   );
   gpc606_5 gpc257 (
      {stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258], stage0_5[259]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[83],stage1_7[91],stage1_6[122],stage1_5[172]}
   );
   gpc606_5 gpc258 (
      {stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264], stage0_5[265]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[84],stage1_7[92],stage1_6[123],stage1_5[173]}
   );
   gpc606_5 gpc259 (
      {stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270], stage0_5[271]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[85],stage1_7[93],stage1_6[124],stage1_5[174]}
   );
   gpc615_5 gpc260 (
      {stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276]},
      {stage0_6[294]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[86],stage1_7[94],stage1_6[125],stage1_5[175]}
   );
   gpc615_5 gpc261 (
      {stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_6[295]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[87],stage1_7[95],stage1_6[126],stage1_5[176]}
   );
   gpc615_5 gpc262 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286]},
      {stage0_6[296]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[88],stage1_7[96],stage1_6[127],stage1_5[177]}
   );
   gpc615_5 gpc263 (
      {stage0_5[287], stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291]},
      {stage0_6[297]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[89],stage1_7[97],stage1_6[128],stage1_5[178]}
   );
   gpc615_5 gpc264 (
      {stage0_5[292], stage0_5[293], stage0_5[294], stage0_5[295], stage0_5[296]},
      {stage0_6[298]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[90],stage1_7[98],stage1_6[129],stage1_5[179]}
   );
   gpc615_5 gpc265 (
      {stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300], stage0_5[301]},
      {stage0_6[299]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[91],stage1_7[99],stage1_6[130],stage1_5[180]}
   );
   gpc615_5 gpc266 (
      {stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306]},
      {stage0_6[300]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[92],stage1_7[100],stage1_6[131],stage1_5[181]}
   );
   gpc615_5 gpc267 (
      {stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_6[301]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[93],stage1_7[101],stage1_6[132],stage1_5[182]}
   );
   gpc615_5 gpc268 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316]},
      {stage0_6[302]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[94],stage1_7[102],stage1_6[133],stage1_5[183]}
   );
   gpc615_5 gpc269 (
      {stage0_5[317], stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321]},
      {stage0_6[303]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[95],stage1_7[103],stage1_6[134],stage1_5[184]}
   );
   gpc615_5 gpc270 (
      {stage0_5[322], stage0_5[323], stage0_5[324], stage0_5[325], stage0_5[326]},
      {stage0_6[304]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[96],stage1_7[104],stage1_6[135],stage1_5[185]}
   );
   gpc615_5 gpc271 (
      {stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330], stage0_5[331]},
      {stage0_6[305]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[97],stage1_7[105],stage1_6[136],stage1_5[186]}
   );
   gpc615_5 gpc272 (
      {stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336]},
      {stage0_6[306]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[98],stage1_7[106],stage1_6[137],stage1_5[187]}
   );
   gpc615_5 gpc273 (
      {stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage0_7[300]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[50],stage1_8[99],stage1_7[107],stage1_6[138]}
   );
   gpc615_5 gpc274 (
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316]},
      {stage0_7[301]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[51],stage1_8[100],stage1_7[108],stage1_6[139]}
   );
   gpc615_5 gpc275 (
      {stage0_6[317], stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321]},
      {stage0_7[302]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[52],stage1_8[101],stage1_7[109],stage1_6[140]}
   );
   gpc615_5 gpc276 (
      {stage0_6[322], stage0_6[323], stage0_6[324], stage0_6[325], stage0_6[326]},
      {stage0_7[303]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[53],stage1_8[102],stage1_7[110],stage1_6[141]}
   );
   gpc615_5 gpc277 (
      {stage0_6[327], stage0_6[328], stage0_6[329], stage0_6[330], stage0_6[331]},
      {stage0_7[304]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[54],stage1_8[103],stage1_7[111],stage1_6[142]}
   );
   gpc615_5 gpc278 (
      {stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335], stage0_6[336]},
      {stage0_7[305]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[55],stage1_8[104],stage1_7[112],stage1_6[143]}
   );
   gpc615_5 gpc279 (
      {stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage0_7[306]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[56],stage1_8[105],stage1_7[113],stage1_6[144]}
   );
   gpc615_5 gpc280 (
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346]},
      {stage0_7[307]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[57],stage1_8[106],stage1_7[114],stage1_6[145]}
   );
   gpc615_5 gpc281 (
      {stage0_6[347], stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351]},
      {stage0_7[308]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[58],stage1_8[107],stage1_7[115],stage1_6[146]}
   );
   gpc615_5 gpc282 (
      {stage0_6[352], stage0_6[353], stage0_6[354], stage0_6[355], stage0_6[356]},
      {stage0_7[309]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[59],stage1_8[108],stage1_7[116],stage1_6[147]}
   );
   gpc615_5 gpc283 (
      {stage0_6[357], stage0_6[358], stage0_6[359], stage0_6[360], stage0_6[361]},
      {stage0_7[310]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[60],stage1_8[109],stage1_7[117],stage1_6[148]}
   );
   gpc615_5 gpc284 (
      {stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365], stage0_6[366]},
      {stage0_7[311]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[61],stage1_8[110],stage1_7[118],stage1_6[149]}
   );
   gpc615_5 gpc285 (
      {stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage0_7[312]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[62],stage1_8[111],stage1_7[119],stage1_6[150]}
   );
   gpc615_5 gpc286 (
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376]},
      {stage0_7[313]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[63],stage1_8[112],stage1_7[120],stage1_6[151]}
   );
   gpc615_5 gpc287 (
      {stage0_6[377], stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381]},
      {stage0_7[314]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[64],stage1_8[113],stage1_7[121],stage1_6[152]}
   );
   gpc615_5 gpc288 (
      {stage0_6[382], stage0_6[383], stage0_6[384], stage0_6[385], stage0_6[386]},
      {stage0_7[315]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[65],stage1_8[114],stage1_7[122],stage1_6[153]}
   );
   gpc615_5 gpc289 (
      {stage0_6[387], stage0_6[388], stage0_6[389], stage0_6[390], stage0_6[391]},
      {stage0_7[316]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[66],stage1_8[115],stage1_7[123],stage1_6[154]}
   );
   gpc615_5 gpc290 (
      {stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395], stage0_6[396]},
      {stage0_7[317]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[67],stage1_8[116],stage1_7[124],stage1_6[155]}
   );
   gpc615_5 gpc291 (
      {stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage0_7[318]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[68],stage1_8[117],stage1_7[125],stage1_6[156]}
   );
   gpc615_5 gpc292 (
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406]},
      {stage0_7[319]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[69],stage1_8[118],stage1_7[126],stage1_6[157]}
   );
   gpc615_5 gpc293 (
      {stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411]},
      {stage0_7[320]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[70],stage1_8[119],stage1_7[127],stage1_6[158]}
   );
   gpc615_5 gpc294 (
      {stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415], stage0_6[416]},
      {stage0_7[321]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[71],stage1_8[120],stage1_7[128],stage1_6[159]}
   );
   gpc615_5 gpc295 (
      {stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420], stage0_6[421]},
      {stage0_7[322]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[72],stage1_8[121],stage1_7[129],stage1_6[160]}
   );
   gpc615_5 gpc296 (
      {stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425], stage0_6[426]},
      {stage0_7[323]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[73],stage1_8[122],stage1_7[130],stage1_6[161]}
   );
   gpc615_5 gpc297 (
      {stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage0_7[324]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[74],stage1_8[123],stage1_7[131],stage1_6[162]}
   );
   gpc615_5 gpc298 (
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436]},
      {stage0_7[325]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[75],stage1_8[124],stage1_7[132],stage1_6[163]}
   );
   gpc615_5 gpc299 (
      {stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441]},
      {stage0_7[326]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[76],stage1_8[125],stage1_7[133],stage1_6[164]}
   );
   gpc615_5 gpc300 (
      {stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445], stage0_6[446]},
      {stage0_7[327]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[77],stage1_8[126],stage1_7[134],stage1_6[165]}
   );
   gpc615_5 gpc301 (
      {stage0_6[447], stage0_6[448], stage0_6[449], stage0_6[450], stage0_6[451]},
      {stage0_7[328]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[78],stage1_8[127],stage1_7[135],stage1_6[166]}
   );
   gpc615_5 gpc302 (
      {stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455], stage0_6[456]},
      {stage0_7[329]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[79],stage1_8[128],stage1_7[136],stage1_6[167]}
   );
   gpc615_5 gpc303 (
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334]},
      {stage0_8[180]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[30],stage1_9[80],stage1_8[129],stage1_7[137]}
   );
   gpc615_5 gpc304 (
      {stage0_7[335], stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339]},
      {stage0_8[181]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[31],stage1_9[81],stage1_8[130],stage1_7[138]}
   );
   gpc615_5 gpc305 (
      {stage0_7[340], stage0_7[341], stage0_7[342], stage0_7[343], stage0_7[344]},
      {stage0_8[182]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[32],stage1_9[82],stage1_8[131],stage1_7[139]}
   );
   gpc615_5 gpc306 (
      {stage0_7[345], stage0_7[346], stage0_7[347], stage0_7[348], stage0_7[349]},
      {stage0_8[183]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[33],stage1_9[83],stage1_8[132],stage1_7[140]}
   );
   gpc615_5 gpc307 (
      {stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353], stage0_7[354]},
      {stage0_8[184]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[34],stage1_9[84],stage1_8[133],stage1_7[141]}
   );
   gpc615_5 gpc308 (
      {stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage0_8[185]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[35],stage1_9[85],stage1_8[134],stage1_7[142]}
   );
   gpc615_5 gpc309 (
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364]},
      {stage0_8[186]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[36],stage1_9[86],stage1_8[135],stage1_7[143]}
   );
   gpc615_5 gpc310 (
      {stage0_7[365], stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369]},
      {stage0_8[187]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[37],stage1_9[87],stage1_8[136],stage1_7[144]}
   );
   gpc615_5 gpc311 (
      {stage0_7[370], stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374]},
      {stage0_8[188]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[38],stage1_9[88],stage1_8[137],stage1_7[145]}
   );
   gpc615_5 gpc312 (
      {stage0_7[375], stage0_7[376], stage0_7[377], stage0_7[378], stage0_7[379]},
      {stage0_8[189]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[39],stage1_9[89],stage1_8[138],stage1_7[146]}
   );
   gpc615_5 gpc313 (
      {stage0_7[380], stage0_7[381], stage0_7[382], stage0_7[383], stage0_7[384]},
      {stage0_8[190]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[40],stage1_9[90],stage1_8[139],stage1_7[147]}
   );
   gpc615_5 gpc314 (
      {stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389]},
      {stage0_8[191]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[41],stage1_9[91],stage1_8[140],stage1_7[148]}
   );
   gpc615_5 gpc315 (
      {stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394]},
      {stage0_8[192]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[42],stage1_9[92],stage1_8[141],stage1_7[149]}
   );
   gpc615_5 gpc316 (
      {stage0_7[395], stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399]},
      {stage0_8[193]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[43],stage1_9[93],stage1_8[142],stage1_7[150]}
   );
   gpc615_5 gpc317 (
      {stage0_7[400], stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404]},
      {stage0_8[194]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[44],stage1_9[94],stage1_8[143],stage1_7[151]}
   );
   gpc615_5 gpc318 (
      {stage0_7[405], stage0_7[406], stage0_7[407], stage0_7[408], stage0_7[409]},
      {stage0_8[195]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[45],stage1_9[95],stage1_8[144],stage1_7[152]}
   );
   gpc615_5 gpc319 (
      {stage0_7[410], stage0_7[411], stage0_7[412], stage0_7[413], stage0_7[414]},
      {stage0_8[196]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[46],stage1_9[96],stage1_8[145],stage1_7[153]}
   );
   gpc615_5 gpc320 (
      {stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419]},
      {stage0_8[197]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[47],stage1_9[97],stage1_8[146],stage1_7[154]}
   );
   gpc615_5 gpc321 (
      {stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424]},
      {stage0_8[198]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[48],stage1_9[98],stage1_8[147],stage1_7[155]}
   );
   gpc606_5 gpc322 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[19],stage1_10[49],stage1_9[99],stage1_8[148]}
   );
   gpc606_5 gpc323 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[20],stage1_10[50],stage1_9[100],stage1_8[149]}
   );
   gpc606_5 gpc324 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[21],stage1_10[51],stage1_9[101],stage1_8[150]}
   );
   gpc606_5 gpc325 (
      {stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[22],stage1_10[52],stage1_9[102],stage1_8[151]}
   );
   gpc606_5 gpc326 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[23],stage1_10[53],stage1_9[103],stage1_8[152]}
   );
   gpc606_5 gpc327 (
      {stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[24],stage1_10[54],stage1_9[104],stage1_8[153]}
   );
   gpc606_5 gpc328 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[25],stage1_10[55],stage1_9[105],stage1_8[154]}
   );
   gpc606_5 gpc329 (
      {stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[26],stage1_10[56],stage1_9[106],stage1_8[155]}
   );
   gpc606_5 gpc330 (
      {stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[27],stage1_10[57],stage1_9[107],stage1_8[156]}
   );
   gpc606_5 gpc331 (
      {stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[28],stage1_10[58],stage1_9[108],stage1_8[157]}
   );
   gpc606_5 gpc332 (
      {stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[29],stage1_10[59],stage1_9[109],stage1_8[158]}
   );
   gpc606_5 gpc333 (
      {stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[30],stage1_10[60],stage1_9[110],stage1_8[159]}
   );
   gpc606_5 gpc334 (
      {stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[31],stage1_10[61],stage1_9[111],stage1_8[160]}
   );
   gpc606_5 gpc335 (
      {stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[32],stage1_10[62],stage1_9[112],stage1_8[161]}
   );
   gpc606_5 gpc336 (
      {stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[33],stage1_10[63],stage1_9[113],stage1_8[162]}
   );
   gpc606_5 gpc337 (
      {stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[34],stage1_10[64],stage1_9[114],stage1_8[163]}
   );
   gpc606_5 gpc338 (
      {stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[35],stage1_10[65],stage1_9[115],stage1_8[164]}
   );
   gpc606_5 gpc339 (
      {stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[36],stage1_10[66],stage1_9[116],stage1_8[165]}
   );
   gpc606_5 gpc340 (
      {stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[37],stage1_10[67],stage1_9[117],stage1_8[166]}
   );
   gpc606_5 gpc341 (
      {stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[38],stage1_10[68],stage1_9[118],stage1_8[167]}
   );
   gpc606_5 gpc342 (
      {stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[39],stage1_10[69],stage1_9[119],stage1_8[168]}
   );
   gpc606_5 gpc343 (
      {stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[40],stage1_10[70],stage1_9[120],stage1_8[169]}
   );
   gpc606_5 gpc344 (
      {stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[41],stage1_10[71],stage1_9[121],stage1_8[170]}
   );
   gpc606_5 gpc345 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[42],stage1_10[72],stage1_9[122],stage1_8[171]}
   );
   gpc606_5 gpc346 (
      {stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[43],stage1_10[73],stage1_9[123],stage1_8[172]}
   );
   gpc606_5 gpc347 (
      {stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[44],stage1_10[74],stage1_9[124],stage1_8[173]}
   );
   gpc606_5 gpc348 (
      {stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[45],stage1_10[75],stage1_9[125],stage1_8[174]}
   );
   gpc606_5 gpc349 (
      {stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[46],stage1_10[76],stage1_9[126],stage1_8[175]}
   );
   gpc606_5 gpc350 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[47],stage1_10[77],stage1_9[127],stage1_8[176]}
   );
   gpc606_5 gpc351 (
      {stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[48],stage1_10[78],stage1_9[128],stage1_8[177]}
   );
   gpc606_5 gpc352 (
      {stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[49],stage1_10[79],stage1_9[129],stage1_8[178]}
   );
   gpc606_5 gpc353 (
      {stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[50],stage1_10[80],stage1_9[130],stage1_8[179]}
   );
   gpc606_5 gpc354 (
      {stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[51],stage1_10[81],stage1_9[131],stage1_8[180]}
   );
   gpc606_5 gpc355 (
      {stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[52],stage1_10[82],stage1_9[132],stage1_8[181]}
   );
   gpc606_5 gpc356 (
      {stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[53],stage1_10[83],stage1_9[133],stage1_8[182]}
   );
   gpc606_5 gpc357 (
      {stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[54],stage1_10[84],stage1_9[134],stage1_8[183]}
   );
   gpc606_5 gpc358 (
      {stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[55],stage1_10[85],stage1_9[135],stage1_8[184]}
   );
   gpc606_5 gpc359 (
      {stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[56],stage1_10[86],stage1_9[136],stage1_8[185]}
   );
   gpc606_5 gpc360 (
      {stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[57],stage1_10[87],stage1_9[137],stage1_8[186]}
   );
   gpc606_5 gpc361 (
      {stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[58],stage1_10[88],stage1_9[138],stage1_8[187]}
   );
   gpc606_5 gpc362 (
      {stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[59],stage1_10[89],stage1_9[139],stage1_8[188]}
   );
   gpc606_5 gpc363 (
      {stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[60],stage1_10[90],stage1_9[140],stage1_8[189]}
   );
   gpc606_5 gpc364 (
      {stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[61],stage1_10[91],stage1_9[141],stage1_8[190]}
   );
   gpc606_5 gpc365 (
      {stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[62],stage1_10[92],stage1_9[142],stage1_8[191]}
   );
   gpc606_5 gpc366 (
      {stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[63],stage1_10[93],stage1_9[143],stage1_8[192]}
   );
   gpc606_5 gpc367 (
      {stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[64],stage1_10[94],stage1_9[144],stage1_8[193]}
   );
   gpc606_5 gpc368 (
      {stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[65],stage1_10[95],stage1_9[145],stage1_8[194]}
   );
   gpc615_5 gpc369 (
      {stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_9[114]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[66],stage1_10[96],stage1_9[146],stage1_8[195]}
   );
   gpc606_5 gpc370 (
      {stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[48],stage1_11[67],stage1_10[97],stage1_9[147]}
   );
   gpc606_5 gpc371 (
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[49],stage1_11[68],stage1_10[98],stage1_9[148]}
   );
   gpc606_5 gpc372 (
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[50],stage1_11[69],stage1_10[99],stage1_9[149]}
   );
   gpc606_5 gpc373 (
      {stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[51],stage1_11[70],stage1_10[100],stage1_9[150]}
   );
   gpc606_5 gpc374 (
      {stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[52],stage1_11[71],stage1_10[101],stage1_9[151]}
   );
   gpc606_5 gpc375 (
      {stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[53],stage1_11[72],stage1_10[102],stage1_9[152]}
   );
   gpc606_5 gpc376 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[54],stage1_11[73],stage1_10[103],stage1_9[153]}
   );
   gpc606_5 gpc377 (
      {stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161], stage0_9[162]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[55],stage1_11[74],stage1_10[104],stage1_9[154]}
   );
   gpc606_5 gpc378 (
      {stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[56],stage1_11[75],stage1_10[105],stage1_9[155]}
   );
   gpc606_5 gpc379 (
      {stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[57],stage1_11[76],stage1_10[106],stage1_9[156]}
   );
   gpc606_5 gpc380 (
      {stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[58],stage1_11[77],stage1_10[107],stage1_9[157]}
   );
   gpc606_5 gpc381 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185], stage0_9[186]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[59],stage1_11[78],stage1_10[108],stage1_9[158]}
   );
   gpc606_5 gpc382 (
      {stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191], stage0_9[192]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[60],stage1_11[79],stage1_10[109],stage1_9[159]}
   );
   gpc606_5 gpc383 (
      {stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[61],stage1_11[80],stage1_10[110],stage1_9[160]}
   );
   gpc606_5 gpc384 (
      {stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[62],stage1_11[81],stage1_10[111],stage1_9[161]}
   );
   gpc606_5 gpc385 (
      {stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[63],stage1_11[82],stage1_10[112],stage1_9[162]}
   );
   gpc606_5 gpc386 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215], stage0_9[216]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[64],stage1_11[83],stage1_10[113],stage1_9[163]}
   );
   gpc606_5 gpc387 (
      {stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221], stage0_9[222]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[65],stage1_11[84],stage1_10[114],stage1_9[164]}
   );
   gpc606_5 gpc388 (
      {stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[66],stage1_11[85],stage1_10[115],stage1_9[165]}
   );
   gpc606_5 gpc389 (
      {stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[67],stage1_11[86],stage1_10[116],stage1_9[166]}
   );
   gpc606_5 gpc390 (
      {stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[68],stage1_11[87],stage1_10[117],stage1_9[167]}
   );
   gpc606_5 gpc391 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245], stage0_9[246]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[69],stage1_11[88],stage1_10[118],stage1_9[168]}
   );
   gpc606_5 gpc392 (
      {stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251], stage0_9[252]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[70],stage1_11[89],stage1_10[119],stage1_9[169]}
   );
   gpc606_5 gpc393 (
      {stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257], stage0_9[258]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[71],stage1_11[90],stage1_10[120],stage1_9[170]}
   );
   gpc606_5 gpc394 (
      {stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[72],stage1_11[91],stage1_10[121],stage1_9[171]}
   );
   gpc606_5 gpc395 (
      {stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[73],stage1_11[92],stage1_10[122],stage1_9[172]}
   );
   gpc606_5 gpc396 (
      {stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275], stage0_9[276]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[74],stage1_11[93],stage1_10[123],stage1_9[173]}
   );
   gpc606_5 gpc397 (
      {stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281], stage0_9[282]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[75],stage1_11[94],stage1_10[124],stage1_9[174]}
   );
   gpc606_5 gpc398 (
      {stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287], stage0_9[288]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[76],stage1_11[95],stage1_10[125],stage1_9[175]}
   );
   gpc606_5 gpc399 (
      {stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[77],stage1_11[96],stage1_10[126],stage1_9[176]}
   );
   gpc606_5 gpc400 (
      {stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[78],stage1_11[97],stage1_10[127],stage1_9[177]}
   );
   gpc606_5 gpc401 (
      {stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305], stage0_9[306]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[79],stage1_11[98],stage1_10[128],stage1_9[178]}
   );
   gpc606_5 gpc402 (
      {stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311], stage0_9[312]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[80],stage1_11[99],stage1_10[129],stage1_9[179]}
   );
   gpc606_5 gpc403 (
      {stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317], stage0_9[318]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[81],stage1_11[100],stage1_10[130],stage1_9[180]}
   );
   gpc606_5 gpc404 (
      {stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[82],stage1_11[101],stage1_10[131],stage1_9[181]}
   );
   gpc606_5 gpc405 (
      {stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[83],stage1_11[102],stage1_10[132],stage1_9[182]}
   );
   gpc606_5 gpc406 (
      {stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335], stage0_9[336]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[84],stage1_11[103],stage1_10[133],stage1_9[183]}
   );
   gpc606_5 gpc407 (
      {stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341], stage0_9[342]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[85],stage1_11[104],stage1_10[134],stage1_9[184]}
   );
   gpc606_5 gpc408 (
      {stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347], stage0_9[348]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[86],stage1_11[105],stage1_10[135],stage1_9[185]}
   );
   gpc606_5 gpc409 (
      {stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[87],stage1_11[106],stage1_10[136],stage1_9[186]}
   );
   gpc606_5 gpc410 (
      {stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[88],stage1_11[107],stage1_10[137],stage1_9[187]}
   );
   gpc606_5 gpc411 (
      {stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365], stage0_9[366]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[89],stage1_11[108],stage1_10[138],stage1_9[188]}
   );
   gpc606_5 gpc412 (
      {stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371], stage0_9[372]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[90],stage1_11[109],stage1_10[139],stage1_9[189]}
   );
   gpc606_5 gpc413 (
      {stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377], stage0_9[378]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[91],stage1_11[110],stage1_10[140],stage1_9[190]}
   );
   gpc606_5 gpc414 (
      {stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[92],stage1_11[111],stage1_10[141],stage1_9[191]}
   );
   gpc606_5 gpc415 (
      {stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[93],stage1_11[112],stage1_10[142],stage1_9[192]}
   );
   gpc606_5 gpc416 (
      {stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395], stage0_9[396]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[94],stage1_11[113],stage1_10[143],stage1_9[193]}
   );
   gpc606_5 gpc417 (
      {stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401], stage0_9[402]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[95],stage1_11[114],stage1_10[144],stage1_9[194]}
   );
   gpc606_5 gpc418 (
      {stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407], stage0_9[408]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[96],stage1_11[115],stage1_10[145],stage1_9[195]}
   );
   gpc606_5 gpc419 (
      {stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413], stage0_9[414]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[97],stage1_11[116],stage1_10[146],stage1_9[196]}
   );
   gpc606_5 gpc420 (
      {stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419], stage0_9[420]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[98],stage1_11[117],stage1_10[147],stage1_9[197]}
   );
   gpc615_5 gpc421 (
      {stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_10[288]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[99],stage1_11[118],stage1_10[148],stage1_9[198]}
   );
   gpc615_5 gpc422 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430]},
      {stage0_10[289]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[100],stage1_11[119],stage1_10[149],stage1_9[199]}
   );
   gpc615_5 gpc423 (
      {stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_10[290]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[101],stage1_11[120],stage1_10[150],stage1_9[200]}
   );
   gpc615_5 gpc424 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440]},
      {stage0_10[291]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[102],stage1_11[121],stage1_10[151],stage1_9[201]}
   );
   gpc615_5 gpc425 (
      {stage0_9[441], stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445]},
      {stage0_10[292]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[103],stage1_11[122],stage1_10[152],stage1_9[202]}
   );
   gpc615_5 gpc426 (
      {stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449], stage0_9[450]},
      {stage0_10[293]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[104],stage1_11[123],stage1_10[153],stage1_9[203]}
   );
   gpc615_5 gpc427 (
      {stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_10[294]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[105],stage1_11[124],stage1_10[154],stage1_9[204]}
   );
   gpc615_5 gpc428 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460]},
      {stage0_10[295]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[106],stage1_11[125],stage1_10[155],stage1_9[205]}
   );
   gpc615_5 gpc429 (
      {stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_10[296]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[107],stage1_11[126],stage1_10[156],stage1_9[206]}
   );
   gpc615_5 gpc430 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470]},
      {stage0_10[297]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[108],stage1_11[127],stage1_10[157],stage1_9[207]}
   );
   gpc615_5 gpc431 (
      {stage0_9[471], stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475]},
      {stage0_10[298]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[109],stage1_11[128],stage1_10[158],stage1_9[208]}
   );
   gpc615_5 gpc432 (
      {stage0_9[476], stage0_9[477], stage0_9[478], stage0_9[479], stage0_9[480]},
      {stage0_10[299]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[110],stage1_11[129],stage1_10[159],stage1_9[209]}
   );
   gpc615_5 gpc433 (
      {stage0_9[481], stage0_9[482], stage0_9[483], stage0_9[484], stage0_9[485]},
      {stage0_10[300]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[111],stage1_11[130],stage1_10[160],stage1_9[210]}
   );
   gpc615_5 gpc434 (
      {stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage0_11[384]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[64],stage1_12[112],stage1_11[131],stage1_10[161]}
   );
   gpc615_5 gpc435 (
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310]},
      {stage0_11[385]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[65],stage1_12[113],stage1_11[132],stage1_10[162]}
   );
   gpc615_5 gpc436 (
      {stage0_10[311], stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315]},
      {stage0_11[386]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[66],stage1_12[114],stage1_11[133],stage1_10[163]}
   );
   gpc615_5 gpc437 (
      {stage0_10[316], stage0_10[317], stage0_10[318], stage0_10[319], stage0_10[320]},
      {stage0_11[387]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[67],stage1_12[115],stage1_11[134],stage1_10[164]}
   );
   gpc615_5 gpc438 (
      {stage0_10[321], stage0_10[322], stage0_10[323], stage0_10[324], stage0_10[325]},
      {stage0_11[388]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[68],stage1_12[116],stage1_11[135],stage1_10[165]}
   );
   gpc615_5 gpc439 (
      {stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329], stage0_10[330]},
      {stage0_11[389]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[69],stage1_12[117],stage1_11[136],stage1_10[166]}
   );
   gpc615_5 gpc440 (
      {stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage0_11[390]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[70],stage1_12[118],stage1_11[137],stage1_10[167]}
   );
   gpc615_5 gpc441 (
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340]},
      {stage0_11[391]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[71],stage1_12[119],stage1_11[138],stage1_10[168]}
   );
   gpc615_5 gpc442 (
      {stage0_10[341], stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345]},
      {stage0_11[392]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[72],stage1_12[120],stage1_11[139],stage1_10[169]}
   );
   gpc615_5 gpc443 (
      {stage0_10[346], stage0_10[347], stage0_10[348], stage0_10[349], stage0_10[350]},
      {stage0_11[393]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[73],stage1_12[121],stage1_11[140],stage1_10[170]}
   );
   gpc615_5 gpc444 (
      {stage0_10[351], stage0_10[352], stage0_10[353], stage0_10[354], stage0_10[355]},
      {stage0_11[394]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[74],stage1_12[122],stage1_11[141],stage1_10[171]}
   );
   gpc615_5 gpc445 (
      {stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359], stage0_10[360]},
      {stage0_11[395]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[75],stage1_12[123],stage1_11[142],stage1_10[172]}
   );
   gpc615_5 gpc446 (
      {stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage0_11[396]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[76],stage1_12[124],stage1_11[143],stage1_10[173]}
   );
   gpc615_5 gpc447 (
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370]},
      {stage0_11[397]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[77],stage1_12[125],stage1_11[144],stage1_10[174]}
   );
   gpc615_5 gpc448 (
      {stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_11[398]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[78],stage1_12[126],stage1_11[145],stage1_10[175]}
   );
   gpc615_5 gpc449 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380]},
      {stage0_11[399]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[79],stage1_12[127],stage1_11[146],stage1_10[176]}
   );
   gpc2135_5 gpc450 (
      {stage0_11[400], stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404]},
      {stage0_12[96], stage0_12[97], stage0_12[98]},
      {stage0_13[0]},
      {stage0_14[0], stage0_14[1]},
      {stage1_15[0],stage1_14[16],stage1_13[80],stage1_12[128],stage1_11[147]}
   );
   gpc606_5 gpc451 (
      {stage0_11[405], stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5], stage0_13[6]},
      {stage1_15[1],stage1_14[17],stage1_13[81],stage1_12[129],stage1_11[148]}
   );
   gpc606_5 gpc452 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415], stage0_11[416]},
      {stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12]},
      {stage1_15[2],stage1_14[18],stage1_13[82],stage1_12[130],stage1_11[149]}
   );
   gpc606_5 gpc453 (
      {stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420], stage0_11[421], stage0_11[422]},
      {stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18]},
      {stage1_15[3],stage1_14[19],stage1_13[83],stage1_12[131],stage1_11[150]}
   );
   gpc606_5 gpc454 (
      {stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104]},
      {stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7]},
      {stage1_16[0],stage1_15[4],stage1_14[20],stage1_13[84],stage1_12[132]}
   );
   gpc606_5 gpc455 (
      {stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110]},
      {stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13]},
      {stage1_16[1],stage1_15[5],stage1_14[21],stage1_13[85],stage1_12[133]}
   );
   gpc606_5 gpc456 (
      {stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116]},
      {stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19]},
      {stage1_16[2],stage1_15[6],stage1_14[22],stage1_13[86],stage1_12[134]}
   );
   gpc606_5 gpc457 (
      {stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25]},
      {stage1_16[3],stage1_15[7],stage1_14[23],stage1_13[87],stage1_12[135]}
   );
   gpc606_5 gpc458 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128]},
      {stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31]},
      {stage1_16[4],stage1_15[8],stage1_14[24],stage1_13[88],stage1_12[136]}
   );
   gpc606_5 gpc459 (
      {stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134]},
      {stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36], stage0_14[37]},
      {stage1_16[5],stage1_15[9],stage1_14[25],stage1_13[89],stage1_12[137]}
   );
   gpc606_5 gpc460 (
      {stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140]},
      {stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42], stage0_14[43]},
      {stage1_16[6],stage1_15[10],stage1_14[26],stage1_13[90],stage1_12[138]}
   );
   gpc606_5 gpc461 (
      {stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146]},
      {stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49]},
      {stage1_16[7],stage1_15[11],stage1_14[27],stage1_13[91],stage1_12[139]}
   );
   gpc606_5 gpc462 (
      {stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152]},
      {stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55]},
      {stage1_16[8],stage1_15[12],stage1_14[28],stage1_13[92],stage1_12[140]}
   );
   gpc606_5 gpc463 (
      {stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158]},
      {stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60], stage0_14[61]},
      {stage1_16[9],stage1_15[13],stage1_14[29],stage1_13[93],stage1_12[141]}
   );
   gpc606_5 gpc464 (
      {stage0_12[159], stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164]},
      {stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67]},
      {stage1_16[10],stage1_15[14],stage1_14[30],stage1_13[94],stage1_12[142]}
   );
   gpc606_5 gpc465 (
      {stage0_12[165], stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169], stage0_12[170]},
      {stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73]},
      {stage1_16[11],stage1_15[15],stage1_14[31],stage1_13[95],stage1_12[143]}
   );
   gpc606_5 gpc466 (
      {stage0_12[171], stage0_12[172], stage0_12[173], stage0_12[174], stage0_12[175], stage0_12[176]},
      {stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79]},
      {stage1_16[12],stage1_15[16],stage1_14[32],stage1_13[96],stage1_12[144]}
   );
   gpc606_5 gpc467 (
      {stage0_12[177], stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182]},
      {stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83], stage0_14[84], stage0_14[85]},
      {stage1_16[13],stage1_15[17],stage1_14[33],stage1_13[97],stage1_12[145]}
   );
   gpc606_5 gpc468 (
      {stage0_12[183], stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188]},
      {stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89], stage0_14[90], stage0_14[91]},
      {stage1_16[14],stage1_15[18],stage1_14[34],stage1_13[98],stage1_12[146]}
   );
   gpc606_5 gpc469 (
      {stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194]},
      {stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95], stage0_14[96], stage0_14[97]},
      {stage1_16[15],stage1_15[19],stage1_14[35],stage1_13[99],stage1_12[147]}
   );
   gpc606_5 gpc470 (
      {stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199], stage0_12[200]},
      {stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102], stage0_14[103]},
      {stage1_16[16],stage1_15[20],stage1_14[36],stage1_13[100],stage1_12[148]}
   );
   gpc606_5 gpc471 (
      {stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205], stage0_12[206]},
      {stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108], stage0_14[109]},
      {stage1_16[17],stage1_15[21],stage1_14[37],stage1_13[101],stage1_12[149]}
   );
   gpc606_5 gpc472 (
      {stage0_12[207], stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212]},
      {stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113], stage0_14[114], stage0_14[115]},
      {stage1_16[18],stage1_15[22],stage1_14[38],stage1_13[102],stage1_12[150]}
   );
   gpc606_5 gpc473 (
      {stage0_12[213], stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218]},
      {stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119], stage0_14[120], stage0_14[121]},
      {stage1_16[19],stage1_15[23],stage1_14[39],stage1_13[103],stage1_12[151]}
   );
   gpc606_5 gpc474 (
      {stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223], stage0_12[224]},
      {stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126], stage0_14[127]},
      {stage1_16[20],stage1_15[24],stage1_14[40],stage1_13[104],stage1_12[152]}
   );
   gpc606_5 gpc475 (
      {stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229], stage0_12[230]},
      {stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132], stage0_14[133]},
      {stage1_16[21],stage1_15[25],stage1_14[41],stage1_13[105],stage1_12[153]}
   );
   gpc606_5 gpc476 (
      {stage0_12[231], stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236]},
      {stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage1_16[22],stage1_15[26],stage1_14[42],stage1_13[106],stage1_12[154]}
   );
   gpc606_5 gpc477 (
      {stage0_12[237], stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242]},
      {stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143], stage0_14[144], stage0_14[145]},
      {stage1_16[23],stage1_15[27],stage1_14[43],stage1_13[107],stage1_12[155]}
   );
   gpc606_5 gpc478 (
      {stage0_12[243], stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248]},
      {stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149], stage0_14[150], stage0_14[151]},
      {stage1_16[24],stage1_15[28],stage1_14[44],stage1_13[108],stage1_12[156]}
   );
   gpc606_5 gpc479 (
      {stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254]},
      {stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156], stage0_14[157]},
      {stage1_16[25],stage1_15[29],stage1_14[45],stage1_13[109],stage1_12[157]}
   );
   gpc606_5 gpc480 (
      {stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258], stage0_12[259], stage0_12[260]},
      {stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161], stage0_14[162], stage0_14[163]},
      {stage1_16[26],stage1_15[30],stage1_14[46],stage1_13[110],stage1_12[158]}
   );
   gpc606_5 gpc481 (
      {stage0_12[261], stage0_12[262], stage0_12[263], stage0_12[264], stage0_12[265], stage0_12[266]},
      {stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167], stage0_14[168], stage0_14[169]},
      {stage1_16[27],stage1_15[31],stage1_14[47],stage1_13[111],stage1_12[159]}
   );
   gpc606_5 gpc482 (
      {stage0_12[267], stage0_12[268], stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272]},
      {stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173], stage0_14[174], stage0_14[175]},
      {stage1_16[28],stage1_15[32],stage1_14[48],stage1_13[112],stage1_12[160]}
   );
   gpc606_5 gpc483 (
      {stage0_12[273], stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278]},
      {stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179], stage0_14[180], stage0_14[181]},
      {stage1_16[29],stage1_15[33],stage1_14[49],stage1_13[113],stage1_12[161]}
   );
   gpc606_5 gpc484 (
      {stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283], stage0_12[284]},
      {stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185], stage0_14[186], stage0_14[187]},
      {stage1_16[30],stage1_15[34],stage1_14[50],stage1_13[114],stage1_12[162]}
   );
   gpc606_5 gpc485 (
      {stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288], stage0_12[289], stage0_12[290]},
      {stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191], stage0_14[192], stage0_14[193]},
      {stage1_16[31],stage1_15[35],stage1_14[51],stage1_13[115],stage1_12[163]}
   );
   gpc606_5 gpc486 (
      {stage0_12[291], stage0_12[292], stage0_12[293], stage0_12[294], stage0_12[295], stage0_12[296]},
      {stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197], stage0_14[198], stage0_14[199]},
      {stage1_16[32],stage1_15[36],stage1_14[52],stage1_13[116],stage1_12[164]}
   );
   gpc606_5 gpc487 (
      {stage0_12[297], stage0_12[298], stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302]},
      {stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203], stage0_14[204], stage0_14[205]},
      {stage1_16[33],stage1_15[37],stage1_14[53],stage1_13[117],stage1_12[165]}
   );
   gpc606_5 gpc488 (
      {stage0_12[303], stage0_12[304], stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308]},
      {stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209], stage0_14[210], stage0_14[211]},
      {stage1_16[34],stage1_15[38],stage1_14[54],stage1_13[118],stage1_12[166]}
   );
   gpc606_5 gpc489 (
      {stage0_12[309], stage0_12[310], stage0_12[311], stage0_12[312], stage0_12[313], stage0_12[314]},
      {stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215], stage0_14[216], stage0_14[217]},
      {stage1_16[35],stage1_15[39],stage1_14[55],stage1_13[119],stage1_12[167]}
   );
   gpc606_5 gpc490 (
      {stage0_12[315], stage0_12[316], stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320]},
      {stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221], stage0_14[222], stage0_14[223]},
      {stage1_16[36],stage1_15[40],stage1_14[56],stage1_13[120],stage1_12[168]}
   );
   gpc615_5 gpc491 (
      {stage0_12[321], stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325]},
      {stage0_13[19]},
      {stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227], stage0_14[228], stage0_14[229]},
      {stage1_16[37],stage1_15[41],stage1_14[57],stage1_13[121],stage1_12[169]}
   );
   gpc615_5 gpc492 (
      {stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330]},
      {stage0_13[20]},
      {stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233], stage0_14[234], stage0_14[235]},
      {stage1_16[38],stage1_15[42],stage1_14[58],stage1_13[122],stage1_12[170]}
   );
   gpc615_5 gpc493 (
      {stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_13[21]},
      {stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239], stage0_14[240], stage0_14[241]},
      {stage1_16[39],stage1_15[43],stage1_14[59],stage1_13[123],stage1_12[171]}
   );
   gpc615_5 gpc494 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340]},
      {stage0_13[22]},
      {stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245], stage0_14[246], stage0_14[247]},
      {stage1_16[40],stage1_15[44],stage1_14[60],stage1_13[124],stage1_12[172]}
   );
   gpc615_5 gpc495 (
      {stage0_12[341], stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345]},
      {stage0_13[23]},
      {stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251], stage0_14[252], stage0_14[253]},
      {stage1_16[41],stage1_15[45],stage1_14[61],stage1_13[125],stage1_12[173]}
   );
   gpc615_5 gpc496 (
      {stage0_12[346], stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350]},
      {stage0_13[24]},
      {stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257], stage0_14[258], stage0_14[259]},
      {stage1_16[42],stage1_15[46],stage1_14[62],stage1_13[126],stage1_12[174]}
   );
   gpc615_5 gpc497 (
      {stage0_12[351], stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355]},
      {stage0_13[25]},
      {stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263], stage0_14[264], stage0_14[265]},
      {stage1_16[43],stage1_15[47],stage1_14[63],stage1_13[127],stage1_12[175]}
   );
   gpc615_5 gpc498 (
      {stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360]},
      {stage0_13[26]},
      {stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269], stage0_14[270], stage0_14[271]},
      {stage1_16[44],stage1_15[48],stage1_14[64],stage1_13[128],stage1_12[176]}
   );
   gpc615_5 gpc499 (
      {stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_13[27]},
      {stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275], stage0_14[276], stage0_14[277]},
      {stage1_16[45],stage1_15[49],stage1_14[65],stage1_13[129],stage1_12[177]}
   );
   gpc615_5 gpc500 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370]},
      {stage0_13[28]},
      {stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281], stage0_14[282], stage0_14[283]},
      {stage1_16[46],stage1_15[50],stage1_14[66],stage1_13[130],stage1_12[178]}
   );
   gpc615_5 gpc501 (
      {stage0_12[371], stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375]},
      {stage0_13[29]},
      {stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287], stage0_14[288], stage0_14[289]},
      {stage1_16[47],stage1_15[51],stage1_14[67],stage1_13[131],stage1_12[179]}
   );
   gpc615_5 gpc502 (
      {stage0_12[376], stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380]},
      {stage0_13[30]},
      {stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293], stage0_14[294], stage0_14[295]},
      {stage1_16[48],stage1_15[52],stage1_14[68],stage1_13[132],stage1_12[180]}
   );
   gpc615_5 gpc503 (
      {stage0_12[381], stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385]},
      {stage0_13[31]},
      {stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299], stage0_14[300], stage0_14[301]},
      {stage1_16[49],stage1_15[53],stage1_14[69],stage1_13[133],stage1_12[181]}
   );
   gpc615_5 gpc504 (
      {stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390]},
      {stage0_13[32]},
      {stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305], stage0_14[306], stage0_14[307]},
      {stage1_16[50],stage1_15[54],stage1_14[70],stage1_13[134],stage1_12[182]}
   );
   gpc615_5 gpc505 (
      {stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_13[33]},
      {stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311], stage0_14[312], stage0_14[313]},
      {stage1_16[51],stage1_15[55],stage1_14[71],stage1_13[135],stage1_12[183]}
   );
   gpc615_5 gpc506 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400]},
      {stage0_13[34]},
      {stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317], stage0_14[318], stage0_14[319]},
      {stage1_16[52],stage1_15[56],stage1_14[72],stage1_13[136],stage1_12[184]}
   );
   gpc615_5 gpc507 (
      {stage0_12[401], stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405]},
      {stage0_13[35]},
      {stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323], stage0_14[324], stage0_14[325]},
      {stage1_16[53],stage1_15[57],stage1_14[73],stage1_13[137],stage1_12[185]}
   );
   gpc615_5 gpc508 (
      {stage0_12[406], stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410]},
      {stage0_13[36]},
      {stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329], stage0_14[330], stage0_14[331]},
      {stage1_16[54],stage1_15[58],stage1_14[74],stage1_13[138],stage1_12[186]}
   );
   gpc615_5 gpc509 (
      {stage0_12[411], stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415]},
      {stage0_13[37]},
      {stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335], stage0_14[336], stage0_14[337]},
      {stage1_16[55],stage1_15[59],stage1_14[75],stage1_13[139],stage1_12[187]}
   );
   gpc615_5 gpc510 (
      {stage0_12[416], stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420]},
      {stage0_13[38]},
      {stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341], stage0_14[342], stage0_14[343]},
      {stage1_16[56],stage1_15[60],stage1_14[76],stage1_13[140],stage1_12[188]}
   );
   gpc615_5 gpc511 (
      {stage0_12[421], stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425]},
      {stage0_13[39]},
      {stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347], stage0_14[348], stage0_14[349]},
      {stage1_16[57],stage1_15[61],stage1_14[77],stage1_13[141],stage1_12[189]}
   );
   gpc615_5 gpc512 (
      {stage0_12[426], stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430]},
      {stage0_13[40]},
      {stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353], stage0_14[354], stage0_14[355]},
      {stage1_16[58],stage1_15[62],stage1_14[78],stage1_13[142],stage1_12[190]}
   );
   gpc615_5 gpc513 (
      {stage0_12[431], stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435]},
      {stage0_13[41]},
      {stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359], stage0_14[360], stage0_14[361]},
      {stage1_16[59],stage1_15[63],stage1_14[79],stage1_13[143],stage1_12[191]}
   );
   gpc615_5 gpc514 (
      {stage0_12[436], stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440]},
      {stage0_13[42]},
      {stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365], stage0_14[366], stage0_14[367]},
      {stage1_16[60],stage1_15[64],stage1_14[80],stage1_13[144],stage1_12[192]}
   );
   gpc615_5 gpc515 (
      {stage0_12[441], stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445]},
      {stage0_13[43]},
      {stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371], stage0_14[372], stage0_14[373]},
      {stage1_16[61],stage1_15[65],stage1_14[81],stage1_13[145],stage1_12[193]}
   );
   gpc615_5 gpc516 (
      {stage0_12[446], stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450]},
      {stage0_13[44]},
      {stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377], stage0_14[378], stage0_14[379]},
      {stage1_16[62],stage1_15[66],stage1_14[82],stage1_13[146],stage1_12[194]}
   );
   gpc615_5 gpc517 (
      {stage0_12[451], stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455]},
      {stage0_13[45]},
      {stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383], stage0_14[384], stage0_14[385]},
      {stage1_16[63],stage1_15[67],stage1_14[83],stage1_13[147],stage1_12[195]}
   );
   gpc615_5 gpc518 (
      {stage0_12[456], stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460]},
      {stage0_13[46]},
      {stage0_14[386], stage0_14[387], stage0_14[388], stage0_14[389], stage0_14[390], stage0_14[391]},
      {stage1_16[64],stage1_15[68],stage1_14[84],stage1_13[148],stage1_12[196]}
   );
   gpc615_5 gpc519 (
      {stage0_12[461], stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465]},
      {stage0_13[47]},
      {stage0_14[392], stage0_14[393], stage0_14[394], stage0_14[395], stage0_14[396], stage0_14[397]},
      {stage1_16[65],stage1_15[69],stage1_14[85],stage1_13[149],stage1_12[197]}
   );
   gpc615_5 gpc520 (
      {stage0_12[466], stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470]},
      {stage0_13[48]},
      {stage0_14[398], stage0_14[399], stage0_14[400], stage0_14[401], stage0_14[402], stage0_14[403]},
      {stage1_16[66],stage1_15[70],stage1_14[86],stage1_13[150],stage1_12[198]}
   );
   gpc615_5 gpc521 (
      {stage0_12[471], stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475]},
      {stage0_13[49]},
      {stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407], stage0_14[408], stage0_14[409]},
      {stage1_16[67],stage1_15[71],stage1_14[87],stage1_13[151],stage1_12[199]}
   );
   gpc615_5 gpc522 (
      {stage0_12[476], stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480]},
      {stage0_13[50]},
      {stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413], stage0_14[414], stage0_14[415]},
      {stage1_16[68],stage1_15[72],stage1_14[88],stage1_13[152],stage1_12[200]}
   );
   gpc615_5 gpc523 (
      {stage0_12[481], stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485]},
      {stage0_13[51]},
      {stage0_14[416], stage0_14[417], stage0_14[418], stage0_14[419], stage0_14[420], stage0_14[421]},
      {stage1_16[69],stage1_15[73],stage1_14[89],stage1_13[153],stage1_12[201]}
   );
   gpc606_5 gpc524 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[70],stage1_15[74],stage1_14[90],stage1_13[154]}
   );
   gpc606_5 gpc525 (
      {stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[71],stage1_15[75],stage1_14[91],stage1_13[155]}
   );
   gpc606_5 gpc526 (
      {stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[72],stage1_15[76],stage1_14[92],stage1_13[156]}
   );
   gpc606_5 gpc527 (
      {stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[73],stage1_15[77],stage1_14[93],stage1_13[157]}
   );
   gpc606_5 gpc528 (
      {stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[74],stage1_15[78],stage1_14[94],stage1_13[158]}
   );
   gpc606_5 gpc529 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[75],stage1_15[79],stage1_14[95],stage1_13[159]}
   );
   gpc606_5 gpc530 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[76],stage1_15[80],stage1_14[96],stage1_13[160]}
   );
   gpc606_5 gpc531 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[77],stage1_15[81],stage1_14[97],stage1_13[161]}
   );
   gpc606_5 gpc532 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[78],stage1_15[82],stage1_14[98],stage1_13[162]}
   );
   gpc606_5 gpc533 (
      {stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[79],stage1_15[83],stage1_14[99],stage1_13[163]}
   );
   gpc606_5 gpc534 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[80],stage1_15[84],stage1_14[100],stage1_13[164]}
   );
   gpc606_5 gpc535 (
      {stage0_13[118], stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[81],stage1_15[85],stage1_14[101],stage1_13[165]}
   );
   gpc606_5 gpc536 (
      {stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[82],stage1_15[86],stage1_14[102],stage1_13[166]}
   );
   gpc606_5 gpc537 (
      {stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[83],stage1_15[87],stage1_14[103],stage1_13[167]}
   );
   gpc606_5 gpc538 (
      {stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[84],stage1_15[88],stage1_14[104],stage1_13[168]}
   );
   gpc606_5 gpc539 (
      {stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[85],stage1_15[89],stage1_14[105],stage1_13[169]}
   );
   gpc606_5 gpc540 (
      {stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[86],stage1_15[90],stage1_14[106],stage1_13[170]}
   );
   gpc606_5 gpc541 (
      {stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[87],stage1_15[91],stage1_14[107],stage1_13[171]}
   );
   gpc606_5 gpc542 (
      {stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[88],stage1_15[92],stage1_14[108],stage1_13[172]}
   );
   gpc606_5 gpc543 (
      {stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[89],stage1_15[93],stage1_14[109],stage1_13[173]}
   );
   gpc606_5 gpc544 (
      {stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[90],stage1_15[94],stage1_14[110],stage1_13[174]}
   );
   gpc606_5 gpc545 (
      {stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[91],stage1_15[95],stage1_14[111],stage1_13[175]}
   );
   gpc606_5 gpc546 (
      {stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[92],stage1_15[96],stage1_14[112],stage1_13[176]}
   );
   gpc606_5 gpc547 (
      {stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[93],stage1_15[97],stage1_14[113],stage1_13[177]}
   );
   gpc606_5 gpc548 (
      {stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[94],stage1_15[98],stage1_14[114],stage1_13[178]}
   );
   gpc606_5 gpc549 (
      {stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[95],stage1_15[99],stage1_14[115],stage1_13[179]}
   );
   gpc606_5 gpc550 (
      {stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[96],stage1_15[100],stage1_14[116],stage1_13[180]}
   );
   gpc606_5 gpc551 (
      {stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[97],stage1_15[101],stage1_14[117],stage1_13[181]}
   );
   gpc606_5 gpc552 (
      {stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[98],stage1_15[102],stage1_14[118],stage1_13[182]}
   );
   gpc615_5 gpc553 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[422]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[99],stage1_15[103],stage1_14[119],stage1_13[183]}
   );
   gpc615_5 gpc554 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[423]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[100],stage1_15[104],stage1_14[120],stage1_13[184]}
   );
   gpc615_5 gpc555 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[424]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[101],stage1_15[105],stage1_14[121],stage1_13[185]}
   );
   gpc615_5 gpc556 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[425]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[102],stage1_15[106],stage1_14[122],stage1_13[186]}
   );
   gpc615_5 gpc557 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[426]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[103],stage1_15[107],stage1_14[123],stage1_13[187]}
   );
   gpc615_5 gpc558 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[427]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[104],stage1_15[108],stage1_14[124],stage1_13[188]}
   );
   gpc615_5 gpc559 (
      {stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_14[428]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[105],stage1_15[109],stage1_14[125],stage1_13[189]}
   );
   gpc615_5 gpc560 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265]},
      {stage0_14[429]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[106],stage1_15[110],stage1_14[126],stage1_13[190]}
   );
   gpc615_5 gpc561 (
      {stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270]},
      {stage0_14[430]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[107],stage1_15[111],stage1_14[127],stage1_13[191]}
   );
   gpc615_5 gpc562 (
      {stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_14[431]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[108],stage1_15[112],stage1_14[128],stage1_13[192]}
   );
   gpc615_5 gpc563 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280]},
      {stage0_14[432]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[109],stage1_15[113],stage1_14[129],stage1_13[193]}
   );
   gpc615_5 gpc564 (
      {stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285]},
      {stage0_14[433]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[110],stage1_15[114],stage1_14[130],stage1_13[194]}
   );
   gpc615_5 gpc565 (
      {stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_14[434]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[111],stage1_15[115],stage1_14[131],stage1_13[195]}
   );
   gpc615_5 gpc566 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295]},
      {stage0_14[435]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[112],stage1_15[116],stage1_14[132],stage1_13[196]}
   );
   gpc615_5 gpc567 (
      {stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300]},
      {stage0_14[436]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[113],stage1_15[117],stage1_14[133],stage1_13[197]}
   );
   gpc615_5 gpc568 (
      {stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_14[437]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[114],stage1_15[118],stage1_14[134],stage1_13[198]}
   );
   gpc615_5 gpc569 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310]},
      {stage0_14[438]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[115],stage1_15[119],stage1_14[135],stage1_13[199]}
   );
   gpc615_5 gpc570 (
      {stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315]},
      {stage0_14[439]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[116],stage1_15[120],stage1_14[136],stage1_13[200]}
   );
   gpc615_5 gpc571 (
      {stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_14[440]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[117],stage1_15[121],stage1_14[137],stage1_13[201]}
   );
   gpc615_5 gpc572 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325]},
      {stage0_14[441]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[118],stage1_15[122],stage1_14[138],stage1_13[202]}
   );
   gpc615_5 gpc573 (
      {stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330]},
      {stage0_14[442]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[119],stage1_15[123],stage1_14[139],stage1_13[203]}
   );
   gpc615_5 gpc574 (
      {stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_14[443]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[120],stage1_15[124],stage1_14[140],stage1_13[204]}
   );
   gpc615_5 gpc575 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340]},
      {stage0_14[444]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[121],stage1_15[125],stage1_14[141],stage1_13[205]}
   );
   gpc615_5 gpc576 (
      {stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345]},
      {stage0_14[445]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[122],stage1_15[126],stage1_14[142],stage1_13[206]}
   );
   gpc615_5 gpc577 (
      {stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_14[446]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[123],stage1_15[127],stage1_14[143],stage1_13[207]}
   );
   gpc615_5 gpc578 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355]},
      {stage0_14[447]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[124],stage1_15[128],stage1_14[144],stage1_13[208]}
   );
   gpc615_5 gpc579 (
      {stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360]},
      {stage0_14[448]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[125],stage1_15[129],stage1_14[145],stage1_13[209]}
   );
   gpc615_5 gpc580 (
      {stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_14[449]},
      {stage0_15[336], stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage1_17[56],stage1_16[126],stage1_15[130],stage1_14[146],stage1_13[210]}
   );
   gpc615_5 gpc581 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370]},
      {stage0_14[450]},
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347]},
      {stage1_17[57],stage1_16[127],stage1_15[131],stage1_14[147],stage1_13[211]}
   );
   gpc615_5 gpc582 (
      {stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375]},
      {stage0_14[451]},
      {stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage1_17[58],stage1_16[128],stage1_15[132],stage1_14[148],stage1_13[212]}
   );
   gpc615_5 gpc583 (
      {stage0_13[376], stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380]},
      {stage0_14[452]},
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage1_17[59],stage1_16[129],stage1_15[133],stage1_14[149],stage1_13[213]}
   );
   gpc615_5 gpc584 (
      {stage0_13[381], stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385]},
      {stage0_14[453]},
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage1_17[60],stage1_16[130],stage1_15[134],stage1_14[150],stage1_13[214]}
   );
   gpc615_5 gpc585 (
      {stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390]},
      {stage0_14[454]},
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage1_17[61],stage1_16[131],stage1_15[135],stage1_14[151],stage1_13[215]}
   );
   gpc615_5 gpc586 (
      {stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_14[455]},
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377]},
      {stage1_17[62],stage1_16[132],stage1_15[136],stage1_14[152],stage1_13[216]}
   );
   gpc615_5 gpc587 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400]},
      {stage0_14[456]},
      {stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage1_17[63],stage1_16[133],stage1_15[137],stage1_14[153],stage1_13[217]}
   );
   gpc615_5 gpc588 (
      {stage0_13[401], stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405]},
      {stage0_14[457]},
      {stage0_15[384], stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389]},
      {stage1_17[64],stage1_16[134],stage1_15[138],stage1_14[154],stage1_13[218]}
   );
   gpc615_5 gpc589 (
      {stage0_13[406], stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410]},
      {stage0_14[458]},
      {stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395]},
      {stage1_17[65],stage1_16[135],stage1_15[139],stage1_14[155],stage1_13[219]}
   );
   gpc615_5 gpc590 (
      {stage0_13[411], stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415]},
      {stage0_14[459]},
      {stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400], stage0_15[401]},
      {stage1_17[66],stage1_16[136],stage1_15[140],stage1_14[156],stage1_13[220]}
   );
   gpc615_5 gpc591 (
      {stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420]},
      {stage0_14[460]},
      {stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405], stage0_15[406], stage0_15[407]},
      {stage1_17[67],stage1_16[137],stage1_15[141],stage1_14[157],stage1_13[221]}
   );
   gpc615_5 gpc592 (
      {stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_14[461]},
      {stage0_15[408], stage0_15[409], stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413]},
      {stage1_17[68],stage1_16[138],stage1_15[142],stage1_14[158],stage1_13[222]}
   );
   gpc615_5 gpc593 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430]},
      {stage0_14[462]},
      {stage0_15[414], stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419]},
      {stage1_17[69],stage1_16[139],stage1_15[143],stage1_14[159],stage1_13[223]}
   );
   gpc615_5 gpc594 (
      {stage0_13[431], stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435]},
      {stage0_14[463]},
      {stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425]},
      {stage1_17[70],stage1_16[140],stage1_15[144],stage1_14[160],stage1_13[224]}
   );
   gpc615_5 gpc595 (
      {stage0_13[436], stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440]},
      {stage0_14[464]},
      {stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430], stage0_15[431]},
      {stage1_17[71],stage1_16[141],stage1_15[145],stage1_14[161],stage1_13[225]}
   );
   gpc615_5 gpc596 (
      {stage0_13[441], stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445]},
      {stage0_14[465]},
      {stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435], stage0_15[436], stage0_15[437]},
      {stage1_17[72],stage1_16[142],stage1_15[146],stage1_14[162],stage1_13[226]}
   );
   gpc615_5 gpc597 (
      {stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450]},
      {stage0_14[466]},
      {stage0_15[438], stage0_15[439], stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443]},
      {stage1_17[73],stage1_16[143],stage1_15[147],stage1_14[163],stage1_13[227]}
   );
   gpc615_5 gpc598 (
      {stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_14[467]},
      {stage0_15[444], stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449]},
      {stage1_17[74],stage1_16[144],stage1_15[148],stage1_14[164],stage1_13[228]}
   );
   gpc615_5 gpc599 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460]},
      {stage0_14[468]},
      {stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455]},
      {stage1_17[75],stage1_16[145],stage1_15[149],stage1_14[165],stage1_13[229]}
   );
   gpc615_5 gpc600 (
      {stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465]},
      {stage0_14[469]},
      {stage0_15[456], stage0_15[457], stage0_15[458], stage0_15[459], stage0_15[460], stage0_15[461]},
      {stage1_17[76],stage1_16[146],stage1_15[150],stage1_14[166],stage1_13[230]}
   );
   gpc615_5 gpc601 (
      {stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_14[470]},
      {stage0_15[462], stage0_15[463], stage0_15[464], stage0_15[465], stage0_15[466], stage0_15[467]},
      {stage1_17[77],stage1_16[147],stage1_15[151],stage1_14[167],stage1_13[231]}
   );
   gpc615_5 gpc602 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475]},
      {stage0_14[471]},
      {stage0_15[468], stage0_15[469], stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473]},
      {stage1_17[78],stage1_16[148],stage1_15[152],stage1_14[168],stage1_13[232]}
   );
   gpc615_5 gpc603 (
      {stage0_13[476], stage0_13[477], stage0_13[478], stage0_13[479], stage0_13[480]},
      {stage0_14[472]},
      {stage0_15[474], stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478], stage0_15[479]},
      {stage1_17[79],stage1_16[149],stage1_15[153],stage1_14[169],stage1_13[233]}
   );
   gpc615_5 gpc604 (
      {stage0_13[481], stage0_13[482], stage0_13[483], stage0_13[484], stage0_13[485]},
      {stage0_14[473]},
      {stage0_15[480], stage0_15[481], stage0_15[482], stage0_15[483], stage0_15[484], stage0_15[485]},
      {stage1_17[80],stage1_16[150],stage1_15[154],stage1_14[170],stage1_13[234]}
   );
   gpc1_1 gpc605 (
      {stage0_0[423]},
      {stage1_0[85]}
   );
   gpc1_1 gpc606 (
      {stage0_0[424]},
      {stage1_0[86]}
   );
   gpc1_1 gpc607 (
      {stage0_0[425]},
      {stage1_0[87]}
   );
   gpc1_1 gpc608 (
      {stage0_0[426]},
      {stage1_0[88]}
   );
   gpc1_1 gpc609 (
      {stage0_0[427]},
      {stage1_0[89]}
   );
   gpc1_1 gpc610 (
      {stage0_0[428]},
      {stage1_0[90]}
   );
   gpc1_1 gpc611 (
      {stage0_0[429]},
      {stage1_0[91]}
   );
   gpc1_1 gpc612 (
      {stage0_0[430]},
      {stage1_0[92]}
   );
   gpc1_1 gpc613 (
      {stage0_0[431]},
      {stage1_0[93]}
   );
   gpc1_1 gpc614 (
      {stage0_0[432]},
      {stage1_0[94]}
   );
   gpc1_1 gpc615 (
      {stage0_0[433]},
      {stage1_0[95]}
   );
   gpc1_1 gpc616 (
      {stage0_0[434]},
      {stage1_0[96]}
   );
   gpc1_1 gpc617 (
      {stage0_0[435]},
      {stage1_0[97]}
   );
   gpc1_1 gpc618 (
      {stage0_0[436]},
      {stage1_0[98]}
   );
   gpc1_1 gpc619 (
      {stage0_0[437]},
      {stage1_0[99]}
   );
   gpc1_1 gpc620 (
      {stage0_0[438]},
      {stage1_0[100]}
   );
   gpc1_1 gpc621 (
      {stage0_0[439]},
      {stage1_0[101]}
   );
   gpc1_1 gpc622 (
      {stage0_0[440]},
      {stage1_0[102]}
   );
   gpc1_1 gpc623 (
      {stage0_0[441]},
      {stage1_0[103]}
   );
   gpc1_1 gpc624 (
      {stage0_0[442]},
      {stage1_0[104]}
   );
   gpc1_1 gpc625 (
      {stage0_0[443]},
      {stage1_0[105]}
   );
   gpc1_1 gpc626 (
      {stage0_0[444]},
      {stage1_0[106]}
   );
   gpc1_1 gpc627 (
      {stage0_0[445]},
      {stage1_0[107]}
   );
   gpc1_1 gpc628 (
      {stage0_0[446]},
      {stage1_0[108]}
   );
   gpc1_1 gpc629 (
      {stage0_0[447]},
      {stage1_0[109]}
   );
   gpc1_1 gpc630 (
      {stage0_0[448]},
      {stage1_0[110]}
   );
   gpc1_1 gpc631 (
      {stage0_0[449]},
      {stage1_0[111]}
   );
   gpc1_1 gpc632 (
      {stage0_0[450]},
      {stage1_0[112]}
   );
   gpc1_1 gpc633 (
      {stage0_0[451]},
      {stage1_0[113]}
   );
   gpc1_1 gpc634 (
      {stage0_0[452]},
      {stage1_0[114]}
   );
   gpc1_1 gpc635 (
      {stage0_0[453]},
      {stage1_0[115]}
   );
   gpc1_1 gpc636 (
      {stage0_0[454]},
      {stage1_0[116]}
   );
   gpc1_1 gpc637 (
      {stage0_0[455]},
      {stage1_0[117]}
   );
   gpc1_1 gpc638 (
      {stage0_0[456]},
      {stage1_0[118]}
   );
   gpc1_1 gpc639 (
      {stage0_0[457]},
      {stage1_0[119]}
   );
   gpc1_1 gpc640 (
      {stage0_0[458]},
      {stage1_0[120]}
   );
   gpc1_1 gpc641 (
      {stage0_0[459]},
      {stage1_0[121]}
   );
   gpc1_1 gpc642 (
      {stage0_0[460]},
      {stage1_0[122]}
   );
   gpc1_1 gpc643 (
      {stage0_0[461]},
      {stage1_0[123]}
   );
   gpc1_1 gpc644 (
      {stage0_0[462]},
      {stage1_0[124]}
   );
   gpc1_1 gpc645 (
      {stage0_0[463]},
      {stage1_0[125]}
   );
   gpc1_1 gpc646 (
      {stage0_0[464]},
      {stage1_0[126]}
   );
   gpc1_1 gpc647 (
      {stage0_0[465]},
      {stage1_0[127]}
   );
   gpc1_1 gpc648 (
      {stage0_0[466]},
      {stage1_0[128]}
   );
   gpc1_1 gpc649 (
      {stage0_0[467]},
      {stage1_0[129]}
   );
   gpc1_1 gpc650 (
      {stage0_0[468]},
      {stage1_0[130]}
   );
   gpc1_1 gpc651 (
      {stage0_0[469]},
      {stage1_0[131]}
   );
   gpc1_1 gpc652 (
      {stage0_0[470]},
      {stage1_0[132]}
   );
   gpc1_1 gpc653 (
      {stage0_0[471]},
      {stage1_0[133]}
   );
   gpc1_1 gpc654 (
      {stage0_0[472]},
      {stage1_0[134]}
   );
   gpc1_1 gpc655 (
      {stage0_0[473]},
      {stage1_0[135]}
   );
   gpc1_1 gpc656 (
      {stage0_0[474]},
      {stage1_0[136]}
   );
   gpc1_1 gpc657 (
      {stage0_0[475]},
      {stage1_0[137]}
   );
   gpc1_1 gpc658 (
      {stage0_0[476]},
      {stage1_0[138]}
   );
   gpc1_1 gpc659 (
      {stage0_0[477]},
      {stage1_0[139]}
   );
   gpc1_1 gpc660 (
      {stage0_0[478]},
      {stage1_0[140]}
   );
   gpc1_1 gpc661 (
      {stage0_0[479]},
      {stage1_0[141]}
   );
   gpc1_1 gpc662 (
      {stage0_0[480]},
      {stage1_0[142]}
   );
   gpc1_1 gpc663 (
      {stage0_0[481]},
      {stage1_0[143]}
   );
   gpc1_1 gpc664 (
      {stage0_0[482]},
      {stage1_0[144]}
   );
   gpc1_1 gpc665 (
      {stage0_0[483]},
      {stage1_0[145]}
   );
   gpc1_1 gpc666 (
      {stage0_0[484]},
      {stage1_0[146]}
   );
   gpc1_1 gpc667 (
      {stage0_0[485]},
      {stage1_0[147]}
   );
   gpc1_1 gpc668 (
      {stage0_2[484]},
      {stage1_2[166]}
   );
   gpc1_1 gpc669 (
      {stage0_2[485]},
      {stage1_2[167]}
   );
   gpc1_1 gpc670 (
      {stage0_3[416]},
      {stage1_3[174]}
   );
   gpc1_1 gpc671 (
      {stage0_3[417]},
      {stage1_3[175]}
   );
   gpc1_1 gpc672 (
      {stage0_3[418]},
      {stage1_3[176]}
   );
   gpc1_1 gpc673 (
      {stage0_3[419]},
      {stage1_3[177]}
   );
   gpc1_1 gpc674 (
      {stage0_3[420]},
      {stage1_3[178]}
   );
   gpc1_1 gpc675 (
      {stage0_3[421]},
      {stage1_3[179]}
   );
   gpc1_1 gpc676 (
      {stage0_3[422]},
      {stage1_3[180]}
   );
   gpc1_1 gpc677 (
      {stage0_3[423]},
      {stage1_3[181]}
   );
   gpc1_1 gpc678 (
      {stage0_3[424]},
      {stage1_3[182]}
   );
   gpc1_1 gpc679 (
      {stage0_3[425]},
      {stage1_3[183]}
   );
   gpc1_1 gpc680 (
      {stage0_3[426]},
      {stage1_3[184]}
   );
   gpc1_1 gpc681 (
      {stage0_3[427]},
      {stage1_3[185]}
   );
   gpc1_1 gpc682 (
      {stage0_3[428]},
      {stage1_3[186]}
   );
   gpc1_1 gpc683 (
      {stage0_3[429]},
      {stage1_3[187]}
   );
   gpc1_1 gpc684 (
      {stage0_3[430]},
      {stage1_3[188]}
   );
   gpc1_1 gpc685 (
      {stage0_3[431]},
      {stage1_3[189]}
   );
   gpc1_1 gpc686 (
      {stage0_3[432]},
      {stage1_3[190]}
   );
   gpc1_1 gpc687 (
      {stage0_3[433]},
      {stage1_3[191]}
   );
   gpc1_1 gpc688 (
      {stage0_3[434]},
      {stage1_3[192]}
   );
   gpc1_1 gpc689 (
      {stage0_3[435]},
      {stage1_3[193]}
   );
   gpc1_1 gpc690 (
      {stage0_3[436]},
      {stage1_3[194]}
   );
   gpc1_1 gpc691 (
      {stage0_3[437]},
      {stage1_3[195]}
   );
   gpc1_1 gpc692 (
      {stage0_3[438]},
      {stage1_3[196]}
   );
   gpc1_1 gpc693 (
      {stage0_3[439]},
      {stage1_3[197]}
   );
   gpc1_1 gpc694 (
      {stage0_3[440]},
      {stage1_3[198]}
   );
   gpc1_1 gpc695 (
      {stage0_3[441]},
      {stage1_3[199]}
   );
   gpc1_1 gpc696 (
      {stage0_3[442]},
      {stage1_3[200]}
   );
   gpc1_1 gpc697 (
      {stage0_3[443]},
      {stage1_3[201]}
   );
   gpc1_1 gpc698 (
      {stage0_3[444]},
      {stage1_3[202]}
   );
   gpc1_1 gpc699 (
      {stage0_3[445]},
      {stage1_3[203]}
   );
   gpc1_1 gpc700 (
      {stage0_3[446]},
      {stage1_3[204]}
   );
   gpc1_1 gpc701 (
      {stage0_3[447]},
      {stage1_3[205]}
   );
   gpc1_1 gpc702 (
      {stage0_3[448]},
      {stage1_3[206]}
   );
   gpc1_1 gpc703 (
      {stage0_3[449]},
      {stage1_3[207]}
   );
   gpc1_1 gpc704 (
      {stage0_3[450]},
      {stage1_3[208]}
   );
   gpc1_1 gpc705 (
      {stage0_3[451]},
      {stage1_3[209]}
   );
   gpc1_1 gpc706 (
      {stage0_3[452]},
      {stage1_3[210]}
   );
   gpc1_1 gpc707 (
      {stage0_3[453]},
      {stage1_3[211]}
   );
   gpc1_1 gpc708 (
      {stage0_3[454]},
      {stage1_3[212]}
   );
   gpc1_1 gpc709 (
      {stage0_3[455]},
      {stage1_3[213]}
   );
   gpc1_1 gpc710 (
      {stage0_3[456]},
      {stage1_3[214]}
   );
   gpc1_1 gpc711 (
      {stage0_3[457]},
      {stage1_3[215]}
   );
   gpc1_1 gpc712 (
      {stage0_3[458]},
      {stage1_3[216]}
   );
   gpc1_1 gpc713 (
      {stage0_3[459]},
      {stage1_3[217]}
   );
   gpc1_1 gpc714 (
      {stage0_3[460]},
      {stage1_3[218]}
   );
   gpc1_1 gpc715 (
      {stage0_3[461]},
      {stage1_3[219]}
   );
   gpc1_1 gpc716 (
      {stage0_3[462]},
      {stage1_3[220]}
   );
   gpc1_1 gpc717 (
      {stage0_3[463]},
      {stage1_3[221]}
   );
   gpc1_1 gpc718 (
      {stage0_3[464]},
      {stage1_3[222]}
   );
   gpc1_1 gpc719 (
      {stage0_3[465]},
      {stage1_3[223]}
   );
   gpc1_1 gpc720 (
      {stage0_3[466]},
      {stage1_3[224]}
   );
   gpc1_1 gpc721 (
      {stage0_3[467]},
      {stage1_3[225]}
   );
   gpc1_1 gpc722 (
      {stage0_3[468]},
      {stage1_3[226]}
   );
   gpc1_1 gpc723 (
      {stage0_3[469]},
      {stage1_3[227]}
   );
   gpc1_1 gpc724 (
      {stage0_3[470]},
      {stage1_3[228]}
   );
   gpc1_1 gpc725 (
      {stage0_3[471]},
      {stage1_3[229]}
   );
   gpc1_1 gpc726 (
      {stage0_3[472]},
      {stage1_3[230]}
   );
   gpc1_1 gpc727 (
      {stage0_3[473]},
      {stage1_3[231]}
   );
   gpc1_1 gpc728 (
      {stage0_3[474]},
      {stage1_3[232]}
   );
   gpc1_1 gpc729 (
      {stage0_3[475]},
      {stage1_3[233]}
   );
   gpc1_1 gpc730 (
      {stage0_3[476]},
      {stage1_3[234]}
   );
   gpc1_1 gpc731 (
      {stage0_3[477]},
      {stage1_3[235]}
   );
   gpc1_1 gpc732 (
      {stage0_3[478]},
      {stage1_3[236]}
   );
   gpc1_1 gpc733 (
      {stage0_3[479]},
      {stage1_3[237]}
   );
   gpc1_1 gpc734 (
      {stage0_3[480]},
      {stage1_3[238]}
   );
   gpc1_1 gpc735 (
      {stage0_3[481]},
      {stage1_3[239]}
   );
   gpc1_1 gpc736 (
      {stage0_3[482]},
      {stage1_3[240]}
   );
   gpc1_1 gpc737 (
      {stage0_3[483]},
      {stage1_3[241]}
   );
   gpc1_1 gpc738 (
      {stage0_3[484]},
      {stage1_3[242]}
   );
   gpc1_1 gpc739 (
      {stage0_3[485]},
      {stage1_3[243]}
   );
   gpc1_1 gpc740 (
      {stage0_5[337]},
      {stage1_5[188]}
   );
   gpc1_1 gpc741 (
      {stage0_5[338]},
      {stage1_5[189]}
   );
   gpc1_1 gpc742 (
      {stage0_5[339]},
      {stage1_5[190]}
   );
   gpc1_1 gpc743 (
      {stage0_5[340]},
      {stage1_5[191]}
   );
   gpc1_1 gpc744 (
      {stage0_5[341]},
      {stage1_5[192]}
   );
   gpc1_1 gpc745 (
      {stage0_5[342]},
      {stage1_5[193]}
   );
   gpc1_1 gpc746 (
      {stage0_5[343]},
      {stage1_5[194]}
   );
   gpc1_1 gpc747 (
      {stage0_5[344]},
      {stage1_5[195]}
   );
   gpc1_1 gpc748 (
      {stage0_5[345]},
      {stage1_5[196]}
   );
   gpc1_1 gpc749 (
      {stage0_5[346]},
      {stage1_5[197]}
   );
   gpc1_1 gpc750 (
      {stage0_5[347]},
      {stage1_5[198]}
   );
   gpc1_1 gpc751 (
      {stage0_5[348]},
      {stage1_5[199]}
   );
   gpc1_1 gpc752 (
      {stage0_5[349]},
      {stage1_5[200]}
   );
   gpc1_1 gpc753 (
      {stage0_5[350]},
      {stage1_5[201]}
   );
   gpc1_1 gpc754 (
      {stage0_5[351]},
      {stage1_5[202]}
   );
   gpc1_1 gpc755 (
      {stage0_5[352]},
      {stage1_5[203]}
   );
   gpc1_1 gpc756 (
      {stage0_5[353]},
      {stage1_5[204]}
   );
   gpc1_1 gpc757 (
      {stage0_5[354]},
      {stage1_5[205]}
   );
   gpc1_1 gpc758 (
      {stage0_5[355]},
      {stage1_5[206]}
   );
   gpc1_1 gpc759 (
      {stage0_5[356]},
      {stage1_5[207]}
   );
   gpc1_1 gpc760 (
      {stage0_5[357]},
      {stage1_5[208]}
   );
   gpc1_1 gpc761 (
      {stage0_5[358]},
      {stage1_5[209]}
   );
   gpc1_1 gpc762 (
      {stage0_5[359]},
      {stage1_5[210]}
   );
   gpc1_1 gpc763 (
      {stage0_5[360]},
      {stage1_5[211]}
   );
   gpc1_1 gpc764 (
      {stage0_5[361]},
      {stage1_5[212]}
   );
   gpc1_1 gpc765 (
      {stage0_5[362]},
      {stage1_5[213]}
   );
   gpc1_1 gpc766 (
      {stage0_5[363]},
      {stage1_5[214]}
   );
   gpc1_1 gpc767 (
      {stage0_5[364]},
      {stage1_5[215]}
   );
   gpc1_1 gpc768 (
      {stage0_5[365]},
      {stage1_5[216]}
   );
   gpc1_1 gpc769 (
      {stage0_5[366]},
      {stage1_5[217]}
   );
   gpc1_1 gpc770 (
      {stage0_5[367]},
      {stage1_5[218]}
   );
   gpc1_1 gpc771 (
      {stage0_5[368]},
      {stage1_5[219]}
   );
   gpc1_1 gpc772 (
      {stage0_5[369]},
      {stage1_5[220]}
   );
   gpc1_1 gpc773 (
      {stage0_5[370]},
      {stage1_5[221]}
   );
   gpc1_1 gpc774 (
      {stage0_5[371]},
      {stage1_5[222]}
   );
   gpc1_1 gpc775 (
      {stage0_5[372]},
      {stage1_5[223]}
   );
   gpc1_1 gpc776 (
      {stage0_5[373]},
      {stage1_5[224]}
   );
   gpc1_1 gpc777 (
      {stage0_5[374]},
      {stage1_5[225]}
   );
   gpc1_1 gpc778 (
      {stage0_5[375]},
      {stage1_5[226]}
   );
   gpc1_1 gpc779 (
      {stage0_5[376]},
      {stage1_5[227]}
   );
   gpc1_1 gpc780 (
      {stage0_5[377]},
      {stage1_5[228]}
   );
   gpc1_1 gpc781 (
      {stage0_5[378]},
      {stage1_5[229]}
   );
   gpc1_1 gpc782 (
      {stage0_5[379]},
      {stage1_5[230]}
   );
   gpc1_1 gpc783 (
      {stage0_5[380]},
      {stage1_5[231]}
   );
   gpc1_1 gpc784 (
      {stage0_5[381]},
      {stage1_5[232]}
   );
   gpc1_1 gpc785 (
      {stage0_5[382]},
      {stage1_5[233]}
   );
   gpc1_1 gpc786 (
      {stage0_5[383]},
      {stage1_5[234]}
   );
   gpc1_1 gpc787 (
      {stage0_5[384]},
      {stage1_5[235]}
   );
   gpc1_1 gpc788 (
      {stage0_5[385]},
      {stage1_5[236]}
   );
   gpc1_1 gpc789 (
      {stage0_5[386]},
      {stage1_5[237]}
   );
   gpc1_1 gpc790 (
      {stage0_5[387]},
      {stage1_5[238]}
   );
   gpc1_1 gpc791 (
      {stage0_5[388]},
      {stage1_5[239]}
   );
   gpc1_1 gpc792 (
      {stage0_5[389]},
      {stage1_5[240]}
   );
   gpc1_1 gpc793 (
      {stage0_5[390]},
      {stage1_5[241]}
   );
   gpc1_1 gpc794 (
      {stage0_5[391]},
      {stage1_5[242]}
   );
   gpc1_1 gpc795 (
      {stage0_5[392]},
      {stage1_5[243]}
   );
   gpc1_1 gpc796 (
      {stage0_5[393]},
      {stage1_5[244]}
   );
   gpc1_1 gpc797 (
      {stage0_5[394]},
      {stage1_5[245]}
   );
   gpc1_1 gpc798 (
      {stage0_5[395]},
      {stage1_5[246]}
   );
   gpc1_1 gpc799 (
      {stage0_5[396]},
      {stage1_5[247]}
   );
   gpc1_1 gpc800 (
      {stage0_5[397]},
      {stage1_5[248]}
   );
   gpc1_1 gpc801 (
      {stage0_5[398]},
      {stage1_5[249]}
   );
   gpc1_1 gpc802 (
      {stage0_5[399]},
      {stage1_5[250]}
   );
   gpc1_1 gpc803 (
      {stage0_5[400]},
      {stage1_5[251]}
   );
   gpc1_1 gpc804 (
      {stage0_5[401]},
      {stage1_5[252]}
   );
   gpc1_1 gpc805 (
      {stage0_5[402]},
      {stage1_5[253]}
   );
   gpc1_1 gpc806 (
      {stage0_5[403]},
      {stage1_5[254]}
   );
   gpc1_1 gpc807 (
      {stage0_5[404]},
      {stage1_5[255]}
   );
   gpc1_1 gpc808 (
      {stage0_5[405]},
      {stage1_5[256]}
   );
   gpc1_1 gpc809 (
      {stage0_5[406]},
      {stage1_5[257]}
   );
   gpc1_1 gpc810 (
      {stage0_5[407]},
      {stage1_5[258]}
   );
   gpc1_1 gpc811 (
      {stage0_5[408]},
      {stage1_5[259]}
   );
   gpc1_1 gpc812 (
      {stage0_5[409]},
      {stage1_5[260]}
   );
   gpc1_1 gpc813 (
      {stage0_5[410]},
      {stage1_5[261]}
   );
   gpc1_1 gpc814 (
      {stage0_5[411]},
      {stage1_5[262]}
   );
   gpc1_1 gpc815 (
      {stage0_5[412]},
      {stage1_5[263]}
   );
   gpc1_1 gpc816 (
      {stage0_5[413]},
      {stage1_5[264]}
   );
   gpc1_1 gpc817 (
      {stage0_5[414]},
      {stage1_5[265]}
   );
   gpc1_1 gpc818 (
      {stage0_5[415]},
      {stage1_5[266]}
   );
   gpc1_1 gpc819 (
      {stage0_5[416]},
      {stage1_5[267]}
   );
   gpc1_1 gpc820 (
      {stage0_5[417]},
      {stage1_5[268]}
   );
   gpc1_1 gpc821 (
      {stage0_5[418]},
      {stage1_5[269]}
   );
   gpc1_1 gpc822 (
      {stage0_5[419]},
      {stage1_5[270]}
   );
   gpc1_1 gpc823 (
      {stage0_5[420]},
      {stage1_5[271]}
   );
   gpc1_1 gpc824 (
      {stage0_5[421]},
      {stage1_5[272]}
   );
   gpc1_1 gpc825 (
      {stage0_5[422]},
      {stage1_5[273]}
   );
   gpc1_1 gpc826 (
      {stage0_5[423]},
      {stage1_5[274]}
   );
   gpc1_1 gpc827 (
      {stage0_5[424]},
      {stage1_5[275]}
   );
   gpc1_1 gpc828 (
      {stage0_5[425]},
      {stage1_5[276]}
   );
   gpc1_1 gpc829 (
      {stage0_5[426]},
      {stage1_5[277]}
   );
   gpc1_1 gpc830 (
      {stage0_5[427]},
      {stage1_5[278]}
   );
   gpc1_1 gpc831 (
      {stage0_5[428]},
      {stage1_5[279]}
   );
   gpc1_1 gpc832 (
      {stage0_5[429]},
      {stage1_5[280]}
   );
   gpc1_1 gpc833 (
      {stage0_5[430]},
      {stage1_5[281]}
   );
   gpc1_1 gpc834 (
      {stage0_5[431]},
      {stage1_5[282]}
   );
   gpc1_1 gpc835 (
      {stage0_5[432]},
      {stage1_5[283]}
   );
   gpc1_1 gpc836 (
      {stage0_5[433]},
      {stage1_5[284]}
   );
   gpc1_1 gpc837 (
      {stage0_5[434]},
      {stage1_5[285]}
   );
   gpc1_1 gpc838 (
      {stage0_5[435]},
      {stage1_5[286]}
   );
   gpc1_1 gpc839 (
      {stage0_5[436]},
      {stage1_5[287]}
   );
   gpc1_1 gpc840 (
      {stage0_5[437]},
      {stage1_5[288]}
   );
   gpc1_1 gpc841 (
      {stage0_5[438]},
      {stage1_5[289]}
   );
   gpc1_1 gpc842 (
      {stage0_5[439]},
      {stage1_5[290]}
   );
   gpc1_1 gpc843 (
      {stage0_5[440]},
      {stage1_5[291]}
   );
   gpc1_1 gpc844 (
      {stage0_5[441]},
      {stage1_5[292]}
   );
   gpc1_1 gpc845 (
      {stage0_5[442]},
      {stage1_5[293]}
   );
   gpc1_1 gpc846 (
      {stage0_5[443]},
      {stage1_5[294]}
   );
   gpc1_1 gpc847 (
      {stage0_5[444]},
      {stage1_5[295]}
   );
   gpc1_1 gpc848 (
      {stage0_5[445]},
      {stage1_5[296]}
   );
   gpc1_1 gpc849 (
      {stage0_5[446]},
      {stage1_5[297]}
   );
   gpc1_1 gpc850 (
      {stage0_5[447]},
      {stage1_5[298]}
   );
   gpc1_1 gpc851 (
      {stage0_5[448]},
      {stage1_5[299]}
   );
   gpc1_1 gpc852 (
      {stage0_5[449]},
      {stage1_5[300]}
   );
   gpc1_1 gpc853 (
      {stage0_5[450]},
      {stage1_5[301]}
   );
   gpc1_1 gpc854 (
      {stage0_5[451]},
      {stage1_5[302]}
   );
   gpc1_1 gpc855 (
      {stage0_5[452]},
      {stage1_5[303]}
   );
   gpc1_1 gpc856 (
      {stage0_5[453]},
      {stage1_5[304]}
   );
   gpc1_1 gpc857 (
      {stage0_5[454]},
      {stage1_5[305]}
   );
   gpc1_1 gpc858 (
      {stage0_5[455]},
      {stage1_5[306]}
   );
   gpc1_1 gpc859 (
      {stage0_5[456]},
      {stage1_5[307]}
   );
   gpc1_1 gpc860 (
      {stage0_5[457]},
      {stage1_5[308]}
   );
   gpc1_1 gpc861 (
      {stage0_5[458]},
      {stage1_5[309]}
   );
   gpc1_1 gpc862 (
      {stage0_5[459]},
      {stage1_5[310]}
   );
   gpc1_1 gpc863 (
      {stage0_5[460]},
      {stage1_5[311]}
   );
   gpc1_1 gpc864 (
      {stage0_5[461]},
      {stage1_5[312]}
   );
   gpc1_1 gpc865 (
      {stage0_5[462]},
      {stage1_5[313]}
   );
   gpc1_1 gpc866 (
      {stage0_5[463]},
      {stage1_5[314]}
   );
   gpc1_1 gpc867 (
      {stage0_5[464]},
      {stage1_5[315]}
   );
   gpc1_1 gpc868 (
      {stage0_5[465]},
      {stage1_5[316]}
   );
   gpc1_1 gpc869 (
      {stage0_5[466]},
      {stage1_5[317]}
   );
   gpc1_1 gpc870 (
      {stage0_5[467]},
      {stage1_5[318]}
   );
   gpc1_1 gpc871 (
      {stage0_5[468]},
      {stage1_5[319]}
   );
   gpc1_1 gpc872 (
      {stage0_5[469]},
      {stage1_5[320]}
   );
   gpc1_1 gpc873 (
      {stage0_5[470]},
      {stage1_5[321]}
   );
   gpc1_1 gpc874 (
      {stage0_5[471]},
      {stage1_5[322]}
   );
   gpc1_1 gpc875 (
      {stage0_5[472]},
      {stage1_5[323]}
   );
   gpc1_1 gpc876 (
      {stage0_5[473]},
      {stage1_5[324]}
   );
   gpc1_1 gpc877 (
      {stage0_5[474]},
      {stage1_5[325]}
   );
   gpc1_1 gpc878 (
      {stage0_5[475]},
      {stage1_5[326]}
   );
   gpc1_1 gpc879 (
      {stage0_5[476]},
      {stage1_5[327]}
   );
   gpc1_1 gpc880 (
      {stage0_5[477]},
      {stage1_5[328]}
   );
   gpc1_1 gpc881 (
      {stage0_5[478]},
      {stage1_5[329]}
   );
   gpc1_1 gpc882 (
      {stage0_5[479]},
      {stage1_5[330]}
   );
   gpc1_1 gpc883 (
      {stage0_5[480]},
      {stage1_5[331]}
   );
   gpc1_1 gpc884 (
      {stage0_5[481]},
      {stage1_5[332]}
   );
   gpc1_1 gpc885 (
      {stage0_5[482]},
      {stage1_5[333]}
   );
   gpc1_1 gpc886 (
      {stage0_5[483]},
      {stage1_5[334]}
   );
   gpc1_1 gpc887 (
      {stage0_5[484]},
      {stage1_5[335]}
   );
   gpc1_1 gpc888 (
      {stage0_5[485]},
      {stage1_5[336]}
   );
   gpc1_1 gpc889 (
      {stage0_6[457]},
      {stage1_6[168]}
   );
   gpc1_1 gpc890 (
      {stage0_6[458]},
      {stage1_6[169]}
   );
   gpc1_1 gpc891 (
      {stage0_6[459]},
      {stage1_6[170]}
   );
   gpc1_1 gpc892 (
      {stage0_6[460]},
      {stage1_6[171]}
   );
   gpc1_1 gpc893 (
      {stage0_6[461]},
      {stage1_6[172]}
   );
   gpc1_1 gpc894 (
      {stage0_6[462]},
      {stage1_6[173]}
   );
   gpc1_1 gpc895 (
      {stage0_6[463]},
      {stage1_6[174]}
   );
   gpc1_1 gpc896 (
      {stage0_6[464]},
      {stage1_6[175]}
   );
   gpc1_1 gpc897 (
      {stage0_6[465]},
      {stage1_6[176]}
   );
   gpc1_1 gpc898 (
      {stage0_6[466]},
      {stage1_6[177]}
   );
   gpc1_1 gpc899 (
      {stage0_6[467]},
      {stage1_6[178]}
   );
   gpc1_1 gpc900 (
      {stage0_6[468]},
      {stage1_6[179]}
   );
   gpc1_1 gpc901 (
      {stage0_6[469]},
      {stage1_6[180]}
   );
   gpc1_1 gpc902 (
      {stage0_6[470]},
      {stage1_6[181]}
   );
   gpc1_1 gpc903 (
      {stage0_6[471]},
      {stage1_6[182]}
   );
   gpc1_1 gpc904 (
      {stage0_6[472]},
      {stage1_6[183]}
   );
   gpc1_1 gpc905 (
      {stage0_6[473]},
      {stage1_6[184]}
   );
   gpc1_1 gpc906 (
      {stage0_6[474]},
      {stage1_6[185]}
   );
   gpc1_1 gpc907 (
      {stage0_6[475]},
      {stage1_6[186]}
   );
   gpc1_1 gpc908 (
      {stage0_6[476]},
      {stage1_6[187]}
   );
   gpc1_1 gpc909 (
      {stage0_6[477]},
      {stage1_6[188]}
   );
   gpc1_1 gpc910 (
      {stage0_6[478]},
      {stage1_6[189]}
   );
   gpc1_1 gpc911 (
      {stage0_6[479]},
      {stage1_6[190]}
   );
   gpc1_1 gpc912 (
      {stage0_6[480]},
      {stage1_6[191]}
   );
   gpc1_1 gpc913 (
      {stage0_6[481]},
      {stage1_6[192]}
   );
   gpc1_1 gpc914 (
      {stage0_6[482]},
      {stage1_6[193]}
   );
   gpc1_1 gpc915 (
      {stage0_6[483]},
      {stage1_6[194]}
   );
   gpc1_1 gpc916 (
      {stage0_6[484]},
      {stage1_6[195]}
   );
   gpc1_1 gpc917 (
      {stage0_6[485]},
      {stage1_6[196]}
   );
   gpc1_1 gpc918 (
      {stage0_7[425]},
      {stage1_7[156]}
   );
   gpc1_1 gpc919 (
      {stage0_7[426]},
      {stage1_7[157]}
   );
   gpc1_1 gpc920 (
      {stage0_7[427]},
      {stage1_7[158]}
   );
   gpc1_1 gpc921 (
      {stage0_7[428]},
      {stage1_7[159]}
   );
   gpc1_1 gpc922 (
      {stage0_7[429]},
      {stage1_7[160]}
   );
   gpc1_1 gpc923 (
      {stage0_7[430]},
      {stage1_7[161]}
   );
   gpc1_1 gpc924 (
      {stage0_7[431]},
      {stage1_7[162]}
   );
   gpc1_1 gpc925 (
      {stage0_7[432]},
      {stage1_7[163]}
   );
   gpc1_1 gpc926 (
      {stage0_7[433]},
      {stage1_7[164]}
   );
   gpc1_1 gpc927 (
      {stage0_7[434]},
      {stage1_7[165]}
   );
   gpc1_1 gpc928 (
      {stage0_7[435]},
      {stage1_7[166]}
   );
   gpc1_1 gpc929 (
      {stage0_7[436]},
      {stage1_7[167]}
   );
   gpc1_1 gpc930 (
      {stage0_7[437]},
      {stage1_7[168]}
   );
   gpc1_1 gpc931 (
      {stage0_7[438]},
      {stage1_7[169]}
   );
   gpc1_1 gpc932 (
      {stage0_7[439]},
      {stage1_7[170]}
   );
   gpc1_1 gpc933 (
      {stage0_7[440]},
      {stage1_7[171]}
   );
   gpc1_1 gpc934 (
      {stage0_7[441]},
      {stage1_7[172]}
   );
   gpc1_1 gpc935 (
      {stage0_7[442]},
      {stage1_7[173]}
   );
   gpc1_1 gpc936 (
      {stage0_7[443]},
      {stage1_7[174]}
   );
   gpc1_1 gpc937 (
      {stage0_7[444]},
      {stage1_7[175]}
   );
   gpc1_1 gpc938 (
      {stage0_7[445]},
      {stage1_7[176]}
   );
   gpc1_1 gpc939 (
      {stage0_7[446]},
      {stage1_7[177]}
   );
   gpc1_1 gpc940 (
      {stage0_7[447]},
      {stage1_7[178]}
   );
   gpc1_1 gpc941 (
      {stage0_7[448]},
      {stage1_7[179]}
   );
   gpc1_1 gpc942 (
      {stage0_7[449]},
      {stage1_7[180]}
   );
   gpc1_1 gpc943 (
      {stage0_7[450]},
      {stage1_7[181]}
   );
   gpc1_1 gpc944 (
      {stage0_7[451]},
      {stage1_7[182]}
   );
   gpc1_1 gpc945 (
      {stage0_7[452]},
      {stage1_7[183]}
   );
   gpc1_1 gpc946 (
      {stage0_7[453]},
      {stage1_7[184]}
   );
   gpc1_1 gpc947 (
      {stage0_7[454]},
      {stage1_7[185]}
   );
   gpc1_1 gpc948 (
      {stage0_7[455]},
      {stage1_7[186]}
   );
   gpc1_1 gpc949 (
      {stage0_7[456]},
      {stage1_7[187]}
   );
   gpc1_1 gpc950 (
      {stage0_7[457]},
      {stage1_7[188]}
   );
   gpc1_1 gpc951 (
      {stage0_7[458]},
      {stage1_7[189]}
   );
   gpc1_1 gpc952 (
      {stage0_7[459]},
      {stage1_7[190]}
   );
   gpc1_1 gpc953 (
      {stage0_7[460]},
      {stage1_7[191]}
   );
   gpc1_1 gpc954 (
      {stage0_7[461]},
      {stage1_7[192]}
   );
   gpc1_1 gpc955 (
      {stage0_7[462]},
      {stage1_7[193]}
   );
   gpc1_1 gpc956 (
      {stage0_7[463]},
      {stage1_7[194]}
   );
   gpc1_1 gpc957 (
      {stage0_7[464]},
      {stage1_7[195]}
   );
   gpc1_1 gpc958 (
      {stage0_7[465]},
      {stage1_7[196]}
   );
   gpc1_1 gpc959 (
      {stage0_7[466]},
      {stage1_7[197]}
   );
   gpc1_1 gpc960 (
      {stage0_7[467]},
      {stage1_7[198]}
   );
   gpc1_1 gpc961 (
      {stage0_7[468]},
      {stage1_7[199]}
   );
   gpc1_1 gpc962 (
      {stage0_7[469]},
      {stage1_7[200]}
   );
   gpc1_1 gpc963 (
      {stage0_7[470]},
      {stage1_7[201]}
   );
   gpc1_1 gpc964 (
      {stage0_7[471]},
      {stage1_7[202]}
   );
   gpc1_1 gpc965 (
      {stage0_7[472]},
      {stage1_7[203]}
   );
   gpc1_1 gpc966 (
      {stage0_7[473]},
      {stage1_7[204]}
   );
   gpc1_1 gpc967 (
      {stage0_7[474]},
      {stage1_7[205]}
   );
   gpc1_1 gpc968 (
      {stage0_7[475]},
      {stage1_7[206]}
   );
   gpc1_1 gpc969 (
      {stage0_7[476]},
      {stage1_7[207]}
   );
   gpc1_1 gpc970 (
      {stage0_7[477]},
      {stage1_7[208]}
   );
   gpc1_1 gpc971 (
      {stage0_7[478]},
      {stage1_7[209]}
   );
   gpc1_1 gpc972 (
      {stage0_7[479]},
      {stage1_7[210]}
   );
   gpc1_1 gpc973 (
      {stage0_7[480]},
      {stage1_7[211]}
   );
   gpc1_1 gpc974 (
      {stage0_7[481]},
      {stage1_7[212]}
   );
   gpc1_1 gpc975 (
      {stage0_7[482]},
      {stage1_7[213]}
   );
   gpc1_1 gpc976 (
      {stage0_7[483]},
      {stage1_7[214]}
   );
   gpc1_1 gpc977 (
      {stage0_7[484]},
      {stage1_7[215]}
   );
   gpc1_1 gpc978 (
      {stage0_7[485]},
      {stage1_7[216]}
   );
   gpc1_1 gpc979 (
      {stage0_10[381]},
      {stage1_10[177]}
   );
   gpc1_1 gpc980 (
      {stage0_10[382]},
      {stage1_10[178]}
   );
   gpc1_1 gpc981 (
      {stage0_10[383]},
      {stage1_10[179]}
   );
   gpc1_1 gpc982 (
      {stage0_10[384]},
      {stage1_10[180]}
   );
   gpc1_1 gpc983 (
      {stage0_10[385]},
      {stage1_10[181]}
   );
   gpc1_1 gpc984 (
      {stage0_10[386]},
      {stage1_10[182]}
   );
   gpc1_1 gpc985 (
      {stage0_10[387]},
      {stage1_10[183]}
   );
   gpc1_1 gpc986 (
      {stage0_10[388]},
      {stage1_10[184]}
   );
   gpc1_1 gpc987 (
      {stage0_10[389]},
      {stage1_10[185]}
   );
   gpc1_1 gpc988 (
      {stage0_10[390]},
      {stage1_10[186]}
   );
   gpc1_1 gpc989 (
      {stage0_10[391]},
      {stage1_10[187]}
   );
   gpc1_1 gpc990 (
      {stage0_10[392]},
      {stage1_10[188]}
   );
   gpc1_1 gpc991 (
      {stage0_10[393]},
      {stage1_10[189]}
   );
   gpc1_1 gpc992 (
      {stage0_10[394]},
      {stage1_10[190]}
   );
   gpc1_1 gpc993 (
      {stage0_10[395]},
      {stage1_10[191]}
   );
   gpc1_1 gpc994 (
      {stage0_10[396]},
      {stage1_10[192]}
   );
   gpc1_1 gpc995 (
      {stage0_10[397]},
      {stage1_10[193]}
   );
   gpc1_1 gpc996 (
      {stage0_10[398]},
      {stage1_10[194]}
   );
   gpc1_1 gpc997 (
      {stage0_10[399]},
      {stage1_10[195]}
   );
   gpc1_1 gpc998 (
      {stage0_10[400]},
      {stage1_10[196]}
   );
   gpc1_1 gpc999 (
      {stage0_10[401]},
      {stage1_10[197]}
   );
   gpc1_1 gpc1000 (
      {stage0_10[402]},
      {stage1_10[198]}
   );
   gpc1_1 gpc1001 (
      {stage0_10[403]},
      {stage1_10[199]}
   );
   gpc1_1 gpc1002 (
      {stage0_10[404]},
      {stage1_10[200]}
   );
   gpc1_1 gpc1003 (
      {stage0_10[405]},
      {stage1_10[201]}
   );
   gpc1_1 gpc1004 (
      {stage0_10[406]},
      {stage1_10[202]}
   );
   gpc1_1 gpc1005 (
      {stage0_10[407]},
      {stage1_10[203]}
   );
   gpc1_1 gpc1006 (
      {stage0_10[408]},
      {stage1_10[204]}
   );
   gpc1_1 gpc1007 (
      {stage0_10[409]},
      {stage1_10[205]}
   );
   gpc1_1 gpc1008 (
      {stage0_10[410]},
      {stage1_10[206]}
   );
   gpc1_1 gpc1009 (
      {stage0_10[411]},
      {stage1_10[207]}
   );
   gpc1_1 gpc1010 (
      {stage0_10[412]},
      {stage1_10[208]}
   );
   gpc1_1 gpc1011 (
      {stage0_10[413]},
      {stage1_10[209]}
   );
   gpc1_1 gpc1012 (
      {stage0_10[414]},
      {stage1_10[210]}
   );
   gpc1_1 gpc1013 (
      {stage0_10[415]},
      {stage1_10[211]}
   );
   gpc1_1 gpc1014 (
      {stage0_10[416]},
      {stage1_10[212]}
   );
   gpc1_1 gpc1015 (
      {stage0_10[417]},
      {stage1_10[213]}
   );
   gpc1_1 gpc1016 (
      {stage0_10[418]},
      {stage1_10[214]}
   );
   gpc1_1 gpc1017 (
      {stage0_10[419]},
      {stage1_10[215]}
   );
   gpc1_1 gpc1018 (
      {stage0_10[420]},
      {stage1_10[216]}
   );
   gpc1_1 gpc1019 (
      {stage0_10[421]},
      {stage1_10[217]}
   );
   gpc1_1 gpc1020 (
      {stage0_10[422]},
      {stage1_10[218]}
   );
   gpc1_1 gpc1021 (
      {stage0_10[423]},
      {stage1_10[219]}
   );
   gpc1_1 gpc1022 (
      {stage0_10[424]},
      {stage1_10[220]}
   );
   gpc1_1 gpc1023 (
      {stage0_10[425]},
      {stage1_10[221]}
   );
   gpc1_1 gpc1024 (
      {stage0_10[426]},
      {stage1_10[222]}
   );
   gpc1_1 gpc1025 (
      {stage0_10[427]},
      {stage1_10[223]}
   );
   gpc1_1 gpc1026 (
      {stage0_10[428]},
      {stage1_10[224]}
   );
   gpc1_1 gpc1027 (
      {stage0_10[429]},
      {stage1_10[225]}
   );
   gpc1_1 gpc1028 (
      {stage0_10[430]},
      {stage1_10[226]}
   );
   gpc1_1 gpc1029 (
      {stage0_10[431]},
      {stage1_10[227]}
   );
   gpc1_1 gpc1030 (
      {stage0_10[432]},
      {stage1_10[228]}
   );
   gpc1_1 gpc1031 (
      {stage0_10[433]},
      {stage1_10[229]}
   );
   gpc1_1 gpc1032 (
      {stage0_10[434]},
      {stage1_10[230]}
   );
   gpc1_1 gpc1033 (
      {stage0_10[435]},
      {stage1_10[231]}
   );
   gpc1_1 gpc1034 (
      {stage0_10[436]},
      {stage1_10[232]}
   );
   gpc1_1 gpc1035 (
      {stage0_10[437]},
      {stage1_10[233]}
   );
   gpc1_1 gpc1036 (
      {stage0_10[438]},
      {stage1_10[234]}
   );
   gpc1_1 gpc1037 (
      {stage0_10[439]},
      {stage1_10[235]}
   );
   gpc1_1 gpc1038 (
      {stage0_10[440]},
      {stage1_10[236]}
   );
   gpc1_1 gpc1039 (
      {stage0_10[441]},
      {stage1_10[237]}
   );
   gpc1_1 gpc1040 (
      {stage0_10[442]},
      {stage1_10[238]}
   );
   gpc1_1 gpc1041 (
      {stage0_10[443]},
      {stage1_10[239]}
   );
   gpc1_1 gpc1042 (
      {stage0_10[444]},
      {stage1_10[240]}
   );
   gpc1_1 gpc1043 (
      {stage0_10[445]},
      {stage1_10[241]}
   );
   gpc1_1 gpc1044 (
      {stage0_10[446]},
      {stage1_10[242]}
   );
   gpc1_1 gpc1045 (
      {stage0_10[447]},
      {stage1_10[243]}
   );
   gpc1_1 gpc1046 (
      {stage0_10[448]},
      {stage1_10[244]}
   );
   gpc1_1 gpc1047 (
      {stage0_10[449]},
      {stage1_10[245]}
   );
   gpc1_1 gpc1048 (
      {stage0_10[450]},
      {stage1_10[246]}
   );
   gpc1_1 gpc1049 (
      {stage0_10[451]},
      {stage1_10[247]}
   );
   gpc1_1 gpc1050 (
      {stage0_10[452]},
      {stage1_10[248]}
   );
   gpc1_1 gpc1051 (
      {stage0_10[453]},
      {stage1_10[249]}
   );
   gpc1_1 gpc1052 (
      {stage0_10[454]},
      {stage1_10[250]}
   );
   gpc1_1 gpc1053 (
      {stage0_10[455]},
      {stage1_10[251]}
   );
   gpc1_1 gpc1054 (
      {stage0_10[456]},
      {stage1_10[252]}
   );
   gpc1_1 gpc1055 (
      {stage0_10[457]},
      {stage1_10[253]}
   );
   gpc1_1 gpc1056 (
      {stage0_10[458]},
      {stage1_10[254]}
   );
   gpc1_1 gpc1057 (
      {stage0_10[459]},
      {stage1_10[255]}
   );
   gpc1_1 gpc1058 (
      {stage0_10[460]},
      {stage1_10[256]}
   );
   gpc1_1 gpc1059 (
      {stage0_10[461]},
      {stage1_10[257]}
   );
   gpc1_1 gpc1060 (
      {stage0_10[462]},
      {stage1_10[258]}
   );
   gpc1_1 gpc1061 (
      {stage0_10[463]},
      {stage1_10[259]}
   );
   gpc1_1 gpc1062 (
      {stage0_10[464]},
      {stage1_10[260]}
   );
   gpc1_1 gpc1063 (
      {stage0_10[465]},
      {stage1_10[261]}
   );
   gpc1_1 gpc1064 (
      {stage0_10[466]},
      {stage1_10[262]}
   );
   gpc1_1 gpc1065 (
      {stage0_10[467]},
      {stage1_10[263]}
   );
   gpc1_1 gpc1066 (
      {stage0_10[468]},
      {stage1_10[264]}
   );
   gpc1_1 gpc1067 (
      {stage0_10[469]},
      {stage1_10[265]}
   );
   gpc1_1 gpc1068 (
      {stage0_10[470]},
      {stage1_10[266]}
   );
   gpc1_1 gpc1069 (
      {stage0_10[471]},
      {stage1_10[267]}
   );
   gpc1_1 gpc1070 (
      {stage0_10[472]},
      {stage1_10[268]}
   );
   gpc1_1 gpc1071 (
      {stage0_10[473]},
      {stage1_10[269]}
   );
   gpc1_1 gpc1072 (
      {stage0_10[474]},
      {stage1_10[270]}
   );
   gpc1_1 gpc1073 (
      {stage0_10[475]},
      {stage1_10[271]}
   );
   gpc1_1 gpc1074 (
      {stage0_10[476]},
      {stage1_10[272]}
   );
   gpc1_1 gpc1075 (
      {stage0_10[477]},
      {stage1_10[273]}
   );
   gpc1_1 gpc1076 (
      {stage0_10[478]},
      {stage1_10[274]}
   );
   gpc1_1 gpc1077 (
      {stage0_10[479]},
      {stage1_10[275]}
   );
   gpc1_1 gpc1078 (
      {stage0_10[480]},
      {stage1_10[276]}
   );
   gpc1_1 gpc1079 (
      {stage0_10[481]},
      {stage1_10[277]}
   );
   gpc1_1 gpc1080 (
      {stage0_10[482]},
      {stage1_10[278]}
   );
   gpc1_1 gpc1081 (
      {stage0_10[483]},
      {stage1_10[279]}
   );
   gpc1_1 gpc1082 (
      {stage0_10[484]},
      {stage1_10[280]}
   );
   gpc1_1 gpc1083 (
      {stage0_10[485]},
      {stage1_10[281]}
   );
   gpc1_1 gpc1084 (
      {stage0_11[423]},
      {stage1_11[151]}
   );
   gpc1_1 gpc1085 (
      {stage0_11[424]},
      {stage1_11[152]}
   );
   gpc1_1 gpc1086 (
      {stage0_11[425]},
      {stage1_11[153]}
   );
   gpc1_1 gpc1087 (
      {stage0_11[426]},
      {stage1_11[154]}
   );
   gpc1_1 gpc1088 (
      {stage0_11[427]},
      {stage1_11[155]}
   );
   gpc1_1 gpc1089 (
      {stage0_11[428]},
      {stage1_11[156]}
   );
   gpc1_1 gpc1090 (
      {stage0_11[429]},
      {stage1_11[157]}
   );
   gpc1_1 gpc1091 (
      {stage0_11[430]},
      {stage1_11[158]}
   );
   gpc1_1 gpc1092 (
      {stage0_11[431]},
      {stage1_11[159]}
   );
   gpc1_1 gpc1093 (
      {stage0_11[432]},
      {stage1_11[160]}
   );
   gpc1_1 gpc1094 (
      {stage0_11[433]},
      {stage1_11[161]}
   );
   gpc1_1 gpc1095 (
      {stage0_11[434]},
      {stage1_11[162]}
   );
   gpc1_1 gpc1096 (
      {stage0_11[435]},
      {stage1_11[163]}
   );
   gpc1_1 gpc1097 (
      {stage0_11[436]},
      {stage1_11[164]}
   );
   gpc1_1 gpc1098 (
      {stage0_11[437]},
      {stage1_11[165]}
   );
   gpc1_1 gpc1099 (
      {stage0_11[438]},
      {stage1_11[166]}
   );
   gpc1_1 gpc1100 (
      {stage0_11[439]},
      {stage1_11[167]}
   );
   gpc1_1 gpc1101 (
      {stage0_11[440]},
      {stage1_11[168]}
   );
   gpc1_1 gpc1102 (
      {stage0_11[441]},
      {stage1_11[169]}
   );
   gpc1_1 gpc1103 (
      {stage0_11[442]},
      {stage1_11[170]}
   );
   gpc1_1 gpc1104 (
      {stage0_11[443]},
      {stage1_11[171]}
   );
   gpc1_1 gpc1105 (
      {stage0_11[444]},
      {stage1_11[172]}
   );
   gpc1_1 gpc1106 (
      {stage0_11[445]},
      {stage1_11[173]}
   );
   gpc1_1 gpc1107 (
      {stage0_11[446]},
      {stage1_11[174]}
   );
   gpc1_1 gpc1108 (
      {stage0_11[447]},
      {stage1_11[175]}
   );
   gpc1_1 gpc1109 (
      {stage0_11[448]},
      {stage1_11[176]}
   );
   gpc1_1 gpc1110 (
      {stage0_11[449]},
      {stage1_11[177]}
   );
   gpc1_1 gpc1111 (
      {stage0_11[450]},
      {stage1_11[178]}
   );
   gpc1_1 gpc1112 (
      {stage0_11[451]},
      {stage1_11[179]}
   );
   gpc1_1 gpc1113 (
      {stage0_11[452]},
      {stage1_11[180]}
   );
   gpc1_1 gpc1114 (
      {stage0_11[453]},
      {stage1_11[181]}
   );
   gpc1_1 gpc1115 (
      {stage0_11[454]},
      {stage1_11[182]}
   );
   gpc1_1 gpc1116 (
      {stage0_11[455]},
      {stage1_11[183]}
   );
   gpc1_1 gpc1117 (
      {stage0_11[456]},
      {stage1_11[184]}
   );
   gpc1_1 gpc1118 (
      {stage0_11[457]},
      {stage1_11[185]}
   );
   gpc1_1 gpc1119 (
      {stage0_11[458]},
      {stage1_11[186]}
   );
   gpc1_1 gpc1120 (
      {stage0_11[459]},
      {stage1_11[187]}
   );
   gpc1_1 gpc1121 (
      {stage0_11[460]},
      {stage1_11[188]}
   );
   gpc1_1 gpc1122 (
      {stage0_11[461]},
      {stage1_11[189]}
   );
   gpc1_1 gpc1123 (
      {stage0_11[462]},
      {stage1_11[190]}
   );
   gpc1_1 gpc1124 (
      {stage0_11[463]},
      {stage1_11[191]}
   );
   gpc1_1 gpc1125 (
      {stage0_11[464]},
      {stage1_11[192]}
   );
   gpc1_1 gpc1126 (
      {stage0_11[465]},
      {stage1_11[193]}
   );
   gpc1_1 gpc1127 (
      {stage0_11[466]},
      {stage1_11[194]}
   );
   gpc1_1 gpc1128 (
      {stage0_11[467]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1129 (
      {stage0_11[468]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1130 (
      {stage0_11[469]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1131 (
      {stage0_11[470]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1132 (
      {stage0_11[471]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1133 (
      {stage0_11[472]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1134 (
      {stage0_11[473]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1135 (
      {stage0_11[474]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1136 (
      {stage0_11[475]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1137 (
      {stage0_11[476]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1138 (
      {stage0_11[477]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1139 (
      {stage0_11[478]},
      {stage1_11[206]}
   );
   gpc1_1 gpc1140 (
      {stage0_11[479]},
      {stage1_11[207]}
   );
   gpc1_1 gpc1141 (
      {stage0_11[480]},
      {stage1_11[208]}
   );
   gpc1_1 gpc1142 (
      {stage0_11[481]},
      {stage1_11[209]}
   );
   gpc1_1 gpc1143 (
      {stage0_11[482]},
      {stage1_11[210]}
   );
   gpc1_1 gpc1144 (
      {stage0_11[483]},
      {stage1_11[211]}
   );
   gpc1_1 gpc1145 (
      {stage0_11[484]},
      {stage1_11[212]}
   );
   gpc1_1 gpc1146 (
      {stage0_11[485]},
      {stage1_11[213]}
   );
   gpc1_1 gpc1147 (
      {stage0_14[474]},
      {stage1_14[171]}
   );
   gpc1_1 gpc1148 (
      {stage0_14[475]},
      {stage1_14[172]}
   );
   gpc1_1 gpc1149 (
      {stage0_14[476]},
      {stage1_14[173]}
   );
   gpc1_1 gpc1150 (
      {stage0_14[477]},
      {stage1_14[174]}
   );
   gpc1_1 gpc1151 (
      {stage0_14[478]},
      {stage1_14[175]}
   );
   gpc1_1 gpc1152 (
      {stage0_14[479]},
      {stage1_14[176]}
   );
   gpc1_1 gpc1153 (
      {stage0_14[480]},
      {stage1_14[177]}
   );
   gpc1_1 gpc1154 (
      {stage0_14[481]},
      {stage1_14[178]}
   );
   gpc1_1 gpc1155 (
      {stage0_14[482]},
      {stage1_14[179]}
   );
   gpc1_1 gpc1156 (
      {stage0_14[483]},
      {stage1_14[180]}
   );
   gpc1_1 gpc1157 (
      {stage0_14[484]},
      {stage1_14[181]}
   );
   gpc1_1 gpc1158 (
      {stage0_14[485]},
      {stage1_14[182]}
   );
   gpc1163_5 gpc1159 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1160 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1161 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1162 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1163 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1164 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1165 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1166 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1167 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1168 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc1169 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc1170 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc1171 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1172 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc1173 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc1174 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc1175 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc1176 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc1177 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc1178 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc1179 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc1180 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101]},
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc1181 (
      {stage1_0[102], stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106], stage1_0[107]},
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc1182 (
      {stage1_0[108], stage1_0[109], stage1_0[110], stage1_0[111], stage1_0[112], stage1_0[113]},
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93]},
      {stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23],stage2_0[23]}
   );
   gpc606_5 gpc1183 (
      {stage1_0[114], stage1_0[115], stage1_0[116], stage1_0[117], stage1_0[118], stage1_0[119]},
      {stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99]},
      {stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24],stage2_0[24]}
   );
   gpc606_5 gpc1184 (
      {stage1_0[120], stage1_0[121], stage1_0[122], stage1_0[123], stage1_0[124], stage1_0[125]},
      {stage1_2[100], stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25],stage2_0[25]}
   );
   gpc606_5 gpc1185 (
      {stage1_0[126], stage1_0[127], stage1_0[128], stage1_0[129], stage1_0[130], stage1_0[131]},
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26],stage2_0[26]}
   );
   gpc606_5 gpc1186 (
      {stage1_0[132], stage1_0[133], stage1_0[134], stage1_0[135], stage1_0[136], stage1_0[137]},
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27],stage2_0[27]}
   );
   gpc606_5 gpc1187 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15]},
      {stage2_5[0],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc1188 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage2_5[1],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc1189 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage2_5[2],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc1190 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage2_5[3],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc1191 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage2_5[4],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc1192 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage2_5[5],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc1193 (
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage2_5[6],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc1194 (
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage2_5[7],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc615_5 gpc1195 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[58]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[8],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc1196 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[59]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[9],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc615_5 gpc1197 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[60]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[10],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc615_5 gpc1198 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[61]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[11],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc1199 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[62]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[12],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc1200 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[63]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[13],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc1201 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[64]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[14],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc1202 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[65]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[15],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc1203 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[16],stage2_4[44],stage2_3[44]}
   );
   gpc615_5 gpc1204 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[17],stage2_4[45],stage2_3[45]}
   );
   gpc615_5 gpc1205 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[50]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[10],stage2_5[18],stage2_4[46],stage2_3[46]}
   );
   gpc615_5 gpc1206 (
      {stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage1_4[51]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[11],stage2_5[19],stage2_4[47],stage2_3[47]}
   );
   gpc615_5 gpc1207 (
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90]},
      {stage1_4[52]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[12],stage2_5[20],stage2_4[48],stage2_3[48]}
   );
   gpc615_5 gpc1208 (
      {stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage1_4[53]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[13],stage2_5[21],stage2_4[49],stage2_3[49]}
   );
   gpc615_5 gpc1209 (
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100]},
      {stage1_4[54]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[14],stage2_5[22],stage2_4[50],stage2_3[50]}
   );
   gpc615_5 gpc1210 (
      {stage1_3[101], stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105]},
      {stage1_4[55]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[15],stage2_5[23],stage2_4[51],stage2_3[51]}
   );
   gpc615_5 gpc1211 (
      {stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109], stage1_3[110]},
      {stage1_4[56]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[16],stage2_5[24],stage2_4[52],stage2_3[52]}
   );
   gpc615_5 gpc1212 (
      {stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage1_4[57]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[17],stage2_5[25],stage2_4[53],stage2_3[53]}
   );
   gpc615_5 gpc1213 (
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120]},
      {stage1_4[58]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[18],stage2_5[26],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc1214 (
      {stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage1_4[59]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[19],stage2_5[27],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc1215 (
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130]},
      {stage1_4[60]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[20],stage2_5[28],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc1216 (
      {stage1_3[131], stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[61]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[21],stage2_5[29],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc1217 (
      {stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139], stage1_3[140]},
      {stage1_4[62]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[22],stage2_5[30],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc1218 (
      {stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage1_4[63]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[23],stage2_5[31],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc1219 (
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150]},
      {stage1_4[64]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[24],stage2_5[32],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc1220 (
      {stage1_3[151], stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155]},
      {stage1_4[65]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[25],stage2_5[33],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc1221 (
      {stage1_3[156], stage1_3[157], stage1_3[158], stage1_3[159], stage1_3[160]},
      {stage1_4[66]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[26],stage2_5[34],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc1222 (
      {stage1_3[161], stage1_3[162], stage1_3[163], stage1_3[164], stage1_3[165]},
      {stage1_4[67]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[27],stage2_5[35],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc1223 (
      {stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169], stage1_3[170]},
      {stage1_4[68]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[28],stage2_5[36],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc1224 (
      {stage1_3[171], stage1_3[172], stage1_3[173], stage1_3[174], stage1_3[175]},
      {stage1_4[69]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage2_7[21],stage2_6[29],stage2_5[37],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc1225 (
      {stage1_3[176], stage1_3[177], stage1_3[178], stage1_3[179], stage1_3[180]},
      {stage1_4[70]},
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage2_7[22],stage2_6[30],stage2_5[38],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc1226 (
      {stage1_3[181], stage1_3[182], stage1_3[183], stage1_3[184], stage1_3[185]},
      {stage1_4[71]},
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage2_7[23],stage2_6[31],stage2_5[39],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc1227 (
      {stage1_3[186], stage1_3[187], stage1_3[188], stage1_3[189], stage1_3[190]},
      {stage1_4[72]},
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage2_7[24],stage2_6[32],stage2_5[40],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc1228 (
      {stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194], stage1_3[195]},
      {stage1_4[73]},
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage2_7[25],stage2_6[33],stage2_5[41],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc1229 (
      {stage1_3[196], stage1_3[197], stage1_3[198], stage1_3[199], stage1_3[200]},
      {stage1_4[74]},
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage2_7[26],stage2_6[34],stage2_5[42],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc1230 (
      {stage1_3[201], stage1_3[202], stage1_3[203], stage1_3[204], stage1_3[205]},
      {stage1_4[75]},
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage2_7[27],stage2_6[35],stage2_5[43],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc1231 (
      {stage1_3[206], stage1_3[207], stage1_3[208], stage1_3[209], stage1_3[210]},
      {stage1_4[76]},
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage2_7[28],stage2_6[36],stage2_5[44],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc1232 (
      {stage1_3[211], stage1_3[212], stage1_3[213], stage1_3[214], stage1_3[215]},
      {stage1_4[77]},
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage2_7[29],stage2_6[37],stage2_5[45],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc1233 (
      {stage1_3[216], stage1_3[217], stage1_3[218], stage1_3[219], stage1_3[220]},
      {stage1_4[78]},
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage2_7[30],stage2_6[38],stage2_5[46],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc1234 (
      {stage1_3[221], stage1_3[222], stage1_3[223], stage1_3[224], stage1_3[225]},
      {stage1_4[79]},
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage2_7[31],stage2_6[39],stage2_5[47],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc1235 (
      {stage1_3[226], stage1_3[227], stage1_3[228], stage1_3[229], stage1_3[230]},
      {stage1_4[80]},
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage2_7[32],stage2_6[40],stage2_5[48],stage2_4[76],stage2_3[76]}
   );
   gpc615_5 gpc1236 (
      {stage1_3[231], stage1_3[232], stage1_3[233], stage1_3[234], stage1_3[235]},
      {stage1_4[81]},
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage2_7[33],stage2_6[41],stage2_5[49],stage2_4[77],stage2_3[77]}
   );
   gpc615_5 gpc1237 (
      {stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_5[204]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[34],stage2_6[42],stage2_5[50],stage2_4[78]}
   );
   gpc615_5 gpc1238 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_5[205]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[35],stage2_6[43],stage2_5[51],stage2_4[79]}
   );
   gpc615_5 gpc1239 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96]},
      {stage1_5[206]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[36],stage2_6[44],stage2_5[52],stage2_4[80]}
   );
   gpc615_5 gpc1240 (
      {stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_5[207]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[37],stage2_6[45],stage2_5[53],stage2_4[81]}
   );
   gpc615_5 gpc1241 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_5[208]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[38],stage2_6[46],stage2_5[54],stage2_4[82]}
   );
   gpc615_5 gpc1242 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111]},
      {stage1_5[209]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[39],stage2_6[47],stage2_5[55],stage2_4[83]}
   );
   gpc615_5 gpc1243 (
      {stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_5[210]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[40],stage2_6[48],stage2_5[56],stage2_4[84]}
   );
   gpc615_5 gpc1244 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_5[211]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[41],stage2_6[49],stage2_5[57],stage2_4[85]}
   );
   gpc615_5 gpc1245 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126]},
      {stage1_5[212]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[42],stage2_6[50],stage2_5[58],stage2_4[86]}
   );
   gpc615_5 gpc1246 (
      {stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130], stage1_4[131]},
      {stage1_5[213]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[43],stage2_6[51],stage2_5[59],stage2_4[87]}
   );
   gpc615_5 gpc1247 (
      {stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135], stage1_4[136]},
      {stage1_5[214]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[44],stage2_6[52],stage2_5[60],stage2_4[88]}
   );
   gpc615_5 gpc1248 (
      {stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141]},
      {stage1_5[215]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[45],stage2_6[53],stage2_5[61],stage2_4[89]}
   );
   gpc615_5 gpc1249 (
      {stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_5[216]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[46],stage2_6[54],stage2_5[62],stage2_4[90]}
   );
   gpc615_5 gpc1250 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151]},
      {stage1_5[217]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[47],stage2_6[55],stage2_5[63],stage2_4[91]}
   );
   gpc615_5 gpc1251 (
      {stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156]},
      {stage1_5[218]},
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage2_8[14],stage2_7[48],stage2_6[56],stage2_5[64],stage2_4[92]}
   );
   gpc615_5 gpc1252 (
      {stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161]},
      {stage1_5[219]},
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage2_8[15],stage2_7[49],stage2_6[57],stage2_5[65],stage2_4[93]}
   );
   gpc615_5 gpc1253 (
      {stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166]},
      {stage1_5[220]},
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage2_8[16],stage2_7[50],stage2_6[58],stage2_5[66],stage2_4[94]}
   );
   gpc615_5 gpc1254 (
      {stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171]},
      {stage1_5[221]},
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage2_8[17],stage2_7[51],stage2_6[59],stage2_5[67],stage2_4[95]}
   );
   gpc615_5 gpc1255 (
      {stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_5[222]},
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage2_8[18],stage2_7[52],stage2_6[60],stage2_5[68],stage2_4[96]}
   );
   gpc615_5 gpc1256 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181]},
      {stage1_5[223]},
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage2_8[19],stage2_7[53],stage2_6[61],stage2_5[69],stage2_4[97]}
   );
   gpc615_5 gpc1257 (
      {stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186]},
      {stage1_5[224]},
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage2_8[20],stage2_7[54],stage2_6[62],stage2_5[70],stage2_4[98]}
   );
   gpc615_5 gpc1258 (
      {stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190], stage1_4[191]},
      {stage1_5[225]},
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage2_8[21],stage2_7[55],stage2_6[63],stage2_5[71],stage2_4[99]}
   );
   gpc615_5 gpc1259 (
      {stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195], stage1_4[196]},
      {stage1_5[226]},
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage2_8[22],stage2_7[56],stage2_6[64],stage2_5[72],stage2_4[100]}
   );
   gpc615_5 gpc1260 (
      {stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200], stage1_4[201]},
      {stage1_5[227]},
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage2_8[23],stage2_7[57],stage2_6[65],stage2_5[73],stage2_4[101]}
   );
   gpc615_5 gpc1261 (
      {stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206]},
      {stage1_5[228]},
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage2_8[24],stage2_7[58],stage2_6[66],stage2_5[74],stage2_4[102]}
   );
   gpc615_5 gpc1262 (
      {stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211]},
      {stage1_5[229]},
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155]},
      {stage2_8[25],stage2_7[59],stage2_6[67],stage2_5[75],stage2_4[103]}
   );
   gpc615_5 gpc1263 (
      {stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_5[230]},
      {stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage2_8[26],stage2_7[60],stage2_6[68],stage2_5[76],stage2_4[104]}
   );
   gpc615_5 gpc1264 (
      {stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221]},
      {stage1_5[231]},
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167]},
      {stage2_8[27],stage2_7[61],stage2_6[69],stage2_5[77],stage2_4[105]}
   );
   gpc606_5 gpc1265 (
      {stage1_5[232], stage1_5[233], stage1_5[234], stage1_5[235], stage1_5[236], stage1_5[237]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[28],stage2_7[62],stage2_6[70],stage2_5[78]}
   );
   gpc606_5 gpc1266 (
      {stage1_5[238], stage1_5[239], stage1_5[240], stage1_5[241], stage1_5[242], stage1_5[243]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[29],stage2_7[63],stage2_6[71],stage2_5[79]}
   );
   gpc606_5 gpc1267 (
      {stage1_5[244], stage1_5[245], stage1_5[246], stage1_5[247], stage1_5[248], stage1_5[249]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[30],stage2_7[64],stage2_6[72],stage2_5[80]}
   );
   gpc606_5 gpc1268 (
      {stage1_5[250], stage1_5[251], stage1_5[252], stage1_5[253], stage1_5[254], stage1_5[255]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[31],stage2_7[65],stage2_6[73],stage2_5[81]}
   );
   gpc606_5 gpc1269 (
      {stage1_5[256], stage1_5[257], stage1_5[258], stage1_5[259], stage1_5[260], stage1_5[261]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[32],stage2_7[66],stage2_6[74],stage2_5[82]}
   );
   gpc606_5 gpc1270 (
      {stage1_5[262], stage1_5[263], stage1_5[264], stage1_5[265], stage1_5[266], stage1_5[267]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[33],stage2_7[67],stage2_6[75],stage2_5[83]}
   );
   gpc606_5 gpc1271 (
      {stage1_5[268], stage1_5[269], stage1_5[270], stage1_5[271], stage1_5[272], stage1_5[273]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[34],stage2_7[68],stage2_6[76],stage2_5[84]}
   );
   gpc606_5 gpc1272 (
      {stage1_5[274], stage1_5[275], stage1_5[276], stage1_5[277], stage1_5[278], stage1_5[279]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[35],stage2_7[69],stage2_6[77],stage2_5[85]}
   );
   gpc606_5 gpc1273 (
      {stage1_5[280], stage1_5[281], stage1_5[282], stage1_5[283], stage1_5[284], stage1_5[285]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[36],stage2_7[70],stage2_6[78],stage2_5[86]}
   );
   gpc606_5 gpc1274 (
      {stage1_5[286], stage1_5[287], stage1_5[288], stage1_5[289], stage1_5[290], stage1_5[291]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[37],stage2_7[71],stage2_6[79],stage2_5[87]}
   );
   gpc606_5 gpc1275 (
      {stage1_5[292], stage1_5[293], stage1_5[294], stage1_5[295], stage1_5[296], stage1_5[297]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[38],stage2_7[72],stage2_6[80],stage2_5[88]}
   );
   gpc606_5 gpc1276 (
      {stage1_5[298], stage1_5[299], stage1_5[300], stage1_5[301], stage1_5[302], stage1_5[303]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[39],stage2_7[73],stage2_6[81],stage2_5[89]}
   );
   gpc606_5 gpc1277 (
      {stage1_5[304], stage1_5[305], stage1_5[306], stage1_5[307], stage1_5[308], stage1_5[309]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[40],stage2_7[74],stage2_6[82],stage2_5[90]}
   );
   gpc606_5 gpc1278 (
      {stage1_5[310], stage1_5[311], stage1_5[312], stage1_5[313], stage1_5[314], stage1_5[315]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[41],stage2_7[75],stage2_6[83],stage2_5[91]}
   );
   gpc606_5 gpc1279 (
      {stage1_5[316], stage1_5[317], stage1_5[318], stage1_5[319], stage1_5[320], stage1_5[321]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[42],stage2_7[76],stage2_6[84],stage2_5[92]}
   );
   gpc606_5 gpc1280 (
      {stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[15],stage2_8[43],stage2_7[77],stage2_6[85]}
   );
   gpc606_5 gpc1281 (
      {stage1_6[174], stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178], stage1_6[179]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[16],stage2_8[44],stage2_7[78],stage2_6[86]}
   );
   gpc606_5 gpc1282 (
      {stage1_6[180], stage1_6[181], stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[17],stage2_8[45],stage2_7[79],stage2_6[87]}
   );
   gpc606_5 gpc1283 (
      {stage1_6[186], stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[18],stage2_8[46],stage2_7[80],stage2_6[88]}
   );
   gpc615_5 gpc1284 (
      {stage1_6[192], stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196]},
      {stage1_7[90]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[19],stage2_8[47],stage2_7[81],stage2_6[89]}
   );
   gpc606_5 gpc1285 (
      {stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[20],stage2_8[48],stage2_7[82]}
   );
   gpc606_5 gpc1286 (
      {stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101], stage1_7[102]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[21],stage2_8[49],stage2_7[83]}
   );
   gpc606_5 gpc1287 (
      {stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[22],stage2_8[50],stage2_7[84]}
   );
   gpc606_5 gpc1288 (
      {stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[23],stage2_8[51],stage2_7[85]}
   );
   gpc606_5 gpc1289 (
      {stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[24],stage2_8[52],stage2_7[86]}
   );
   gpc606_5 gpc1290 (
      {stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[25],stage2_8[53],stage2_7[87]}
   );
   gpc606_5 gpc1291 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131], stage1_7[132]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[11],stage2_9[26],stage2_8[54],stage2_7[88]}
   );
   gpc606_5 gpc1292 (
      {stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136], stage1_7[137], stage1_7[138]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[12],stage2_9[27],stage2_8[55],stage2_7[89]}
   );
   gpc606_5 gpc1293 (
      {stage1_7[139], stage1_7[140], stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[13],stage2_9[28],stage2_8[56],stage2_7[90]}
   );
   gpc606_5 gpc1294 (
      {stage1_7[145], stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[14],stage2_9[29],stage2_8[57],stage2_7[91]}
   );
   gpc606_5 gpc1295 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[15],stage2_9[30],stage2_8[58],stage2_7[92]}
   );
   gpc606_5 gpc1296 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161], stage1_7[162]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[16],stage2_9[31],stage2_8[59],stage2_7[93]}
   );
   gpc606_5 gpc1297 (
      {stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166], stage1_7[167], stage1_7[168]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[17],stage2_9[32],stage2_8[60],stage2_7[94]}
   );
   gpc606_5 gpc1298 (
      {stage1_7[169], stage1_7[170], stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[18],stage2_9[33],stage2_8[61],stage2_7[95]}
   );
   gpc606_5 gpc1299 (
      {stage1_7[175], stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[19],stage2_9[34],stage2_8[62],stage2_7[96]}
   );
   gpc606_5 gpc1300 (
      {stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[20],stage2_9[35],stage2_8[63],stage2_7[97]}
   );
   gpc606_5 gpc1301 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191], stage1_7[192]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[21],stage2_9[36],stage2_8[64],stage2_7[98]}
   );
   gpc606_5 gpc1302 (
      {stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196], stage1_7[197], stage1_7[198]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[22],stage2_9[37],stage2_8[65],stage2_7[99]}
   );
   gpc606_5 gpc1303 (
      {stage1_7[199], stage1_7[200], stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[23],stage2_9[38],stage2_8[66],stage2_7[100]}
   );
   gpc606_5 gpc1304 (
      {stage1_7[205], stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[24],stage2_9[39],stage2_8[67],stage2_7[101]}
   );
   gpc606_5 gpc1305 (
      {stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215], stage1_7[216]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[25],stage2_9[40],stage2_8[68],stage2_7[102]}
   );
   gpc606_5 gpc1306 (
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[21],stage2_10[26],stage2_9[41],stage2_8[69]}
   );
   gpc606_5 gpc1307 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[22],stage2_10[27],stage2_9[42],stage2_8[70]}
   );
   gpc606_5 gpc1308 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[23],stage2_10[28],stage2_9[43],stage2_8[71]}
   );
   gpc606_5 gpc1309 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[24],stage2_10[29],stage2_9[44],stage2_8[72]}
   );
   gpc606_5 gpc1310 (
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[25],stage2_10[30],stage2_9[45],stage2_8[73]}
   );
   gpc606_5 gpc1311 (
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[26],stage2_10[31],stage2_9[46],stage2_8[74]}
   );
   gpc606_5 gpc1312 (
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[27],stage2_10[32],stage2_9[47],stage2_8[75]}
   );
   gpc606_5 gpc1313 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[28],stage2_10[33],stage2_9[48],stage2_8[76]}
   );
   gpc606_5 gpc1314 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[29],stage2_10[34],stage2_9[49],stage2_8[77]}
   );
   gpc606_5 gpc1315 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[30],stage2_10[35],stage2_9[50],stage2_8[78]}
   );
   gpc606_5 gpc1316 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[31],stage2_10[36],stage2_9[51],stage2_8[79]}
   );
   gpc606_5 gpc1317 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[32],stage2_10[37],stage2_9[52],stage2_8[80]}
   );
   gpc606_5 gpc1318 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[33],stage2_10[38],stage2_9[53],stage2_8[81]}
   );
   gpc606_5 gpc1319 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[34],stage2_10[39],stage2_9[54],stage2_8[82]}
   );
   gpc606_5 gpc1320 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[35],stage2_10[40],stage2_9[55],stage2_8[83]}
   );
   gpc606_5 gpc1321 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[36],stage2_10[41],stage2_9[56],stage2_8[84]}
   );
   gpc606_5 gpc1322 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[37],stage2_10[42],stage2_9[57],stage2_8[85]}
   );
   gpc606_5 gpc1323 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[38],stage2_10[43],stage2_9[58],stage2_8[86]}
   );
   gpc606_5 gpc1324 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage2_12[18],stage2_11[39],stage2_10[44],stage2_9[59],stage2_8[87]}
   );
   gpc606_5 gpc1325 (
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage2_12[19],stage2_11[40],stage2_10[45],stage2_9[60],stage2_8[88]}
   );
   gpc606_5 gpc1326 (
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage2_12[20],stage2_11[41],stage2_10[46],stage2_9[61],stage2_8[89]}
   );
   gpc606_5 gpc1327 (
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage2_12[21],stage2_11[42],stage2_10[47],stage2_9[62],stage2_8[90]}
   );
   gpc606_5 gpc1328 (
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage2_12[22],stage2_11[43],stage2_10[48],stage2_9[63],stage2_8[91]}
   );
   gpc606_5 gpc1329 (
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172], stage1_8[173]},
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage2_12[23],stage2_11[44],stage2_10[49],stage2_9[64],stage2_8[92]}
   );
   gpc606_5 gpc1330 (
      {stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177], stage1_8[178], stage1_8[179]},
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage2_12[24],stage2_11[45],stage2_10[50],stage2_9[65],stage2_8[93]}
   );
   gpc615_5 gpc1331 (
      {stage1_8[180], stage1_8[181], stage1_8[182], stage1_8[183], stage1_8[184]},
      {stage1_9[126]},
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage2_12[25],stage2_11[46],stage2_10[51],stage2_9[66],stage2_8[94]}
   );
   gpc606_5 gpc1332 (
      {stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131], stage1_9[132]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[26],stage2_11[47],stage2_10[52],stage2_9[67]}
   );
   gpc606_5 gpc1333 (
      {stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137], stage1_9[138]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[27],stage2_11[48],stage2_10[53],stage2_9[68]}
   );
   gpc606_5 gpc1334 (
      {stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143], stage1_9[144]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[28],stage2_11[49],stage2_10[54],stage2_9[69]}
   );
   gpc606_5 gpc1335 (
      {stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149], stage1_9[150]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[29],stage2_11[50],stage2_10[55],stage2_9[70]}
   );
   gpc606_5 gpc1336 (
      {stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155], stage1_9[156]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[30],stage2_11[51],stage2_10[56],stage2_9[71]}
   );
   gpc606_5 gpc1337 (
      {stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161], stage1_9[162]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[31],stage2_11[52],stage2_10[57],stage2_9[72]}
   );
   gpc606_5 gpc1338 (
      {stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167], stage1_9[168]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[32],stage2_11[53],stage2_10[58],stage2_9[73]}
   );
   gpc606_5 gpc1339 (
      {stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173], stage1_9[174]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[33],stage2_11[54],stage2_10[59],stage2_9[74]}
   );
   gpc606_5 gpc1340 (
      {stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179], stage1_9[180]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[34],stage2_11[55],stage2_10[60],stage2_9[75]}
   );
   gpc606_5 gpc1341 (
      {stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185], stage1_9[186]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[35],stage2_11[56],stage2_10[61],stage2_9[76]}
   );
   gpc606_5 gpc1342 (
      {stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191], stage1_9[192]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[36],stage2_11[57],stage2_10[62],stage2_9[77]}
   );
   gpc606_5 gpc1343 (
      {stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197], stage1_9[198]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[37],stage2_11[58],stage2_10[63],stage2_9[78]}
   );
   gpc606_5 gpc1344 (
      {stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203], stage1_9[204]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[38],stage2_11[59],stage2_10[64],stage2_9[79]}
   );
   gpc606_5 gpc1345 (
      {stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209], stage1_9[210]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[39],stage2_11[60],stage2_10[65],stage2_9[80]}
   );
   gpc606_5 gpc1346 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[14],stage2_12[40],stage2_11[61],stage2_10[66]}
   );
   gpc606_5 gpc1347 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[15],stage2_12[41],stage2_11[62],stage2_10[67]}
   );
   gpc606_5 gpc1348 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[16],stage2_12[42],stage2_11[63],stage2_10[68]}
   );
   gpc606_5 gpc1349 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[17],stage2_12[43],stage2_11[64],stage2_10[69]}
   );
   gpc606_5 gpc1350 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[18],stage2_12[44],stage2_11[65],stage2_10[70]}
   );
   gpc606_5 gpc1351 (
      {stage1_10[186], stage1_10[187], stage1_10[188], stage1_10[189], stage1_10[190], stage1_10[191]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[19],stage2_12[45],stage2_11[66],stage2_10[71]}
   );
   gpc606_5 gpc1352 (
      {stage1_10[192], stage1_10[193], stage1_10[194], stage1_10[195], stage1_10[196], stage1_10[197]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[20],stage2_12[46],stage2_11[67],stage2_10[72]}
   );
   gpc606_5 gpc1353 (
      {stage1_10[198], stage1_10[199], stage1_10[200], stage1_10[201], stage1_10[202], stage1_10[203]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[21],stage2_12[47],stage2_11[68],stage2_10[73]}
   );
   gpc606_5 gpc1354 (
      {stage1_10[204], stage1_10[205], stage1_10[206], stage1_10[207], stage1_10[208], stage1_10[209]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[22],stage2_12[48],stage2_11[69],stage2_10[74]}
   );
   gpc606_5 gpc1355 (
      {stage1_10[210], stage1_10[211], stage1_10[212], stage1_10[213], stage1_10[214], stage1_10[215]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[23],stage2_12[49],stage2_11[70],stage2_10[75]}
   );
   gpc615_5 gpc1356 (
      {stage1_10[216], stage1_10[217], stage1_10[218], stage1_10[219], stage1_10[220]},
      {stage1_11[84]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[24],stage2_12[50],stage2_11[71],stage2_10[76]}
   );
   gpc615_5 gpc1357 (
      {stage1_10[221], stage1_10[222], stage1_10[223], stage1_10[224], stage1_10[225]},
      {stage1_11[85]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[25],stage2_12[51],stage2_11[72],stage2_10[77]}
   );
   gpc615_5 gpc1358 (
      {stage1_10[226], stage1_10[227], stage1_10[228], stage1_10[229], stage1_10[230]},
      {stage1_11[86]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[26],stage2_12[52],stage2_11[73],stage2_10[78]}
   );
   gpc615_5 gpc1359 (
      {stage1_10[231], stage1_10[232], stage1_10[233], stage1_10[234], stage1_10[235]},
      {stage1_11[87]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[27],stage2_12[53],stage2_11[74],stage2_10[79]}
   );
   gpc615_5 gpc1360 (
      {stage1_10[236], stage1_10[237], stage1_10[238], stage1_10[239], stage1_10[240]},
      {stage1_11[88]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[28],stage2_12[54],stage2_11[75],stage2_10[80]}
   );
   gpc615_5 gpc1361 (
      {stage1_10[241], stage1_10[242], stage1_10[243], stage1_10[244], stage1_10[245]},
      {stage1_11[89]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[29],stage2_12[55],stage2_11[76],stage2_10[81]}
   );
   gpc615_5 gpc1362 (
      {stage1_10[246], stage1_10[247], stage1_10[248], stage1_10[249], stage1_10[250]},
      {stage1_11[90]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage2_14[16],stage2_13[30],stage2_12[56],stage2_11[77],stage2_10[82]}
   );
   gpc615_5 gpc1363 (
      {stage1_10[251], stage1_10[252], stage1_10[253], stage1_10[254], stage1_10[255]},
      {stage1_11[91]},
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage2_14[17],stage2_13[31],stage2_12[57],stage2_11[78],stage2_10[83]}
   );
   gpc615_5 gpc1364 (
      {stage1_10[256], stage1_10[257], stage1_10[258], stage1_10[259], stage1_10[260]},
      {stage1_11[92]},
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage2_14[18],stage2_13[32],stage2_12[58],stage2_11[79],stage2_10[84]}
   );
   gpc615_5 gpc1365 (
      {stage1_10[261], stage1_10[262], stage1_10[263], stage1_10[264], stage1_10[265]},
      {stage1_11[93]},
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage2_14[19],stage2_13[33],stage2_12[59],stage2_11[80],stage2_10[85]}
   );
   gpc615_5 gpc1366 (
      {stage1_10[266], stage1_10[267], stage1_10[268], stage1_10[269], stage1_10[270]},
      {stage1_11[94]},
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage2_14[20],stage2_13[34],stage2_12[60],stage2_11[81],stage2_10[86]}
   );
   gpc615_5 gpc1367 (
      {stage1_10[271], stage1_10[272], stage1_10[273], stage1_10[274], stage1_10[275]},
      {stage1_11[95]},
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage2_14[21],stage2_13[35],stage2_12[61],stage2_11[82],stage2_10[87]}
   );
   gpc615_5 gpc1368 (
      {stage1_10[276], stage1_10[277], stage1_10[278], stage1_10[279], stage1_10[280]},
      {stage1_11[96]},
      {stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137]},
      {stage2_14[22],stage2_13[36],stage2_12[62],stage2_11[83],stage2_10[88]}
   );
   gpc606_5 gpc1369 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101], stage1_11[102]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[23],stage2_13[37],stage2_12[63],stage2_11[84]}
   );
   gpc606_5 gpc1370 (
      {stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[24],stage2_13[38],stage2_12[64],stage2_11[85]}
   );
   gpc615_5 gpc1371 (
      {stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage1_12[138]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[25],stage2_13[39],stage2_12[65],stage2_11[86]}
   );
   gpc615_5 gpc1372 (
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118]},
      {stage1_12[139]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[26],stage2_13[40],stage2_12[66],stage2_11[87]}
   );
   gpc615_5 gpc1373 (
      {stage1_11[119], stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123]},
      {stage1_12[140]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[27],stage2_13[41],stage2_12[67],stage2_11[88]}
   );
   gpc615_5 gpc1374 (
      {stage1_11[124], stage1_11[125], stage1_11[126], stage1_11[127], stage1_11[128]},
      {stage1_12[141]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[28],stage2_13[42],stage2_12[68],stage2_11[89]}
   );
   gpc615_5 gpc1375 (
      {stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132], stage1_11[133]},
      {stage1_12[142]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[29],stage2_13[43],stage2_12[69],stage2_11[90]}
   );
   gpc615_5 gpc1376 (
      {stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137], stage1_11[138]},
      {stage1_12[143]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[30],stage2_13[44],stage2_12[70],stage2_11[91]}
   );
   gpc615_5 gpc1377 (
      {stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143]},
      {stage1_12[144]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[31],stage2_13[45],stage2_12[71],stage2_11[92]}
   );
   gpc615_5 gpc1378 (
      {stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147], stage1_11[148]},
      {stage1_12[145]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[32],stage2_13[46],stage2_12[72],stage2_11[93]}
   );
   gpc615_5 gpc1379 (
      {stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152], stage1_11[153]},
      {stage1_12[146]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[33],stage2_13[47],stage2_12[73],stage2_11[94]}
   );
   gpc615_5 gpc1380 (
      {stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157], stage1_11[158]},
      {stage1_12[147]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[34],stage2_13[48],stage2_12[74],stage2_11[95]}
   );
   gpc615_5 gpc1381 (
      {stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162], stage1_11[163]},
      {stage1_12[148]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[35],stage2_13[49],stage2_12[75],stage2_11[96]}
   );
   gpc615_5 gpc1382 (
      {stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167], stage1_11[168]},
      {stage1_12[149]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[36],stage2_13[50],stage2_12[76],stage2_11[97]}
   );
   gpc615_5 gpc1383 (
      {stage1_11[169], stage1_11[170], stage1_11[171], stage1_11[172], stage1_11[173]},
      {stage1_12[150]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[37],stage2_13[51],stage2_12[77],stage2_11[98]}
   );
   gpc615_5 gpc1384 (
      {stage1_11[174], stage1_11[175], stage1_11[176], stage1_11[177], stage1_11[178]},
      {stage1_12[151]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[38],stage2_13[52],stage2_12[78],stage2_11[99]}
   );
   gpc615_5 gpc1385 (
      {stage1_11[179], stage1_11[180], stage1_11[181], stage1_11[182], stage1_11[183]},
      {stage1_12[152]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[39],stage2_13[53],stage2_12[79],stage2_11[100]}
   );
   gpc615_5 gpc1386 (
      {stage1_11[184], stage1_11[185], stage1_11[186], stage1_11[187], stage1_11[188]},
      {stage1_12[153]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[40],stage2_13[54],stage2_12[80],stage2_11[101]}
   );
   gpc615_5 gpc1387 (
      {stage1_11[189], stage1_11[190], stage1_11[191], stage1_11[192], stage1_11[193]},
      {stage1_12[154]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[41],stage2_13[55],stage2_12[81],stage2_11[102]}
   );
   gpc615_5 gpc1388 (
      {stage1_11[194], stage1_11[195], stage1_11[196], stage1_11[197], stage1_11[198]},
      {stage1_12[155]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[42],stage2_13[56],stage2_12[82],stage2_11[103]}
   );
   gpc615_5 gpc1389 (
      {stage1_11[199], stage1_11[200], stage1_11[201], stage1_11[202], stage1_11[203]},
      {stage1_12[156]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[43],stage2_13[57],stage2_12[83],stage2_11[104]}
   );
   gpc615_5 gpc1390 (
      {stage1_11[204], stage1_11[205], stage1_11[206], stage1_11[207], stage1_11[208]},
      {stage1_12[157]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[44],stage2_13[58],stage2_12[84],stage2_11[105]}
   );
   gpc615_5 gpc1391 (
      {stage1_11[209], stage1_11[210], stage1_11[211], stage1_11[212], stage1_11[213]},
      {stage1_12[158]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[45],stage2_13[59],stage2_12[85],stage2_11[106]}
   );
   gpc606_5 gpc1392 (
      {stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[23],stage2_14[46],stage2_13[60],stage2_12[86]}
   );
   gpc606_5 gpc1393 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[24],stage2_14[47],stage2_13[61],stage2_12[87]}
   );
   gpc606_5 gpc1394 (
      {stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174], stage1_12[175], stage1_12[176]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[25],stage2_14[48],stage2_13[62],stage2_12[88]}
   );
   gpc606_5 gpc1395 (
      {stage1_12[177], stage1_12[178], stage1_12[179], stage1_12[180], stage1_12[181], stage1_12[182]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[26],stage2_14[49],stage2_13[63],stage2_12[89]}
   );
   gpc606_5 gpc1396 (
      {stage1_12[183], stage1_12[184], stage1_12[185], stage1_12[186], stage1_12[187], stage1_12[188]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[27],stage2_14[50],stage2_13[64],stage2_12[90]}
   );
   gpc606_5 gpc1397 (
      {stage1_12[189], stage1_12[190], stage1_12[191], stage1_12[192], stage1_12[193], stage1_12[194]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[28],stage2_14[51],stage2_13[65],stage2_12[91]}
   );
   gpc606_5 gpc1398 (
      {stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198], stage1_12[199], stage1_12[200]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[29],stage2_14[52],stage2_13[66],stage2_12[92]}
   );
   gpc606_5 gpc1399 (
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[30],stage2_14[53],stage2_13[67]}
   );
   gpc606_5 gpc1400 (
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[8],stage2_15[31],stage2_14[54],stage2_13[68]}
   );
   gpc615_5 gpc1401 (
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154]},
      {stage1_14[42]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[9],stage2_15[32],stage2_14[55],stage2_13[69]}
   );
   gpc615_5 gpc1402 (
      {stage1_13[155], stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159]},
      {stage1_14[43]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[10],stage2_15[33],stage2_14[56],stage2_13[70]}
   );
   gpc615_5 gpc1403 (
      {stage1_13[160], stage1_13[161], stage1_13[162], stage1_13[163], stage1_13[164]},
      {stage1_14[44]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[11],stage2_15[34],stage2_14[57],stage2_13[71]}
   );
   gpc615_5 gpc1404 (
      {stage1_13[165], stage1_13[166], stage1_13[167], stage1_13[168], stage1_13[169]},
      {stage1_14[45]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[12],stage2_15[35],stage2_14[58],stage2_13[72]}
   );
   gpc615_5 gpc1405 (
      {stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173], stage1_13[174]},
      {stage1_14[46]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[13],stage2_15[36],stage2_14[59],stage2_13[73]}
   );
   gpc615_5 gpc1406 (
      {stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_14[47]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[14],stage2_15[37],stage2_14[60],stage2_13[74]}
   );
   gpc615_5 gpc1407 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184]},
      {stage1_14[48]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[15],stage2_15[38],stage2_14[61],stage2_13[75]}
   );
   gpc615_5 gpc1408 (
      {stage1_13[185], stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189]},
      {stage1_14[49]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[16],stage2_15[39],stage2_14[62],stage2_13[76]}
   );
   gpc615_5 gpc1409 (
      {stage1_13[190], stage1_13[191], stage1_13[192], stage1_13[193], stage1_13[194]},
      {stage1_14[50]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[17],stage2_15[40],stage2_14[63],stage2_13[77]}
   );
   gpc615_5 gpc1410 (
      {stage1_13[195], stage1_13[196], stage1_13[197], stage1_13[198], stage1_13[199]},
      {stage1_14[51]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[18],stage2_15[41],stage2_14[64],stage2_13[78]}
   );
   gpc615_5 gpc1411 (
      {stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203], stage1_13[204]},
      {stage1_14[52]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[19],stage2_15[42],stage2_14[65],stage2_13[79]}
   );
   gpc615_5 gpc1412 (
      {stage1_13[205], stage1_13[206], stage1_13[207], stage1_13[208], stage1_13[209]},
      {stage1_14[53]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[20],stage2_15[43],stage2_14[66],stage2_13[80]}
   );
   gpc615_5 gpc1413 (
      {stage1_13[210], stage1_13[211], stage1_13[212], stage1_13[213], stage1_13[214]},
      {stage1_14[54]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[21],stage2_15[44],stage2_14[67],stage2_13[81]}
   );
   gpc615_5 gpc1414 (
      {stage1_13[215], stage1_13[216], stage1_13[217], stage1_13[218], stage1_13[219]},
      {stage1_14[55]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[22],stage2_15[45],stage2_14[68],stage2_13[82]}
   );
   gpc615_5 gpc1415 (
      {stage1_13[220], stage1_13[221], stage1_13[222], stage1_13[223], stage1_13[224]},
      {stage1_14[56]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[23],stage2_15[46],stage2_14[69],stage2_13[83]}
   );
   gpc615_5 gpc1416 (
      {stage1_13[225], stage1_13[226], stage1_13[227], stage1_13[228], stage1_13[229]},
      {stage1_14[57]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[24],stage2_15[47],stage2_14[70],stage2_13[84]}
   );
   gpc615_5 gpc1417 (
      {stage1_13[230], stage1_13[231], stage1_13[232], stage1_13[233], stage1_13[234]},
      {stage1_14[58]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[25],stage2_15[48],stage2_14[71],stage2_13[85]}
   );
   gpc606_5 gpc1418 (
      {stage1_14[59], stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[19],stage2_16[26],stage2_15[49],stage2_14[72]}
   );
   gpc606_5 gpc1419 (
      {stage1_14[65], stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[20],stage2_16[27],stage2_15[50],stage2_14[73]}
   );
   gpc606_5 gpc1420 (
      {stage1_14[71], stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[21],stage2_16[28],stage2_15[51],stage2_14[74]}
   );
   gpc606_5 gpc1421 (
      {stage1_14[77], stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[22],stage2_16[29],stage2_15[52],stage2_14[75]}
   );
   gpc606_5 gpc1422 (
      {stage1_14[83], stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[23],stage2_16[30],stage2_15[53],stage2_14[76]}
   );
   gpc606_5 gpc1423 (
      {stage1_14[89], stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[24],stage2_16[31],stage2_15[54],stage2_14[77]}
   );
   gpc606_5 gpc1424 (
      {stage1_14[95], stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[25],stage2_16[32],stage2_15[55],stage2_14[78]}
   );
   gpc606_5 gpc1425 (
      {stage1_14[101], stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[26],stage2_16[33],stage2_15[56],stage2_14[79]}
   );
   gpc606_5 gpc1426 (
      {stage1_14[107], stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[27],stage2_16[34],stage2_15[57],stage2_14[80]}
   );
   gpc606_5 gpc1427 (
      {stage1_14[113], stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[28],stage2_16[35],stage2_15[58],stage2_14[81]}
   );
   gpc615_5 gpc1428 (
      {stage1_14[119], stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123]},
      {stage1_15[114]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[29],stage2_16[36],stage2_15[59],stage2_14[82]}
   );
   gpc615_5 gpc1429 (
      {stage1_14[124], stage1_14[125], stage1_14[126], stage1_14[127], stage1_14[128]},
      {stage1_15[115]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[30],stage2_16[37],stage2_15[60],stage2_14[83]}
   );
   gpc615_5 gpc1430 (
      {stage1_14[129], stage1_14[130], stage1_14[131], stage1_14[132], stage1_14[133]},
      {stage1_15[116]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[31],stage2_16[38],stage2_15[61],stage2_14[84]}
   );
   gpc615_5 gpc1431 (
      {stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138]},
      {stage1_15[117]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[32],stage2_16[39],stage2_15[62],stage2_14[85]}
   );
   gpc615_5 gpc1432 (
      {stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage1_15[118]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[33],stage2_16[40],stage2_15[63],stage2_14[86]}
   );
   gpc615_5 gpc1433 (
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148]},
      {stage1_15[119]},
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage2_18[15],stage2_17[34],stage2_16[41],stage2_15[64],stage2_14[87]}
   );
   gpc615_5 gpc1434 (
      {stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153]},
      {stage1_15[120]},
      {stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101]},
      {stage2_18[16],stage2_17[35],stage2_16[42],stage2_15[65],stage2_14[88]}
   );
   gpc615_5 gpc1435 (
      {stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157], stage1_14[158]},
      {stage1_15[121]},
      {stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107]},
      {stage2_18[17],stage2_17[36],stage2_16[43],stage2_15[66],stage2_14[89]}
   );
   gpc615_5 gpc1436 (
      {stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163]},
      {stage1_15[122]},
      {stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113]},
      {stage2_18[18],stage2_17[37],stage2_16[44],stage2_15[67],stage2_14[90]}
   );
   gpc615_5 gpc1437 (
      {stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168]},
      {stage1_15[123]},
      {stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119]},
      {stage2_18[19],stage2_17[38],stage2_16[45],stage2_15[68],stage2_14[91]}
   );
   gpc615_5 gpc1438 (
      {stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage1_15[124]},
      {stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125]},
      {stage2_18[20],stage2_17[39],stage2_16[46],stage2_15[69],stage2_14[92]}
   );
   gpc606_5 gpc1439 (
      {stage1_15[125], stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[21],stage2_17[40],stage2_16[47],stage2_15[70]}
   );
   gpc606_5 gpc1440 (
      {stage1_15[131], stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[22],stage2_17[41],stage2_16[48],stage2_15[71]}
   );
   gpc606_5 gpc1441 (
      {stage1_15[137], stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[23],stage2_17[42],stage2_16[49],stage2_15[72]}
   );
   gpc606_5 gpc1442 (
      {stage1_15[143], stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[24],stage2_17[43],stage2_16[50],stage2_15[73]}
   );
   gpc606_5 gpc1443 (
      {stage1_15[149], stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[25],stage2_17[44],stage2_16[51],stage2_15[74]}
   );
   gpc1_1 gpc1444 (
      {stage1_0[138]},
      {stage2_0[28]}
   );
   gpc1_1 gpc1445 (
      {stage1_0[139]},
      {stage2_0[29]}
   );
   gpc1_1 gpc1446 (
      {stage1_0[140]},
      {stage2_0[30]}
   );
   gpc1_1 gpc1447 (
      {stage1_0[141]},
      {stage2_0[31]}
   );
   gpc1_1 gpc1448 (
      {stage1_0[142]},
      {stage2_0[32]}
   );
   gpc1_1 gpc1449 (
      {stage1_0[143]},
      {stage2_0[33]}
   );
   gpc1_1 gpc1450 (
      {stage1_0[144]},
      {stage2_0[34]}
   );
   gpc1_1 gpc1451 (
      {stage1_0[145]},
      {stage2_0[35]}
   );
   gpc1_1 gpc1452 (
      {stage1_0[146]},
      {stage2_0[36]}
   );
   gpc1_1 gpc1453 (
      {stage1_0[147]},
      {stage2_0[37]}
   );
   gpc1_1 gpc1454 (
      {stage1_1[108]},
      {stage2_1[36]}
   );
   gpc1_1 gpc1455 (
      {stage1_1[109]},
      {stage2_1[37]}
   );
   gpc1_1 gpc1456 (
      {stage1_1[110]},
      {stage2_1[38]}
   );
   gpc1_1 gpc1457 (
      {stage1_1[111]},
      {stage2_1[39]}
   );
   gpc1_1 gpc1458 (
      {stage1_1[112]},
      {stage2_1[40]}
   );
   gpc1_1 gpc1459 (
      {stage1_1[113]},
      {stage2_1[41]}
   );
   gpc1_1 gpc1460 (
      {stage1_1[114]},
      {stage2_1[42]}
   );
   gpc1_1 gpc1461 (
      {stage1_1[115]},
      {stage2_1[43]}
   );
   gpc1_1 gpc1462 (
      {stage1_1[116]},
      {stage2_1[44]}
   );
   gpc1_1 gpc1463 (
      {stage1_1[117]},
      {stage2_1[45]}
   );
   gpc1_1 gpc1464 (
      {stage1_1[118]},
      {stage2_1[46]}
   );
   gpc1_1 gpc1465 (
      {stage1_1[119]},
      {stage2_1[47]}
   );
   gpc1_1 gpc1466 (
      {stage1_1[120]},
      {stage2_1[48]}
   );
   gpc1_1 gpc1467 (
      {stage1_1[121]},
      {stage2_1[49]}
   );
   gpc1_1 gpc1468 (
      {stage1_1[122]},
      {stage2_1[50]}
   );
   gpc1_1 gpc1469 (
      {stage1_1[123]},
      {stage2_1[51]}
   );
   gpc1_1 gpc1470 (
      {stage1_1[124]},
      {stage2_1[52]}
   );
   gpc1_1 gpc1471 (
      {stage1_1[125]},
      {stage2_1[53]}
   );
   gpc1_1 gpc1472 (
      {stage1_1[126]},
      {stage2_1[54]}
   );
   gpc1_1 gpc1473 (
      {stage1_1[127]},
      {stage2_1[55]}
   );
   gpc1_1 gpc1474 (
      {stage1_1[128]},
      {stage2_1[56]}
   );
   gpc1_1 gpc1475 (
      {stage1_1[129]},
      {stage2_1[57]}
   );
   gpc1_1 gpc1476 (
      {stage1_1[130]},
      {stage2_1[58]}
   );
   gpc1_1 gpc1477 (
      {stage1_1[131]},
      {stage2_1[59]}
   );
   gpc1_1 gpc1478 (
      {stage1_1[132]},
      {stage2_1[60]}
   );
   gpc1_1 gpc1479 (
      {stage1_1[133]},
      {stage2_1[61]}
   );
   gpc1_1 gpc1480 (
      {stage1_1[134]},
      {stage2_1[62]}
   );
   gpc1_1 gpc1481 (
      {stage1_2[158]},
      {stage2_2[44]}
   );
   gpc1_1 gpc1482 (
      {stage1_2[159]},
      {stage2_2[45]}
   );
   gpc1_1 gpc1483 (
      {stage1_2[160]},
      {stage2_2[46]}
   );
   gpc1_1 gpc1484 (
      {stage1_2[161]},
      {stage2_2[47]}
   );
   gpc1_1 gpc1485 (
      {stage1_2[162]},
      {stage2_2[48]}
   );
   gpc1_1 gpc1486 (
      {stage1_2[163]},
      {stage2_2[49]}
   );
   gpc1_1 gpc1487 (
      {stage1_2[164]},
      {stage2_2[50]}
   );
   gpc1_1 gpc1488 (
      {stage1_2[165]},
      {stage2_2[51]}
   );
   gpc1_1 gpc1489 (
      {stage1_2[166]},
      {stage2_2[52]}
   );
   gpc1_1 gpc1490 (
      {stage1_2[167]},
      {stage2_2[53]}
   );
   gpc1_1 gpc1491 (
      {stage1_3[236]},
      {stage2_3[78]}
   );
   gpc1_1 gpc1492 (
      {stage1_3[237]},
      {stage2_3[79]}
   );
   gpc1_1 gpc1493 (
      {stage1_3[238]},
      {stage2_3[80]}
   );
   gpc1_1 gpc1494 (
      {stage1_3[239]},
      {stage2_3[81]}
   );
   gpc1_1 gpc1495 (
      {stage1_3[240]},
      {stage2_3[82]}
   );
   gpc1_1 gpc1496 (
      {stage1_3[241]},
      {stage2_3[83]}
   );
   gpc1_1 gpc1497 (
      {stage1_3[242]},
      {stage2_3[84]}
   );
   gpc1_1 gpc1498 (
      {stage1_3[243]},
      {stage2_3[85]}
   );
   gpc1_1 gpc1499 (
      {stage1_4[222]},
      {stage2_4[106]}
   );
   gpc1_1 gpc1500 (
      {stage1_5[322]},
      {stage2_5[93]}
   );
   gpc1_1 gpc1501 (
      {stage1_5[323]},
      {stage2_5[94]}
   );
   gpc1_1 gpc1502 (
      {stage1_5[324]},
      {stage2_5[95]}
   );
   gpc1_1 gpc1503 (
      {stage1_5[325]},
      {stage2_5[96]}
   );
   gpc1_1 gpc1504 (
      {stage1_5[326]},
      {stage2_5[97]}
   );
   gpc1_1 gpc1505 (
      {stage1_5[327]},
      {stage2_5[98]}
   );
   gpc1_1 gpc1506 (
      {stage1_5[328]},
      {stage2_5[99]}
   );
   gpc1_1 gpc1507 (
      {stage1_5[329]},
      {stage2_5[100]}
   );
   gpc1_1 gpc1508 (
      {stage1_5[330]},
      {stage2_5[101]}
   );
   gpc1_1 gpc1509 (
      {stage1_5[331]},
      {stage2_5[102]}
   );
   gpc1_1 gpc1510 (
      {stage1_5[332]},
      {stage2_5[103]}
   );
   gpc1_1 gpc1511 (
      {stage1_5[333]},
      {stage2_5[104]}
   );
   gpc1_1 gpc1512 (
      {stage1_5[334]},
      {stage2_5[105]}
   );
   gpc1_1 gpc1513 (
      {stage1_5[335]},
      {stage2_5[106]}
   );
   gpc1_1 gpc1514 (
      {stage1_5[336]},
      {stage2_5[107]}
   );
   gpc1_1 gpc1515 (
      {stage1_8[185]},
      {stage2_8[95]}
   );
   gpc1_1 gpc1516 (
      {stage1_8[186]},
      {stage2_8[96]}
   );
   gpc1_1 gpc1517 (
      {stage1_8[187]},
      {stage2_8[97]}
   );
   gpc1_1 gpc1518 (
      {stage1_8[188]},
      {stage2_8[98]}
   );
   gpc1_1 gpc1519 (
      {stage1_8[189]},
      {stage2_8[99]}
   );
   gpc1_1 gpc1520 (
      {stage1_8[190]},
      {stage2_8[100]}
   );
   gpc1_1 gpc1521 (
      {stage1_8[191]},
      {stage2_8[101]}
   );
   gpc1_1 gpc1522 (
      {stage1_8[192]},
      {stage2_8[102]}
   );
   gpc1_1 gpc1523 (
      {stage1_8[193]},
      {stage2_8[103]}
   );
   gpc1_1 gpc1524 (
      {stage1_8[194]},
      {stage2_8[104]}
   );
   gpc1_1 gpc1525 (
      {stage1_8[195]},
      {stage2_8[105]}
   );
   gpc1_1 gpc1526 (
      {stage1_10[281]},
      {stage2_10[89]}
   );
   gpc1_1 gpc1527 (
      {stage1_12[201]},
      {stage2_12[93]}
   );
   gpc1_1 gpc1528 (
      {stage1_14[174]},
      {stage2_14[93]}
   );
   gpc1_1 gpc1529 (
      {stage1_14[175]},
      {stage2_14[94]}
   );
   gpc1_1 gpc1530 (
      {stage1_14[176]},
      {stage2_14[95]}
   );
   gpc1_1 gpc1531 (
      {stage1_14[177]},
      {stage2_14[96]}
   );
   gpc1_1 gpc1532 (
      {stage1_14[178]},
      {stage2_14[97]}
   );
   gpc1_1 gpc1533 (
      {stage1_14[179]},
      {stage2_14[98]}
   );
   gpc1_1 gpc1534 (
      {stage1_14[180]},
      {stage2_14[99]}
   );
   gpc1_1 gpc1535 (
      {stage1_14[181]},
      {stage2_14[100]}
   );
   gpc1_1 gpc1536 (
      {stage1_14[182]},
      {stage2_14[101]}
   );
   gpc1_1 gpc1537 (
      {stage1_16[126]},
      {stage2_16[52]}
   );
   gpc1_1 gpc1538 (
      {stage1_16[127]},
      {stage2_16[53]}
   );
   gpc1_1 gpc1539 (
      {stage1_16[128]},
      {stage2_16[54]}
   );
   gpc1_1 gpc1540 (
      {stage1_16[129]},
      {stage2_16[55]}
   );
   gpc1_1 gpc1541 (
      {stage1_16[130]},
      {stage2_16[56]}
   );
   gpc1_1 gpc1542 (
      {stage1_16[131]},
      {stage2_16[57]}
   );
   gpc1_1 gpc1543 (
      {stage1_16[132]},
      {stage2_16[58]}
   );
   gpc1_1 gpc1544 (
      {stage1_16[133]},
      {stage2_16[59]}
   );
   gpc1_1 gpc1545 (
      {stage1_16[134]},
      {stage2_16[60]}
   );
   gpc1_1 gpc1546 (
      {stage1_16[135]},
      {stage2_16[61]}
   );
   gpc1_1 gpc1547 (
      {stage1_16[136]},
      {stage2_16[62]}
   );
   gpc1_1 gpc1548 (
      {stage1_16[137]},
      {stage2_16[63]}
   );
   gpc1_1 gpc1549 (
      {stage1_16[138]},
      {stage2_16[64]}
   );
   gpc1_1 gpc1550 (
      {stage1_16[139]},
      {stage2_16[65]}
   );
   gpc1_1 gpc1551 (
      {stage1_16[140]},
      {stage2_16[66]}
   );
   gpc1_1 gpc1552 (
      {stage1_16[141]},
      {stage2_16[67]}
   );
   gpc1_1 gpc1553 (
      {stage1_16[142]},
      {stage2_16[68]}
   );
   gpc1_1 gpc1554 (
      {stage1_16[143]},
      {stage2_16[69]}
   );
   gpc1_1 gpc1555 (
      {stage1_16[144]},
      {stage2_16[70]}
   );
   gpc1_1 gpc1556 (
      {stage1_16[145]},
      {stage2_16[71]}
   );
   gpc1_1 gpc1557 (
      {stage1_16[146]},
      {stage2_16[72]}
   );
   gpc1_1 gpc1558 (
      {stage1_16[147]},
      {stage2_16[73]}
   );
   gpc1_1 gpc1559 (
      {stage1_16[148]},
      {stage2_16[74]}
   );
   gpc1_1 gpc1560 (
      {stage1_16[149]},
      {stage2_16[75]}
   );
   gpc1_1 gpc1561 (
      {stage1_16[150]},
      {stage2_16[76]}
   );
   gpc1_1 gpc1562 (
      {stage1_17[30]},
      {stage2_17[45]}
   );
   gpc1_1 gpc1563 (
      {stage1_17[31]},
      {stage2_17[46]}
   );
   gpc1_1 gpc1564 (
      {stage1_17[32]},
      {stage2_17[47]}
   );
   gpc1_1 gpc1565 (
      {stage1_17[33]},
      {stage2_17[48]}
   );
   gpc1_1 gpc1566 (
      {stage1_17[34]},
      {stage2_17[49]}
   );
   gpc1_1 gpc1567 (
      {stage1_17[35]},
      {stage2_17[50]}
   );
   gpc1_1 gpc1568 (
      {stage1_17[36]},
      {stage2_17[51]}
   );
   gpc1_1 gpc1569 (
      {stage1_17[37]},
      {stage2_17[52]}
   );
   gpc1_1 gpc1570 (
      {stage1_17[38]},
      {stage2_17[53]}
   );
   gpc1_1 gpc1571 (
      {stage1_17[39]},
      {stage2_17[54]}
   );
   gpc1_1 gpc1572 (
      {stage1_17[40]},
      {stage2_17[55]}
   );
   gpc1_1 gpc1573 (
      {stage1_17[41]},
      {stage2_17[56]}
   );
   gpc1_1 gpc1574 (
      {stage1_17[42]},
      {stage2_17[57]}
   );
   gpc1_1 gpc1575 (
      {stage1_17[43]},
      {stage2_17[58]}
   );
   gpc1_1 gpc1576 (
      {stage1_17[44]},
      {stage2_17[59]}
   );
   gpc1_1 gpc1577 (
      {stage1_17[45]},
      {stage2_17[60]}
   );
   gpc1_1 gpc1578 (
      {stage1_17[46]},
      {stage2_17[61]}
   );
   gpc1_1 gpc1579 (
      {stage1_17[47]},
      {stage2_17[62]}
   );
   gpc1_1 gpc1580 (
      {stage1_17[48]},
      {stage2_17[63]}
   );
   gpc1_1 gpc1581 (
      {stage1_17[49]},
      {stage2_17[64]}
   );
   gpc1_1 gpc1582 (
      {stage1_17[50]},
      {stage2_17[65]}
   );
   gpc1_1 gpc1583 (
      {stage1_17[51]},
      {stage2_17[66]}
   );
   gpc1_1 gpc1584 (
      {stage1_17[52]},
      {stage2_17[67]}
   );
   gpc1_1 gpc1585 (
      {stage1_17[53]},
      {stage2_17[68]}
   );
   gpc1_1 gpc1586 (
      {stage1_17[54]},
      {stage2_17[69]}
   );
   gpc1_1 gpc1587 (
      {stage1_17[55]},
      {stage2_17[70]}
   );
   gpc1_1 gpc1588 (
      {stage1_17[56]},
      {stage2_17[71]}
   );
   gpc1_1 gpc1589 (
      {stage1_17[57]},
      {stage2_17[72]}
   );
   gpc1_1 gpc1590 (
      {stage1_17[58]},
      {stage2_17[73]}
   );
   gpc1_1 gpc1591 (
      {stage1_17[59]},
      {stage2_17[74]}
   );
   gpc1_1 gpc1592 (
      {stage1_17[60]},
      {stage2_17[75]}
   );
   gpc1_1 gpc1593 (
      {stage1_17[61]},
      {stage2_17[76]}
   );
   gpc1_1 gpc1594 (
      {stage1_17[62]},
      {stage2_17[77]}
   );
   gpc1_1 gpc1595 (
      {stage1_17[63]},
      {stage2_17[78]}
   );
   gpc1_1 gpc1596 (
      {stage1_17[64]},
      {stage2_17[79]}
   );
   gpc1_1 gpc1597 (
      {stage1_17[65]},
      {stage2_17[80]}
   );
   gpc1_1 gpc1598 (
      {stage1_17[66]},
      {stage2_17[81]}
   );
   gpc1_1 gpc1599 (
      {stage1_17[67]},
      {stage2_17[82]}
   );
   gpc1_1 gpc1600 (
      {stage1_17[68]},
      {stage2_17[83]}
   );
   gpc1_1 gpc1601 (
      {stage1_17[69]},
      {stage2_17[84]}
   );
   gpc1_1 gpc1602 (
      {stage1_17[70]},
      {stage2_17[85]}
   );
   gpc1_1 gpc1603 (
      {stage1_17[71]},
      {stage2_17[86]}
   );
   gpc1_1 gpc1604 (
      {stage1_17[72]},
      {stage2_17[87]}
   );
   gpc1_1 gpc1605 (
      {stage1_17[73]},
      {stage2_17[88]}
   );
   gpc1_1 gpc1606 (
      {stage1_17[74]},
      {stage2_17[89]}
   );
   gpc1_1 gpc1607 (
      {stage1_17[75]},
      {stage2_17[90]}
   );
   gpc1_1 gpc1608 (
      {stage1_17[76]},
      {stage2_17[91]}
   );
   gpc1_1 gpc1609 (
      {stage1_17[77]},
      {stage2_17[92]}
   );
   gpc1_1 gpc1610 (
      {stage1_17[78]},
      {stage2_17[93]}
   );
   gpc1_1 gpc1611 (
      {stage1_17[79]},
      {stage2_17[94]}
   );
   gpc1_1 gpc1612 (
      {stage1_17[80]},
      {stage2_17[95]}
   );
   gpc1163_5 gpc1613 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc1614 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc1615 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[2]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1163_5 gpc1616 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[3]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1617 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc1618 (
      {stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23]},
      {stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc1619 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc1620 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc1621 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc1622 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27]},
      {stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc1623 (
      {stage2_1[48], stage2_1[49], stage2_1[50], stage2_1[51], stage2_1[52], stage2_1[53]},
      {stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10]}
   );
   gpc606_5 gpc1624 (
      {stage2_1[54], stage2_1[55], stage2_1[56], stage2_1[57], stage2_1[58], stage2_1[59]},
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc1625 (
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc606_5 gpc1626 (
      {stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc606_5 gpc1627 (
      {stage2_2[28], stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc1628 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[40]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc1629 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[41]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc615_5 gpc1630 (
      {stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage2_3[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[17],stage3_3[17],stage3_2[17]}
   );
   gpc615_5 gpc1631 (
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53]},
      {stage2_3[43]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc615_5 gpc1632 (
      {stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage2_4[42]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc1633 (
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53]},
      {stage2_4[43]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc1634 (
      {stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58]},
      {stage2_4[44]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc1635 (
      {stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63]},
      {stage2_4[45]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc1636 (
      {stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_4[46]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc606_5 gpc1637 (
      {stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51], stage2_4[52]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[24]}
   );
   gpc606_5 gpc1638 (
      {stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[25]}
   );
   gpc606_5 gpc1639 (
      {stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[26]}
   );
   gpc606_5 gpc1640 (
      {stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[27]}
   );
   gpc606_5 gpc1641 (
      {stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[28]}
   );
   gpc606_5 gpc1642 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[29]}
   );
   gpc606_5 gpc1643 (
      {stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[30]}
   );
   gpc606_5 gpc1644 (
      {stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[31]}
   );
   gpc606_5 gpc1645 (
      {stage2_4[95], stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[32]}
   );
   gpc606_5 gpc1646 (
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[9],stage3_7[14],stage3_6[21],stage3_5[27]}
   );
   gpc606_5 gpc1647 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[10],stage3_7[15],stage3_6[22],stage3_5[28]}
   );
   gpc606_5 gpc1648 (
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[11],stage3_7[16],stage3_6[23],stage3_5[29]}
   );
   gpc606_5 gpc1649 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[12],stage3_7[17],stage3_6[24],stage3_5[30]}
   );
   gpc606_5 gpc1650 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[13],stage3_7[18],stage3_6[25],stage3_5[31]}
   );
   gpc606_5 gpc1651 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[14],stage3_7[19],stage3_6[26],stage3_5[32]}
   );
   gpc606_5 gpc1652 (
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage2_7[36], stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage3_9[6],stage3_8[15],stage3_7[20],stage3_6[27],stage3_5[33]}
   );
   gpc606_5 gpc1653 (
      {stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77]},
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage3_9[7],stage3_8[16],stage3_7[21],stage3_6[28],stage3_5[34]}
   );
   gpc606_5 gpc1654 (
      {stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51], stage2_7[52], stage2_7[53]},
      {stage3_9[8],stage3_8[17],stage3_7[22],stage3_6[29],stage3_5[35]}
   );
   gpc606_5 gpc1655 (
      {stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87], stage2_5[88], stage2_5[89]},
      {stage2_7[54], stage2_7[55], stage2_7[56], stage2_7[57], stage2_7[58], stage2_7[59]},
      {stage3_9[9],stage3_8[18],stage3_7[23],stage3_6[30],stage3_5[36]}
   );
   gpc606_5 gpc1656 (
      {stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93], stage2_5[94], stage2_5[95]},
      {stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65]},
      {stage3_9[10],stage3_8[19],stage3_7[24],stage3_6[31],stage3_5[37]}
   );
   gpc606_5 gpc1657 (
      {stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99], stage2_5[100], stage2_5[101]},
      {stage2_7[66], stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage3_9[11],stage3_8[20],stage3_7[25],stage3_6[32],stage3_5[38]}
   );
   gpc606_5 gpc1658 (
      {stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105], stage2_5[106], stage2_5[107]},
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76], stage2_7[77]},
      {stage3_9[12],stage3_8[21],stage3_7[26],stage3_6[33],stage3_5[39]}
   );
   gpc615_5 gpc1659 (
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58]},
      {stage2_7[78]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[13],stage3_8[22],stage3_7[27],stage3_6[34]}
   );
   gpc615_5 gpc1660 (
      {stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63]},
      {stage2_7[79]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[14],stage3_8[23],stage3_7[28],stage3_6[35]}
   );
   gpc615_5 gpc1661 (
      {stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67], stage2_6[68]},
      {stage2_7[80]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[15],stage3_8[24],stage3_7[29],stage3_6[36]}
   );
   gpc615_5 gpc1662 (
      {stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_7[81]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[16],stage3_8[25],stage3_7[30],stage3_6[37]}
   );
   gpc615_5 gpc1663 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78]},
      {stage2_7[82]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[17],stage3_8[26],stage3_7[31],stage3_6[38]}
   );
   gpc615_5 gpc1664 (
      {stage2_7[83], stage2_7[84], stage2_7[85], stage2_7[86], stage2_7[87]},
      {stage2_8[30]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[5],stage3_9[18],stage3_8[27],stage3_7[32]}
   );
   gpc615_5 gpc1665 (
      {stage2_7[88], stage2_7[89], stage2_7[90], stage2_7[91], stage2_7[92]},
      {stage2_8[31]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[6],stage3_9[19],stage3_8[28],stage3_7[33]}
   );
   gpc615_5 gpc1666 (
      {stage2_7[93], stage2_7[94], stage2_7[95], stage2_7[96], stage2_7[97]},
      {stage2_8[32]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[7],stage3_9[20],stage3_8[29],stage3_7[34]}
   );
   gpc615_5 gpc1667 (
      {stage2_7[98], stage2_7[99], stage2_7[100], stage2_7[101], stage2_7[102]},
      {stage2_8[33]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[8],stage3_9[21],stage3_8[30],stage3_7[35]}
   );
   gpc606_5 gpc1668 (
      {stage2_8[34], stage2_8[35], stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[9],stage3_9[22],stage3_8[31]}
   );
   gpc606_5 gpc1669 (
      {stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[10],stage3_9[23],stage3_8[32]}
   );
   gpc606_5 gpc1670 (
      {stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[11],stage3_9[24],stage3_8[33]}
   );
   gpc606_5 gpc1671 (
      {stage2_8[52], stage2_8[53], stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[12],stage3_9[25],stage3_8[34]}
   );
   gpc606_5 gpc1672 (
      {stage2_8[58], stage2_8[59], stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[13],stage3_9[26],stage3_8[35]}
   );
   gpc606_5 gpc1673 (
      {stage2_8[64], stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[9],stage3_10[14],stage3_9[27],stage3_8[36]}
   );
   gpc606_5 gpc1674 (
      {stage2_8[70], stage2_8[71], stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[10],stage3_10[15],stage3_9[28],stage3_8[37]}
   );
   gpc606_5 gpc1675 (
      {stage2_8[76], stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[11],stage3_10[16],stage3_9[29],stage3_8[38]}
   );
   gpc606_5 gpc1676 (
      {stage2_8[82], stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[8],stage3_11[12],stage3_10[17],stage3_9[30],stage3_8[39]}
   );
   gpc606_5 gpc1677 (
      {stage2_8[88], stage2_8[89], stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[9],stage3_11[13],stage3_10[18],stage3_9[31],stage3_8[40]}
   );
   gpc606_5 gpc1678 (
      {stage2_8[94], stage2_8[95], stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[10],stage3_11[14],stage3_10[19],stage3_9[32],stage3_8[41]}
   );
   gpc207_4 gpc1679 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30]},
      {stage2_11[0], stage2_11[1]},
      {stage3_12[11],stage3_11[15],stage3_10[20],stage3_9[33]}
   );
   gpc207_4 gpc1680 (
      {stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35], stage2_9[36], stage2_9[37]},
      {stage2_11[2], stage2_11[3]},
      {stage3_12[12],stage3_11[16],stage3_10[21],stage3_9[34]}
   );
   gpc606_5 gpc1681 (
      {stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41], stage2_9[42], stage2_9[43]},
      {stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage3_13[0],stage3_12[13],stage3_11[17],stage3_10[22],stage3_9[35]}
   );
   gpc606_5 gpc1682 (
      {stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48], stage2_9[49]},
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15]},
      {stage3_13[1],stage3_12[14],stage3_11[18],stage3_10[23],stage3_9[36]}
   );
   gpc606_5 gpc1683 (
      {stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54], stage2_9[55]},
      {stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage3_13[2],stage3_12[15],stage3_11[19],stage3_10[24],stage3_9[37]}
   );
   gpc606_5 gpc1684 (
      {stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60], stage2_9[61]},
      {stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage3_13[3],stage3_12[16],stage3_11[20],stage3_10[25],stage3_9[38]}
   );
   gpc606_5 gpc1685 (
      {stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65], stage2_9[66], stage2_9[67]},
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage3_13[4],stage3_12[17],stage3_11[21],stage3_10[26],stage3_9[39]}
   );
   gpc606_5 gpc1686 (
      {stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71], stage2_9[72], stage2_9[73]},
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage3_13[5],stage3_12[18],stage3_11[22],stage3_10[27],stage3_9[40]}
   );
   gpc606_5 gpc1687 (
      {stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79]},
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45]},
      {stage3_13[6],stage3_12[19],stage3_11[23],stage3_10[28],stage3_9[41]}
   );
   gpc606_5 gpc1688 (
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[7],stage3_12[20],stage3_11[24],stage3_10[29]}
   );
   gpc615_5 gpc1689 (
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76]},
      {stage2_11[46]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[8],stage3_12[21],stage3_11[25],stage3_10[30]}
   );
   gpc615_5 gpc1690 (
      {stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51]},
      {stage2_12[12]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[9],stage3_12[22],stage3_11[26]}
   );
   gpc615_5 gpc1691 (
      {stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56]},
      {stage2_12[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[10],stage3_12[23],stage3_11[27]}
   );
   gpc615_5 gpc1692 (
      {stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61]},
      {stage2_12[14]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[4],stage3_13[11],stage3_12[24],stage3_11[28]}
   );
   gpc615_5 gpc1693 (
      {stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66]},
      {stage2_12[15]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[5],stage3_13[12],stage3_12[25],stage3_11[29]}
   );
   gpc615_5 gpc1694 (
      {stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage2_12[16]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[6],stage3_13[13],stage3_12[26],stage3_11[30]}
   );
   gpc615_5 gpc1695 (
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76]},
      {stage2_12[17]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[7],stage3_13[14],stage3_12[27],stage3_11[31]}
   );
   gpc615_5 gpc1696 (
      {stage2_11[77], stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81]},
      {stage2_12[18]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[8],stage3_13[15],stage3_12[28],stage3_11[32]}
   );
   gpc615_5 gpc1697 (
      {stage2_11[82], stage2_11[83], stage2_11[84], stage2_11[85], stage2_11[86]},
      {stage2_12[19]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[9],stage3_13[16],stage3_12[29],stage3_11[33]}
   );
   gpc615_5 gpc1698 (
      {stage2_11[87], stage2_11[88], stage2_11[89], stage2_11[90], stage2_11[91]},
      {stage2_12[20]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[10],stage3_13[17],stage3_12[30],stage3_11[34]}
   );
   gpc615_5 gpc1699 (
      {stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96]},
      {stage2_12[21]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[11],stage3_13[18],stage3_12[31],stage3_11[35]}
   );
   gpc615_5 gpc1700 (
      {stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101]},
      {stage2_12[22]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[12],stage3_13[19],stage3_12[32],stage3_11[36]}
   );
   gpc615_5 gpc1701 (
      {stage2_11[102], stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106]},
      {stage2_12[23]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[13],stage3_13[20],stage3_12[33],stage3_11[37]}
   );
   gpc606_5 gpc1702 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[12],stage3_14[14],stage3_13[21],stage3_12[34]}
   );
   gpc606_5 gpc1703 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[13],stage3_14[15],stage3_13[22],stage3_12[35]}
   );
   gpc606_5 gpc1704 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[14],stage3_14[16],stage3_13[23],stage3_12[36]}
   );
   gpc606_5 gpc1705 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[15],stage3_14[17],stage3_13[24],stage3_12[37]}
   );
   gpc606_5 gpc1706 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[16],stage3_14[18],stage3_13[25],stage3_12[38]}
   );
   gpc615_5 gpc1707 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58]},
      {stage2_13[72]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[17],stage3_14[19],stage3_13[26],stage3_12[39]}
   );
   gpc615_5 gpc1708 (
      {stage2_12[59], stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63]},
      {stage2_13[73]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[18],stage3_14[20],stage3_13[27],stage3_12[40]}
   );
   gpc615_5 gpc1709 (
      {stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67], stage2_12[68]},
      {stage2_13[74]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[19],stage3_14[21],stage3_13[28],stage3_12[41]}
   );
   gpc615_5 gpc1710 (
      {stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_13[75]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[20],stage3_14[22],stage3_13[29],stage3_12[42]}
   );
   gpc615_5 gpc1711 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78]},
      {stage2_13[76]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[21],stage3_14[23],stage3_13[30],stage3_12[43]}
   );
   gpc615_5 gpc1712 (
      {stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83]},
      {stage2_13[77]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[22],stage3_14[24],stage3_13[31],stage3_12[44]}
   );
   gpc615_5 gpc1713 (
      {stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88]},
      {stage2_13[78]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[23],stage3_14[25],stage3_13[32],stage3_12[45]}
   );
   gpc615_5 gpc1714 (
      {stage2_12[89], stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93]},
      {stage2_13[79]},
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage3_16[12],stage3_15[24],stage3_14[26],stage3_13[33],stage3_12[46]}
   );
   gpc615_5 gpc1715 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[13],stage3_15[25],stage3_14[27]}
   );
   gpc615_5 gpc1716 (
      {stage2_14[83], stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[14],stage3_15[26],stage3_14[28]}
   );
   gpc615_5 gpc1717 (
      {stage2_14[88], stage2_14[89], stage2_14[90], stage2_14[91], stage2_14[92]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[15],stage3_15[27],stage3_14[29]}
   );
   gpc615_5 gpc1718 (
      {stage2_14[93], stage2_14[94], stage2_14[95], stage2_14[96], stage2_14[97]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[16],stage3_15[28],stage3_14[30]}
   );
   gpc615_5 gpc1719 (
      {stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101], 1'b0},
      {stage2_15[4]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[4],stage3_16[17],stage3_15[29],stage3_14[31]}
   );
   gpc615_5 gpc1720 (
      {stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9]},
      {stage2_16[30]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[5],stage3_17[5],stage3_16[18],stage3_15[30]}
   );
   gpc615_5 gpc1721 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[31]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[6],stage3_17[6],stage3_16[19],stage3_15[31]}
   );
   gpc615_5 gpc1722 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[32]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[7],stage3_17[7],stage3_16[20],stage3_15[32]}
   );
   gpc615_5 gpc1723 (
      {stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23], stage2_15[24]},
      {stage2_16[33]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[8],stage3_17[8],stage3_16[21],stage3_15[33]}
   );
   gpc615_5 gpc1724 (
      {stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage2_16[34]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[9],stage3_17[9],stage3_16[22],stage3_15[34]}
   );
   gpc615_5 gpc1725 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[35]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[10],stage3_17[10],stage3_16[23],stage3_15[35]}
   );
   gpc615_5 gpc1726 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[36]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[11],stage3_17[11],stage3_16[24],stage3_15[36]}
   );
   gpc615_5 gpc1727 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[37]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[12],stage3_17[12],stage3_16[25],stage3_15[37]}
   );
   gpc615_5 gpc1728 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[38]},
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage3_19[8],stage3_18[13],stage3_17[13],stage3_16[26],stage3_15[38]}
   );
   gpc615_5 gpc1729 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[39]},
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage3_19[9],stage3_18[14],stage3_17[14],stage3_16[27],stage3_15[39]}
   );
   gpc615_5 gpc1730 (
      {stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59]},
      {stage2_16[40]},
      {stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65]},
      {stage3_19[10],stage3_18[15],stage3_17[15],stage3_16[28],stage3_15[40]}
   );
   gpc615_5 gpc1731 (
      {stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_16[41]},
      {stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71]},
      {stage3_19[11],stage3_18[16],stage3_17[16],stage3_16[29],stage3_15[41]}
   );
   gpc615_5 gpc1732 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69]},
      {stage2_16[42]},
      {stage2_17[72], stage2_17[73], stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77]},
      {stage3_19[12],stage3_18[17],stage3_17[17],stage3_16[30],stage3_15[42]}
   );
   gpc615_5 gpc1733 (
      {stage2_15[70], stage2_15[71], stage2_15[72], stage2_15[73], stage2_15[74]},
      {stage2_16[43]},
      {stage2_17[78], stage2_17[79], stage2_17[80], stage2_17[81], stage2_17[82], stage2_17[83]},
      {stage3_19[13],stage3_18[18],stage3_17[18],stage3_16[31],stage3_15[43]}
   );
   gpc606_5 gpc1734 (
      {stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47], stage2_16[48], stage2_16[49]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[14],stage3_18[19],stage3_17[19],stage3_16[32]}
   );
   gpc606_5 gpc1735 (
      {stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53], stage2_16[54], stage2_16[55]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[15],stage3_18[20],stage3_17[20],stage3_16[33]}
   );
   gpc606_5 gpc1736 (
      {stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59], stage2_16[60], stage2_16[61]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[16],stage3_18[21],stage3_17[21],stage3_16[34]}
   );
   gpc606_5 gpc1737 (
      {stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65], stage2_16[66], stage2_16[67]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[17],stage3_18[22],stage3_17[22],stage3_16[35]}
   );
   gpc606_5 gpc1738 (
      {stage2_17[84], stage2_17[85], stage2_17[86], stage2_17[87], stage2_17[88], stage2_17[89]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], 1'b0},
      {stage3_21[0],stage3_20[4],stage3_19[18],stage3_18[23],stage3_17[23]}
   );
   gpc1_1 gpc1739 (
      {stage2_0[24]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1740 (
      {stage2_0[25]},
      {stage3_0[7]}
   );
   gpc1_1 gpc1741 (
      {stage2_0[26]},
      {stage3_0[8]}
   );
   gpc1_1 gpc1742 (
      {stage2_0[27]},
      {stage3_0[9]}
   );
   gpc1_1 gpc1743 (
      {stage2_0[28]},
      {stage3_0[10]}
   );
   gpc1_1 gpc1744 (
      {stage2_0[29]},
      {stage3_0[11]}
   );
   gpc1_1 gpc1745 (
      {stage2_0[30]},
      {stage3_0[12]}
   );
   gpc1_1 gpc1746 (
      {stage2_0[31]},
      {stage3_0[13]}
   );
   gpc1_1 gpc1747 (
      {stage2_0[32]},
      {stage3_0[14]}
   );
   gpc1_1 gpc1748 (
      {stage2_0[33]},
      {stage3_0[15]}
   );
   gpc1_1 gpc1749 (
      {stage2_0[34]},
      {stage3_0[16]}
   );
   gpc1_1 gpc1750 (
      {stage2_0[35]},
      {stage3_0[17]}
   );
   gpc1_1 gpc1751 (
      {stage2_0[36]},
      {stage3_0[18]}
   );
   gpc1_1 gpc1752 (
      {stage2_0[37]},
      {stage3_0[19]}
   );
   gpc1_1 gpc1753 (
      {stage2_1[60]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1754 (
      {stage2_1[61]},
      {stage3_1[13]}
   );
   gpc1_1 gpc1755 (
      {stage2_1[62]},
      {stage3_1[14]}
   );
   gpc1_1 gpc1756 (
      {stage2_3[69]},
      {stage3_3[24]}
   );
   gpc1_1 gpc1757 (
      {stage2_3[70]},
      {stage3_3[25]}
   );
   gpc1_1 gpc1758 (
      {stage2_3[71]},
      {stage3_3[26]}
   );
   gpc1_1 gpc1759 (
      {stage2_3[72]},
      {stage3_3[27]}
   );
   gpc1_1 gpc1760 (
      {stage2_3[73]},
      {stage3_3[28]}
   );
   gpc1_1 gpc1761 (
      {stage2_3[74]},
      {stage3_3[29]}
   );
   gpc1_1 gpc1762 (
      {stage2_3[75]},
      {stage3_3[30]}
   );
   gpc1_1 gpc1763 (
      {stage2_3[76]},
      {stage3_3[31]}
   );
   gpc1_1 gpc1764 (
      {stage2_3[77]},
      {stage3_3[32]}
   );
   gpc1_1 gpc1765 (
      {stage2_3[78]},
      {stage3_3[33]}
   );
   gpc1_1 gpc1766 (
      {stage2_3[79]},
      {stage3_3[34]}
   );
   gpc1_1 gpc1767 (
      {stage2_3[80]},
      {stage3_3[35]}
   );
   gpc1_1 gpc1768 (
      {stage2_3[81]},
      {stage3_3[36]}
   );
   gpc1_1 gpc1769 (
      {stage2_3[82]},
      {stage3_3[37]}
   );
   gpc1_1 gpc1770 (
      {stage2_3[83]},
      {stage3_3[38]}
   );
   gpc1_1 gpc1771 (
      {stage2_3[84]},
      {stage3_3[39]}
   );
   gpc1_1 gpc1772 (
      {stage2_3[85]},
      {stage3_3[40]}
   );
   gpc1_1 gpc1773 (
      {stage2_4[101]},
      {stage3_4[33]}
   );
   gpc1_1 gpc1774 (
      {stage2_4[102]},
      {stage3_4[34]}
   );
   gpc1_1 gpc1775 (
      {stage2_4[103]},
      {stage3_4[35]}
   );
   gpc1_1 gpc1776 (
      {stage2_4[104]},
      {stage3_4[36]}
   );
   gpc1_1 gpc1777 (
      {stage2_4[105]},
      {stage3_4[37]}
   );
   gpc1_1 gpc1778 (
      {stage2_4[106]},
      {stage3_4[38]}
   );
   gpc1_1 gpc1779 (
      {stage2_6[79]},
      {stage3_6[39]}
   );
   gpc1_1 gpc1780 (
      {stage2_6[80]},
      {stage3_6[40]}
   );
   gpc1_1 gpc1781 (
      {stage2_6[81]},
      {stage3_6[41]}
   );
   gpc1_1 gpc1782 (
      {stage2_6[82]},
      {stage3_6[42]}
   );
   gpc1_1 gpc1783 (
      {stage2_6[83]},
      {stage3_6[43]}
   );
   gpc1_1 gpc1784 (
      {stage2_6[84]},
      {stage3_6[44]}
   );
   gpc1_1 gpc1785 (
      {stage2_6[85]},
      {stage3_6[45]}
   );
   gpc1_1 gpc1786 (
      {stage2_6[86]},
      {stage3_6[46]}
   );
   gpc1_1 gpc1787 (
      {stage2_6[87]},
      {stage3_6[47]}
   );
   gpc1_1 gpc1788 (
      {stage2_6[88]},
      {stage3_6[48]}
   );
   gpc1_1 gpc1789 (
      {stage2_6[89]},
      {stage3_6[49]}
   );
   gpc1_1 gpc1790 (
      {stage2_8[100]},
      {stage3_8[42]}
   );
   gpc1_1 gpc1791 (
      {stage2_8[101]},
      {stage3_8[43]}
   );
   gpc1_1 gpc1792 (
      {stage2_8[102]},
      {stage3_8[44]}
   );
   gpc1_1 gpc1793 (
      {stage2_8[103]},
      {stage3_8[45]}
   );
   gpc1_1 gpc1794 (
      {stage2_8[104]},
      {stage3_8[46]}
   );
   gpc1_1 gpc1795 (
      {stage2_8[105]},
      {stage3_8[47]}
   );
   gpc1_1 gpc1796 (
      {stage2_9[80]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1797 (
      {stage2_10[77]},
      {stage3_10[31]}
   );
   gpc1_1 gpc1798 (
      {stage2_10[78]},
      {stage3_10[32]}
   );
   gpc1_1 gpc1799 (
      {stage2_10[79]},
      {stage3_10[33]}
   );
   gpc1_1 gpc1800 (
      {stage2_10[80]},
      {stage3_10[34]}
   );
   gpc1_1 gpc1801 (
      {stage2_10[81]},
      {stage3_10[35]}
   );
   gpc1_1 gpc1802 (
      {stage2_10[82]},
      {stage3_10[36]}
   );
   gpc1_1 gpc1803 (
      {stage2_10[83]},
      {stage3_10[37]}
   );
   gpc1_1 gpc1804 (
      {stage2_10[84]},
      {stage3_10[38]}
   );
   gpc1_1 gpc1805 (
      {stage2_10[85]},
      {stage3_10[39]}
   );
   gpc1_1 gpc1806 (
      {stage2_10[86]},
      {stage3_10[40]}
   );
   gpc1_1 gpc1807 (
      {stage2_10[87]},
      {stage3_10[41]}
   );
   gpc1_1 gpc1808 (
      {stage2_10[88]},
      {stage3_10[42]}
   );
   gpc1_1 gpc1809 (
      {stage2_10[89]},
      {stage3_10[43]}
   );
   gpc1_1 gpc1810 (
      {stage2_13[80]},
      {stage3_13[34]}
   );
   gpc1_1 gpc1811 (
      {stage2_13[81]},
      {stage3_13[35]}
   );
   gpc1_1 gpc1812 (
      {stage2_13[82]},
      {stage3_13[36]}
   );
   gpc1_1 gpc1813 (
      {stage2_13[83]},
      {stage3_13[37]}
   );
   gpc1_1 gpc1814 (
      {stage2_13[84]},
      {stage3_13[38]}
   );
   gpc1_1 gpc1815 (
      {stage2_13[85]},
      {stage3_13[39]}
   );
   gpc1_1 gpc1816 (
      {stage2_16[68]},
      {stage3_16[36]}
   );
   gpc1_1 gpc1817 (
      {stage2_16[69]},
      {stage3_16[37]}
   );
   gpc1_1 gpc1818 (
      {stage2_16[70]},
      {stage3_16[38]}
   );
   gpc1_1 gpc1819 (
      {stage2_16[71]},
      {stage3_16[39]}
   );
   gpc1_1 gpc1820 (
      {stage2_16[72]},
      {stage3_16[40]}
   );
   gpc1_1 gpc1821 (
      {stage2_16[73]},
      {stage3_16[41]}
   );
   gpc1_1 gpc1822 (
      {stage2_16[74]},
      {stage3_16[42]}
   );
   gpc1_1 gpc1823 (
      {stage2_16[75]},
      {stage3_16[43]}
   );
   gpc1_1 gpc1824 (
      {stage2_16[76]},
      {stage3_16[44]}
   );
   gpc1_1 gpc1825 (
      {stage2_17[90]},
      {stage3_17[24]}
   );
   gpc1_1 gpc1826 (
      {stage2_17[91]},
      {stage3_17[25]}
   );
   gpc1_1 gpc1827 (
      {stage2_17[92]},
      {stage3_17[26]}
   );
   gpc1_1 gpc1828 (
      {stage2_17[93]},
      {stage3_17[27]}
   );
   gpc1_1 gpc1829 (
      {stage2_17[94]},
      {stage3_17[28]}
   );
   gpc1_1 gpc1830 (
      {stage2_17[95]},
      {stage3_17[29]}
   );
   gpc1_1 gpc1831 (
      {stage2_18[24]},
      {stage3_18[24]}
   );
   gpc1_1 gpc1832 (
      {stage2_18[25]},
      {stage3_18[25]}
   );
   gpc1406_5 gpc1833 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1834 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10], stage3_0[11]},
      {stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1343_5 gpc1835 (
      {stage3_1[0], stage3_1[1], stage3_1[2]},
      {stage3_2[10], stage3_2[11], stage3_2[12], stage3_2[13]},
      {stage3_3[1], stage3_3[2], stage3_3[3]},
      {stage3_4[0]},
      {stage4_5[0],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc1836 (
      {stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8]},
      {stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9]},
      {stage4_5[1],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc615_5 gpc1837 (
      {stage3_1[9], stage3_1[10], stage3_1[11], stage3_1[12], stage3_1[13]},
      {stage3_2[14]},
      {stage3_3[10], stage3_3[11], stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15]},
      {stage4_5[2],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc615_5 gpc1838 (
      {stage3_3[16], stage3_3[17], stage3_3[18], stage3_3[19], stage3_3[20]},
      {stage3_4[1]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[3],stage4_4[5],stage4_3[5]}
   );
   gpc615_5 gpc1839 (
      {stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24], stage3_3[25]},
      {stage3_4[2]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[4],stage4_4[6],stage4_3[6]}
   );
   gpc615_5 gpc1840 (
      {stage3_3[26], stage3_3[27], stage3_3[28], stage3_3[29], stage3_3[30]},
      {stage3_4[3]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[2],stage4_5[5],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc1841 (
      {stage3_3[31], stage3_3[32], stage3_3[33], stage3_3[34], stage3_3[35]},
      {stage3_4[4]},
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage4_7[3],stage4_6[3],stage4_5[6],stage4_4[8],stage4_3[8]}
   );
   gpc615_5 gpc1842 (
      {stage3_3[36], stage3_3[37], stage3_3[38], stage3_3[39], stage3_3[40]},
      {stage3_4[5]},
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage4_7[4],stage4_6[4],stage4_5[7],stage4_4[9],stage4_3[9]}
   );
   gpc1415_5 gpc1843 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[30]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[5],stage4_6[5],stage4_5[8],stage4_4[10]}
   );
   gpc606_5 gpc1844 (
      {stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16]},
      {stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage4_8[1],stage4_7[6],stage4_6[6],stage4_5[9],stage4_4[11]}
   );
   gpc606_5 gpc1845 (
      {stage3_4[17], stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22]},
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage4_8[2],stage4_7[7],stage4_6[7],stage4_5[10],stage4_4[12]}
   );
   gpc615_5 gpc1846 (
      {stage3_4[23], stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27]},
      {stage3_5[31]},
      {stage3_6[16], stage3_6[17], stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21]},
      {stage4_8[3],stage4_7[8],stage4_6[8],stage4_5[11],stage4_4[13]}
   );
   gpc615_5 gpc1847 (
      {stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_5[32]},
      {stage3_6[22], stage3_6[23], stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27]},
      {stage4_8[4],stage4_7[9],stage4_6[9],stage4_5[12],stage4_4[14]}
   );
   gpc615_5 gpc1848 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37]},
      {stage3_5[33]},
      {stage3_6[28], stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage4_8[5],stage4_7[10],stage4_6[10],stage4_5[13],stage4_4[15]}
   );
   gpc606_5 gpc1849 (
      {stage3_5[34], stage3_5[35], stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39]},
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage4_9[0],stage4_8[6],stage4_7[11],stage4_6[11],stage4_5[14]}
   );
   gpc615_5 gpc1850 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[7]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[7],stage4_7[12],stage4_6[12]}
   );
   gpc615_5 gpc1851 (
      {stage3_6[39], stage3_6[40], stage3_6[41], stage3_6[42], stage3_6[43]},
      {stage3_7[8]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[8],stage4_7[13],stage4_6[13]}
   );
   gpc615_5 gpc1852 (
      {stage3_6[44], stage3_6[45], stage3_6[46], stage3_6[47], stage3_6[48]},
      {stage3_7[9]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[3],stage4_8[9],stage4_7[14],stage4_6[14]}
   );
   gpc615_5 gpc1853 (
      {stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_8[18]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[3],stage4_9[4],stage4_8[10],stage4_7[15]}
   );
   gpc615_5 gpc1854 (
      {stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage3_8[19]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[4],stage4_9[5],stage4_8[11],stage4_7[16]}
   );
   gpc615_5 gpc1855 (
      {stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23], stage3_7[24]},
      {stage3_8[20]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[5],stage4_9[6],stage4_8[12],stage4_7[17]}
   );
   gpc615_5 gpc1856 (
      {stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage3_8[21]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[6],stage4_9[7],stage4_8[13],stage4_7[18]}
   );
   gpc615_5 gpc1857 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[22]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[7],stage4_9[8],stage4_8[14],stage4_7[19]}
   );
   gpc606_5 gpc1858 (
      {stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[5],stage4_10[8],stage4_9[9],stage4_8[15]}
   );
   gpc606_5 gpc1859 (
      {stage3_8[29], stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[6],stage4_10[9],stage4_9[10],stage4_8[16]}
   );
   gpc606_5 gpc1860 (
      {stage3_8[35], stage3_8[36], stage3_8[37], stage3_8[38], stage3_8[39], stage3_8[40]},
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage4_12[2],stage4_11[7],stage4_10[10],stage4_9[11],stage4_8[17]}
   );
   gpc606_5 gpc1861 (
      {stage3_8[41], stage3_8[42], stage3_8[43], stage3_8[44], stage3_8[45], stage3_8[46]},
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23]},
      {stage4_12[3],stage4_11[8],stage4_10[11],stage4_9[12],stage4_8[18]}
   );
   gpc606_5 gpc1862 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[4],stage4_11[9],stage4_10[12],stage4_9[13]}
   );
   gpc606_5 gpc1863 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[5],stage4_11[10],stage4_10[13],stage4_9[14]}
   );
   gpc615_5 gpc1864 (
      {stage3_10[24], stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[6],stage4_11[11],stage4_10[14]}
   );
   gpc615_5 gpc1865 (
      {stage3_10[29], stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33]},
      {stage3_11[13]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[3],stage4_12[7],stage4_11[12],stage4_10[15]}
   );
   gpc615_5 gpc1866 (
      {stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38]},
      {stage3_11[14]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[4],stage4_12[8],stage4_11[13],stage4_10[16]}
   );
   gpc615_5 gpc1867 (
      {stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_11[15]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[5],stage4_12[9],stage4_11[14],stage4_10[17]}
   );
   gpc606_5 gpc1868 (
      {stage3_11[16], stage3_11[17], stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[4],stage4_13[6],stage4_12[10],stage4_11[15]}
   );
   gpc606_5 gpc1869 (
      {stage3_11[22], stage3_11[23], stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[5],stage4_13[7],stage4_12[11],stage4_11[16]}
   );
   gpc615_5 gpc1870 (
      {stage3_11[28], stage3_11[29], stage3_11[30], stage3_11[31], stage3_11[32]},
      {stage3_12[24]},
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage4_15[2],stage4_14[6],stage4_13[8],stage4_12[12],stage4_11[17]}
   );
   gpc615_5 gpc1871 (
      {stage3_11[33], stage3_11[34], stage3_11[35], stage3_11[36], stage3_11[37]},
      {stage3_12[25]},
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23]},
      {stage4_15[3],stage4_14[7],stage4_13[9],stage4_12[13],stage4_11[18]}
   );
   gpc117_4 gpc1872 (
      {stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29], stage3_12[30], stage3_12[31], stage3_12[32]},
      {stage3_13[24]},
      {stage3_14[0]},
      {stage4_15[4],stage4_14[8],stage4_13[10],stage4_12[14]}
   );
   gpc606_5 gpc1873 (
      {stage3_12[33], stage3_12[34], stage3_12[35], stage3_12[36], stage3_12[37], stage3_12[38]},
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage4_16[0],stage4_15[5],stage4_14[9],stage4_13[11],stage4_12[15]}
   );
   gpc606_5 gpc1874 (
      {stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[6],stage4_14[10],stage4_13[12]}
   );
   gpc606_5 gpc1875 (
      {stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[7],stage4_14[11],stage4_13[13]}
   );
   gpc606_5 gpc1876 (
      {stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11], stage3_14[12]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[8],stage4_14[12]}
   );
   gpc615_5 gpc1877 (
      {stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage3_15[12]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[9],stage4_14[13]}
   );
   gpc615_5 gpc1878 (
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22]},
      {stage3_15[13]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[10],stage4_14[14]}
   );
   gpc615_5 gpc1879 (
      {stage3_14[23], stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27]},
      {stage3_15[14]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[11],stage4_14[15]}
   );
   gpc606_5 gpc1880 (
      {stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[12]}
   );
   gpc615_5 gpc1881 (
      {stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25]},
      {stage3_16[24]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[5],stage4_17[7],stage4_16[8],stage4_15[13]}
   );
   gpc615_5 gpc1882 (
      {stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30]},
      {stage3_16[25]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[6],stage4_17[8],stage4_16[9],stage4_15[14]}
   );
   gpc606_5 gpc1883 (
      {stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29], stage3_16[30], stage3_16[31]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[7],stage4_17[9],stage4_16[10]}
   );
   gpc606_5 gpc1884 (
      {stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35], stage3_16[36], stage3_16[37]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[8],stage4_17[10],stage4_16[11]}
   );
   gpc606_5 gpc1885 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[2],stage4_19[5],stage4_18[9],stage4_17[11]}
   );
   gpc606_5 gpc1886 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[3],stage4_19[6],stage4_18[10],stage4_17[12]}
   );
   gpc1_1 gpc1887 (
      {stage3_0[12]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1888 (
      {stage3_0[13]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1889 (
      {stage3_0[14]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1890 (
      {stage3_0[15]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1891 (
      {stage3_0[16]},
      {stage4_0[6]}
   );
   gpc1_1 gpc1892 (
      {stage3_0[17]},
      {stage4_0[7]}
   );
   gpc1_1 gpc1893 (
      {stage3_0[18]},
      {stage4_0[8]}
   );
   gpc1_1 gpc1894 (
      {stage3_0[19]},
      {stage4_0[9]}
   );
   gpc1_1 gpc1895 (
      {stage3_1[14]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1896 (
      {stage3_2[15]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1897 (
      {stage3_2[16]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1898 (
      {stage3_2[17]},
      {stage4_2[7]}
   );
   gpc1_1 gpc1899 (
      {stage3_2[18]},
      {stage4_2[8]}
   );
   gpc1_1 gpc1900 (
      {stage3_4[38]},
      {stage4_4[16]}
   );
   gpc1_1 gpc1901 (
      {stage3_6[49]},
      {stage4_6[15]}
   );
   gpc1_1 gpc1902 (
      {stage3_7[35]},
      {stage4_7[20]}
   );
   gpc1_1 gpc1903 (
      {stage3_8[47]},
      {stage4_8[19]}
   );
   gpc1_1 gpc1904 (
      {stage3_9[42]},
      {stage4_9[15]}
   );
   gpc1_1 gpc1905 (
      {stage3_12[39]},
      {stage4_12[16]}
   );
   gpc1_1 gpc1906 (
      {stage3_12[40]},
      {stage4_12[17]}
   );
   gpc1_1 gpc1907 (
      {stage3_12[41]},
      {stage4_12[18]}
   );
   gpc1_1 gpc1908 (
      {stage3_12[42]},
      {stage4_12[19]}
   );
   gpc1_1 gpc1909 (
      {stage3_12[43]},
      {stage4_12[20]}
   );
   gpc1_1 gpc1910 (
      {stage3_12[44]},
      {stage4_12[21]}
   );
   gpc1_1 gpc1911 (
      {stage3_12[45]},
      {stage4_12[22]}
   );
   gpc1_1 gpc1912 (
      {stage3_12[46]},
      {stage4_12[23]}
   );
   gpc1_1 gpc1913 (
      {stage3_13[37]},
      {stage4_13[14]}
   );
   gpc1_1 gpc1914 (
      {stage3_13[38]},
      {stage4_13[15]}
   );
   gpc1_1 gpc1915 (
      {stage3_13[39]},
      {stage4_13[16]}
   );
   gpc1_1 gpc1916 (
      {stage3_14[28]},
      {stage4_14[16]}
   );
   gpc1_1 gpc1917 (
      {stage3_14[29]},
      {stage4_14[17]}
   );
   gpc1_1 gpc1918 (
      {stage3_14[30]},
      {stage4_14[18]}
   );
   gpc1_1 gpc1919 (
      {stage3_14[31]},
      {stage4_14[19]}
   );
   gpc1_1 gpc1920 (
      {stage3_15[31]},
      {stage4_15[15]}
   );
   gpc1_1 gpc1921 (
      {stage3_15[32]},
      {stage4_15[16]}
   );
   gpc1_1 gpc1922 (
      {stage3_15[33]},
      {stage4_15[17]}
   );
   gpc1_1 gpc1923 (
      {stage3_15[34]},
      {stage4_15[18]}
   );
   gpc1_1 gpc1924 (
      {stage3_15[35]},
      {stage4_15[19]}
   );
   gpc1_1 gpc1925 (
      {stage3_15[36]},
      {stage4_15[20]}
   );
   gpc1_1 gpc1926 (
      {stage3_15[37]},
      {stage4_15[21]}
   );
   gpc1_1 gpc1927 (
      {stage3_15[38]},
      {stage4_15[22]}
   );
   gpc1_1 gpc1928 (
      {stage3_15[39]},
      {stage4_15[23]}
   );
   gpc1_1 gpc1929 (
      {stage3_15[40]},
      {stage4_15[24]}
   );
   gpc1_1 gpc1930 (
      {stage3_15[41]},
      {stage4_15[25]}
   );
   gpc1_1 gpc1931 (
      {stage3_15[42]},
      {stage4_15[26]}
   );
   gpc1_1 gpc1932 (
      {stage3_15[43]},
      {stage4_15[27]}
   );
   gpc1_1 gpc1933 (
      {stage3_16[38]},
      {stage4_16[12]}
   );
   gpc1_1 gpc1934 (
      {stage3_16[39]},
      {stage4_16[13]}
   );
   gpc1_1 gpc1935 (
      {stage3_16[40]},
      {stage4_16[14]}
   );
   gpc1_1 gpc1936 (
      {stage3_16[41]},
      {stage4_16[15]}
   );
   gpc1_1 gpc1937 (
      {stage3_16[42]},
      {stage4_16[16]}
   );
   gpc1_1 gpc1938 (
      {stage3_16[43]},
      {stage4_16[17]}
   );
   gpc1_1 gpc1939 (
      {stage3_16[44]},
      {stage4_16[18]}
   );
   gpc1_1 gpc1940 (
      {stage3_18[12]},
      {stage4_18[11]}
   );
   gpc1_1 gpc1941 (
      {stage3_18[13]},
      {stage4_18[12]}
   );
   gpc1_1 gpc1942 (
      {stage3_18[14]},
      {stage4_18[13]}
   );
   gpc1_1 gpc1943 (
      {stage3_18[15]},
      {stage4_18[14]}
   );
   gpc1_1 gpc1944 (
      {stage3_18[16]},
      {stage4_18[15]}
   );
   gpc1_1 gpc1945 (
      {stage3_18[17]},
      {stage4_18[16]}
   );
   gpc1_1 gpc1946 (
      {stage3_18[18]},
      {stage4_18[17]}
   );
   gpc1_1 gpc1947 (
      {stage3_18[19]},
      {stage4_18[18]}
   );
   gpc1_1 gpc1948 (
      {stage3_18[20]},
      {stage4_18[19]}
   );
   gpc1_1 gpc1949 (
      {stage3_18[21]},
      {stage4_18[20]}
   );
   gpc1_1 gpc1950 (
      {stage3_18[22]},
      {stage4_18[21]}
   );
   gpc1_1 gpc1951 (
      {stage3_18[23]},
      {stage4_18[22]}
   );
   gpc1_1 gpc1952 (
      {stage3_18[24]},
      {stage4_18[23]}
   );
   gpc1_1 gpc1953 (
      {stage3_18[25]},
      {stage4_18[24]}
   );
   gpc1_1 gpc1954 (
      {stage3_19[12]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1955 (
      {stage3_19[13]},
      {stage4_19[8]}
   );
   gpc1_1 gpc1956 (
      {stage3_19[14]},
      {stage4_19[9]}
   );
   gpc1_1 gpc1957 (
      {stage3_19[15]},
      {stage4_19[10]}
   );
   gpc1_1 gpc1958 (
      {stage3_19[16]},
      {stage4_19[11]}
   );
   gpc1_1 gpc1959 (
      {stage3_19[17]},
      {stage4_19[12]}
   );
   gpc1_1 gpc1960 (
      {stage3_19[18]},
      {stage4_19[13]}
   );
   gpc1_1 gpc1961 (
      {stage3_20[0]},
      {stage4_20[4]}
   );
   gpc1_1 gpc1962 (
      {stage3_20[1]},
      {stage4_20[5]}
   );
   gpc1_1 gpc1963 (
      {stage3_20[2]},
      {stage4_20[6]}
   );
   gpc1_1 gpc1964 (
      {stage3_20[3]},
      {stage4_20[7]}
   );
   gpc1_1 gpc1965 (
      {stage3_20[4]},
      {stage4_20[8]}
   );
   gpc1_1 gpc1966 (
      {stage3_21[0]},
      {stage4_21[2]}
   );
   gpc615_5 gpc1967 (
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4]},
      {stage4_4[0]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0]}
   );
   gpc2135_5 gpc1968 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[6], stage4_5[7], stage4_5[8]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[1],stage5_6[1],stage5_5[1],stage5_4[1]}
   );
   gpc2135_5 gpc1969 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10]},
      {stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_6[1]},
      {stage4_7[2], stage4_7[3]},
      {stage5_8[1],stage5_7[2],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc2135_5 gpc1970 (
      {stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_5[12], stage4_5[13], stage4_5[14]},
      {stage4_6[2]},
      {stage4_7[4], stage4_7[5]},
      {stage5_8[2],stage5_7[3],stage5_6[3],stage5_5[3],stage5_4[3]}
   );
   gpc615_5 gpc1971 (
      {stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[3],stage5_7[4],stage5_6[4]}
   );
   gpc615_5 gpc1972 (
      {stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12]},
      {stage4_7[7]},
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage5_10[1],stage5_9[1],stage5_8[4],stage5_7[5],stage5_6[5]}
   );
   gpc2116_5 gpc1973 (
      {stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11], stage4_7[12], stage4_7[13]},
      {stage4_8[12]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[5],stage5_7[6]}
   );
   gpc606_5 gpc1974 (
      {stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17], stage4_7[18], stage4_7[19]},
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[6],stage5_7[7]}
   );
   gpc623_5 gpc1975 (
      {stage4_9[7], stage4_9[8], stage4_9[9]},
      {stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[4]}
   );
   gpc623_5 gpc1976 (
      {stage4_9[10], stage4_9[11], stage4_9[12]},
      {stage4_10[4], stage4_10[5]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[5]}
   );
   gpc606_5 gpc1977 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[4],stage5_10[6]}
   );
   gpc606_5 gpc1978 (
      {stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[3],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc7_3 gpc1979 (
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17], stage4_11[18]},
      {stage5_13[4],stage5_12[4],stage5_11[6]}
   );
   gpc606_5 gpc1980 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[5],stage5_12[5]}
   );
   gpc606_5 gpc1981 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[1],stage5_14[3],stage5_13[6],stage5_12[6]}
   );
   gpc606_5 gpc1982 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[2],stage5_15[2],stage5_14[4],stage5_13[7]}
   );
   gpc606_5 gpc1983 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[3],stage5_15[3],stage5_14[5],stage5_13[8]}
   );
   gpc615_5 gpc1984 (
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16]},
      {stage4_14[12]},
      {stage4_15[12], stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17]},
      {stage5_17[2],stage5_16[4],stage5_15[4],stage5_14[6],stage5_13[9]}
   );
   gpc7_3 gpc1985 (
      {stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19]},
      {stage5_16[5],stage5_15[5],stage5_14[7]}
   );
   gpc1163_5 gpc1986 (
      {stage4_15[18], stage4_15[19], stage4_15[20]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0]},
      {stage4_18[0]},
      {stage5_19[0],stage5_18[0],stage5_17[3],stage5_16[6],stage5_15[6]}
   );
   gpc615_5 gpc1987 (
      {stage4_15[21], stage4_15[22], stage4_15[23], stage4_15[24], stage4_15[25]},
      {stage4_16[6]},
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6]},
      {stage5_19[1],stage5_18[1],stage5_17[4],stage5_16[7],stage5_15[7]}
   );
   gpc606_5 gpc1988 (
      {stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12]},
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[0],stage5_19[2],stage5_18[2],stage5_17[5],stage5_16[8]}
   );
   gpc606_5 gpc1989 (
      {stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11], stage4_18[12]},
      {stage5_20[1],stage5_19[3],stage5_18[3],stage5_17[6],stage5_16[9]}
   );
   gpc606_5 gpc1990 (
      {stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11], stage4_17[12]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[2],stage5_19[4],stage5_18[4],stage5_17[7]}
   );
   gpc2135_5 gpc1991 (
      {stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[0]},
      {stage4_21[0], stage4_21[1]},
      {stage5_22[0],stage5_21[1],stage5_20[3],stage5_19[5],stage5_18[5]}
   );
   gpc117_4 gpc1992 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22], stage4_18[23], stage4_18[24]},
      {stage4_19[9]},
      {stage4_20[1]},
      {stage5_21[2],stage5_20[4],stage5_19[6],stage5_18[6]}
   );
   gpc1_1 gpc1993 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1994 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1995 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc1996 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc1997 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc1998 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc1999 (
      {stage4_0[6]},
      {stage5_0[6]}
   );
   gpc1_1 gpc2000 (
      {stage4_0[7]},
      {stage5_0[7]}
   );
   gpc1_1 gpc2001 (
      {stage4_0[8]},
      {stage5_0[8]}
   );
   gpc1_1 gpc2002 (
      {stage4_0[9]},
      {stage5_0[9]}
   );
   gpc1_1 gpc2003 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2004 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2005 (
      {stage4_1[2]},
      {stage5_1[2]}
   );
   gpc1_1 gpc2006 (
      {stage4_1[3]},
      {stage5_1[3]}
   );
   gpc1_1 gpc2007 (
      {stage4_1[4]},
      {stage5_1[4]}
   );
   gpc1_1 gpc2008 (
      {stage4_1[5]},
      {stage5_1[5]}
   );
   gpc1_1 gpc2009 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc2010 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2011 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc2012 (
      {stage4_2[3]},
      {stage5_2[3]}
   );
   gpc1_1 gpc2013 (
      {stage4_2[4]},
      {stage5_2[4]}
   );
   gpc1_1 gpc2014 (
      {stage4_2[5]},
      {stage5_2[5]}
   );
   gpc1_1 gpc2015 (
      {stage4_2[6]},
      {stage5_2[6]}
   );
   gpc1_1 gpc2016 (
      {stage4_2[7]},
      {stage5_2[7]}
   );
   gpc1_1 gpc2017 (
      {stage4_2[8]},
      {stage5_2[8]}
   );
   gpc1_1 gpc2018 (
      {stage4_3[5]},
      {stage5_3[1]}
   );
   gpc1_1 gpc2019 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2020 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2021 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc2022 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc2023 (
      {stage4_4[16]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2024 (
      {stage4_6[13]},
      {stage5_6[6]}
   );
   gpc1_1 gpc2025 (
      {stage4_6[14]},
      {stage5_6[7]}
   );
   gpc1_1 gpc2026 (
      {stage4_6[15]},
      {stage5_6[8]}
   );
   gpc1_1 gpc2027 (
      {stage4_7[20]},
      {stage5_7[8]}
   );
   gpc1_1 gpc2028 (
      {stage4_8[13]},
      {stage5_8[7]}
   );
   gpc1_1 gpc2029 (
      {stage4_8[14]},
      {stage5_8[8]}
   );
   gpc1_1 gpc2030 (
      {stage4_8[15]},
      {stage5_8[9]}
   );
   gpc1_1 gpc2031 (
      {stage4_8[16]},
      {stage5_8[10]}
   );
   gpc1_1 gpc2032 (
      {stage4_8[17]},
      {stage5_8[11]}
   );
   gpc1_1 gpc2033 (
      {stage4_8[18]},
      {stage5_8[12]}
   );
   gpc1_1 gpc2034 (
      {stage4_8[19]},
      {stage5_8[13]}
   );
   gpc1_1 gpc2035 (
      {stage4_9[13]},
      {stage5_9[6]}
   );
   gpc1_1 gpc2036 (
      {stage4_9[14]},
      {stage5_9[7]}
   );
   gpc1_1 gpc2037 (
      {stage4_9[15]},
      {stage5_9[8]}
   );
   gpc1_1 gpc2038 (
      {stage4_15[26]},
      {stage5_15[8]}
   );
   gpc1_1 gpc2039 (
      {stage4_15[27]},
      {stage5_15[9]}
   );
   gpc1_1 gpc2040 (
      {stage4_19[10]},
      {stage5_19[7]}
   );
   gpc1_1 gpc2041 (
      {stage4_19[11]},
      {stage5_19[8]}
   );
   gpc1_1 gpc2042 (
      {stage4_19[12]},
      {stage5_19[9]}
   );
   gpc1_1 gpc2043 (
      {stage4_19[13]},
      {stage5_19[10]}
   );
   gpc1_1 gpc2044 (
      {stage4_20[2]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2045 (
      {stage4_20[3]},
      {stage5_20[6]}
   );
   gpc1_1 gpc2046 (
      {stage4_20[4]},
      {stage5_20[7]}
   );
   gpc1_1 gpc2047 (
      {stage4_20[5]},
      {stage5_20[8]}
   );
   gpc1_1 gpc2048 (
      {stage4_20[6]},
      {stage5_20[9]}
   );
   gpc1_1 gpc2049 (
      {stage4_20[7]},
      {stage5_20[10]}
   );
   gpc1_1 gpc2050 (
      {stage4_20[8]},
      {stage5_20[11]}
   );
   gpc1_1 gpc2051 (
      {stage4_21[2]},
      {stage5_21[3]}
   );
   gpc2135_5 gpc2052 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0]},
      {stage5_3[0], stage5_3[1]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc135_4 gpc2053 (
      {stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4], stage5_2[5]},
      {stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[1],stage6_3[1],stage6_2[1]}
   );
   gpc615_5 gpc2054 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[0]}
   );
   gpc623_5 gpc2055 (
      {stage5_6[5], stage5_6[6], stage5_6[7]},
      {stage5_7[1], stage5_7[2]},
      {stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[1],stage6_6[1]}
   );
   gpc615_5 gpc2056 (
      {stage5_7[3], stage5_7[4], stage5_7[5], stage5_7[6], stage5_7[7]},
      {stage5_8[12]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[2],stage6_9[2],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc2057 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[3]}
   );
   gpc615_5 gpc2058 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], stage5_10[7]},
      {stage5_11[6]},
      {stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[2],stage6_10[4]}
   );
   gpc135_4 gpc2059 (
      {stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[2],stage6_13[2]}
   );
   gpc2135_5 gpc2060 (
      {stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6], stage5_14[7]},
      {stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1]},
      {stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[3]}
   );
   gpc606_5 gpc2061 (
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9]},
      {stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7]},
      {stage6_19[0],stage6_18[1],stage6_17[1],stage6_16[2],stage6_15[2]}
   );
   gpc7_3 gpc2062 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7]},
      {stage6_18[2],stage6_17[2],stage6_16[3]}
   );
   gpc615_5 gpc2063 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[0]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[3]}
   );
   gpc2135_5 gpc2064 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_21[0]},
      {stage5_22[0], 1'b0},
      {stage6_23[0],stage6_22[1],stage6_21[1],stage6_20[1],stage6_19[2]}
   );
   gpc615_5 gpc2065 (
      {stage5_19[6], stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10]},
      {stage5_20[9]},
      {stage5_21[1], stage5_21[2], stage5_21[3], 1'b0, 1'b0, 1'b0},
      {stage6_23[1],stage6_22[2],stage6_21[2],stage6_20[2],stage6_19[3]}
   );
   gpc1_1 gpc2066 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc2067 (
      {stage5_0[6]},
      {stage6_0[2]}
   );
   gpc1_1 gpc2068 (
      {stage5_0[7]},
      {stage6_0[3]}
   );
   gpc1_1 gpc2069 (
      {stage5_0[8]},
      {stage6_0[4]}
   );
   gpc1_1 gpc2070 (
      {stage5_0[9]},
      {stage6_0[5]}
   );
   gpc1_1 gpc2071 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2072 (
      {stage5_1[4]},
      {stage6_1[2]}
   );
   gpc1_1 gpc2073 (
      {stage5_1[5]},
      {stage6_1[3]}
   );
   gpc1_1 gpc2074 (
      {stage5_2[6]},
      {stage6_2[2]}
   );
   gpc1_1 gpc2075 (
      {stage5_2[7]},
      {stage6_2[3]}
   );
   gpc1_1 gpc2076 (
      {stage5_2[8]},
      {stage6_2[4]}
   );
   gpc1_1 gpc2077 (
      {stage5_3[5]},
      {stage6_3[2]}
   );
   gpc1_1 gpc2078 (
      {stage5_4[1]},
      {stage6_4[2]}
   );
   gpc1_1 gpc2079 (
      {stage5_4[2]},
      {stage6_4[3]}
   );
   gpc1_1 gpc2080 (
      {stage5_4[3]},
      {stage6_4[4]}
   );
   gpc1_1 gpc2081 (
      {stage5_4[4]},
      {stage6_4[5]}
   );
   gpc1_1 gpc2082 (
      {stage5_5[0]},
      {stage6_5[1]}
   );
   gpc1_1 gpc2083 (
      {stage5_5[1]},
      {stage6_5[2]}
   );
   gpc1_1 gpc2084 (
      {stage5_5[2]},
      {stage6_5[3]}
   );
   gpc1_1 gpc2085 (
      {stage5_5[3]},
      {stage6_5[4]}
   );
   gpc1_1 gpc2086 (
      {stage5_6[8]},
      {stage6_6[2]}
   );
   gpc1_1 gpc2087 (
      {stage5_7[8]},
      {stage6_7[3]}
   );
   gpc1_1 gpc2088 (
      {stage5_8[13]},
      {stage6_8[3]}
   );
   gpc1_1 gpc2089 (
      {stage5_9[6]},
      {stage6_9[3]}
   );
   gpc1_1 gpc2090 (
      {stage5_9[7]},
      {stage6_9[4]}
   );
   gpc1_1 gpc2091 (
      {stage5_9[8]},
      {stage6_9[5]}
   );
   gpc1_1 gpc2092 (
      {stage5_13[6]},
      {stage6_13[3]}
   );
   gpc1_1 gpc2093 (
      {stage5_13[7]},
      {stage6_13[4]}
   );
   gpc1_1 gpc2094 (
      {stage5_13[8]},
      {stage6_13[5]}
   );
   gpc1_1 gpc2095 (
      {stage5_13[9]},
      {stage6_13[6]}
   );
   gpc1_1 gpc2096 (
      {stage5_16[8]},
      {stage6_16[4]}
   );
   gpc1_1 gpc2097 (
      {stage5_16[9]},
      {stage6_16[5]}
   );
   gpc1_1 gpc2098 (
      {stage5_18[5]},
      {stage6_18[4]}
   );
   gpc1_1 gpc2099 (
      {stage5_18[6]},
      {stage6_18[5]}
   );
   gpc1_1 gpc2100 (
      {stage5_20[10]},
      {stage6_20[3]}
   );
   gpc1_1 gpc2101 (
      {stage5_20[11]},
      {stage6_20[4]}
   );
   gpc2135_5 gpc2102 (
      {stage6_0[0], stage6_0[1], stage6_0[2], stage6_0[3], stage6_0[4]},
      {stage6_1[0], stage6_1[1], stage6_1[2]},
      {stage6_2[0]},
      {stage6_3[0], stage6_3[1]},
      {stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0],stage7_0[0]}
   );
   gpc615_5 gpc2103 (
      {stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4], 1'b0},
      {stage6_3[2]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3], stage6_4[4], stage6_4[5]},
      {stage7_6[0],stage7_5[0],stage7_4[1],stage7_3[1],stage7_2[1]}
   );
   gpc135_4 gpc2104 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], stage6_5[4]},
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0]},
      {stage7_8[0],stage7_7[0],stage7_6[1],stage7_5[1]}
   );
   gpc1343_5 gpc2105 (
      {stage6_7[1], stage6_7[2], stage6_7[3]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3]},
      {stage6_9[0], stage6_9[1], stage6_9[2]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[1],stage7_7[1]}
   );
   gpc1343_5 gpc2106 (
      {stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4]},
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0]},
      {stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1],stage7_9[1]}
   );
   gpc117_4 gpc2107 (
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6]},
      {stage6_14[0]},
      {stage6_15[0]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1]}
   );
   gpc623_5 gpc2108 (
      {stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1],stage7_14[1]}
   );
   gpc1163_5 gpc2109 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_19[0]},
      {stage6_20[0]},
      {stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1]}
   );
   gpc1343_5 gpc2110 (
      {stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[0],stage7_21[1],stage7_20[1],stage7_19[1]}
   );
   gpc623_5 gpc2111 (
      {stage6_22[1], stage6_22[2], 1'b0},
      {stage6_23[0], stage6_23[1]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_24[0],stage7_23[1],stage7_22[1]}
   );
   gpc1_1 gpc2112 (
      {stage6_0[5]},
      {stage7_0[1]}
   );
   gpc1_1 gpc2113 (
      {stage6_1[3]},
      {stage7_1[1]}
   );
   gpc1_1 gpc2114 (
      {stage6_12[1]},
      {stage7_12[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor_CLA486_16 compressor_CLA486_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb3afb6bb74ab01db81096e89b5d488629cfa742586907e4c25f8670c2fad9a0695ab0bb748ea53443deb7748f00303420598b244ce610587d9ca0006b54da5a48b91846836f0dd1dbfd40dfec682bd462680c3fea28d0984337467cea1c50915c1f574d4f3899c7e7e1abfc1cffd25cd583c5d0ae95acf117be735c4fbe47cef0fe8ad66a7fb0404de2fae1fe2f3fd0bf88b67a91a729c9c2dc5f22e789f529bb4d94503ef29981a4b17fa50272aa6b4de3585f5014d01b7a1ae765dc04b57d64a92e37404729be6a846285934f362c2aceb57d527aebac0e3d99d513beea85655c6ee2669db94824595ea1a00f84721bec82f5ab9d69b8e919dab8c09e22b567c1827a46fdf8c1c93555f785fc5ac5869369aa7b51f663d8f5df00d16507607d7e15e927f0840907ca560d762a79dd832b96c291aa77fb88271a7e435453ee5eb61088979b2c573128e86158855a0967b13db446ce167b8dc78f313abe06c9b020532ec7ec7fd570c1b4702135ed60692bd774caf0ca94eb494205ba22a048ff2a49bd6cf96f127c967e9a829bc7bb863a2f72b8401d900a00a069f476d4bca286d1357a40dc83a5b7722a27027db0733495089c1d6602418007fe3e4c938e0bc683b80cba418070c727d1e1477eae1cdfedecaee83690e1da94339ec0d8bf9ce533b3be48d553bd0e03d0fa8f069cb2adcde3e66e322d1426b6a1c287ff7da14cb2250e21f8968fa6ed3dc871c9171b3baec16e496e924be781f4d774570a8caa3d41fce32f46089c5cedc458de2dd22c02719d0b332b8616506dc5716e23eba62ae4ac7c5700bd4b4595d74594a5c71af3aea6e975bc2af359cd48f94c219a2644df48c128149ac2f220b30ff5def5867cf1989e61895936d2a276ec3dec79ac0e44a596903b28dc5723597dc373b21b9aeb8b1f84fc55ba3eaba28d3832318713d87bce101780f51305e222d88ad6a55e2eeb6af268f22edcf742bf7ed4dcecbaa17f006a5ab777bbcae2660613236c931bb3eebe9be6ce6dcc2cd148e845e6e13de6e40225d43341df4ee1e7ce30efaf47ed97b398d4d9251cdf39d0dbd1e82532df403fe7ac7c589c113eaa892abf7c590a6e334c978578fa84bbf79b1ecc60afeeb427da9a1c305ad67ead689769a439154282869df788d5d884f7e99a985a039e025b252391588738c74042fa294652ee49f76bd55c3a9a1c4f6bfd298b9f34fac0168d97bb032fbeb8d72d80913c78411c1a666381d9d6d49f20da5d108e1895c7d8852db1a572782a51a7b38f30730703782c7e1dcb943e33c5bb2b1e1261fea19ebc239647ddbb2292ddd3f5af9ab12db3fde2d7ab72349a0c4e4875241004bf819248e3f35a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h70165821eaec06dbcbf880979b4d916854724e5b7d6112f5dbf8372291577015ed4b4260769d34d198097b63f05a043fc1bfe05a8509dfd63b54ad97d74863795f0ccf3994e7086faa6fc35d7c4383436a64bb0dbfcede2fb6bc8488a4542f4f4685fd35354104ee3395123c318e8edc1d657c5f983aa98829e46eb040d66af7f2238f0bc30e92645935adb1bfcc600b300eed44a8ac230d47f729800c0d5666b4b9a11ca98c30357b1833348a813b74ce9d9f1e61004bf5cbca81b5286b7f0285fdc9d5eeee07e447d7c81d95657efcf4aea0117e2392d2a6563df0350870142aca7597aa99653c9f79252eb39eb4e208a1f27e359360b4228ccb8de1933f980432e25015586ed393c74f58681e6b71babbc6da1e88240b018dc4660ab283f1ab420bbfa3cde36ee5999a5fe68870ad706ac17af16e7d777602c91e91db81c502f5ce51fd417fcb69fc8125b8eeab03f8922a343efa4749e4bcd19b0aab8c555e2debffda528765cf70037238ac5e6fd84cdc9a95e9ec0276c8d9e2180c98202eacc7d86a0c77a291c506ea15947f16386219903c7c921381925f4de9f284608a601e79613008985af0073a04a5c240d0912b0bda1885687877266d93a4679cb9ff8b0eed407f45e484757c5de4b9932ce604babd6be119cdb13f5f3924a3ed3cf22a8bd2ca90e5624085540d6aae5858af216dd7c2be6f24c3a2778c102bcbb5bffec2f22b7f39ad5e9c88eb1c9d6fe88c36598abe863ff079ea98ecbb95884873e34fe590a873379ba4c4f7e8758a0d976c6f2a41961e4117de452b3d8241441113a45abd93b3082340b0db73078f2992c3adf46ae2e7f8ef2077963009f1b18b0c08d85c0e4949dc3f3a2f36a58a9cfad04114f79021f6b44502930bc985b7f367577208313801bd85b42a1964495c3b3e9facd761f3aaff293f08b80c563c5eb0f16409fd788928f8aee2c78947b9974556036189aeee0331d9ef04374acdf4f0521bc003c8e883b4ad854e778d9a6ea1775599d365ba0e0f1477190d688b1b596dc0af4825fa15b59b95180eb682f3008c06176cfb952a898d66c47eb5cab1e43c401261ecd3f15745af08268959bb59b123e1ab4623c0de4bb3104ed0d9ebcfcac9620c9be680da6a4a93c2b245284df0824a19737b4c5a9939a1642143c2afe7bc20faa33ffde91e3d41cf322423ecff40cc24d183a3a5b86a22417988bf86a1ca1040ce4adee5b7c2d33e1b6a70024679bc9d6b449cc7b8ebe1127e90e18608847f4cb6ca601244252b61c3640c631eab10169c86e54c25546f1a8a6da66b3c75dff362135ebd2507bbfb24d51e732d0707bbfdc653532321b2b30af7cbfdb0a026750ee4385871;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd72ce5db684b98b76f0c8781456a53256a1f613a9dbf3a39f90fd9c14d0439016a7d780ad31829d6efddee16b91e911f70d3f97ee34ca89b9aefff9506a3300efa8f1e4dc72d3e1957c39cbfc5f292dc78967576defbc079c2becc3da3ee4610cedbf88d7d6f3b94b519f6c48b6d5351f3853cae3ba1ed7f1c1e51c779ec82d94a49303b7f521e231b9dac9142b7002e6c3c4ecf26b7bd8dfe8dd7a4a704e7884c238a8a8663489efc9812cd841b662e064b4ab1a484392a3361a415ddd4b9c82ac1ab9b828da0429605ca8059b1c74cb552181ec3f3da5badf7f172a68e38cad387ada9b84989262a71adf782dcdd5d17de52170652f692337078d82ff3e86c42fc50c16be86e3e32c36f13f5992720b7e1b86dde2ca86ab765c6f240a059cc9a52004ecfb148acd5f58b0ac696fdceb2773ec8c206739b2232a6114deb1a7c4c2b4a414cd1b7d16c64853061484030ca9ecb0c2c2da4d632922ecf37eb58ca02e5da486e9e00ed4a57b2a7acace0a277a4fd0f5c900fc2d2a78a600b560e982cd737317bc1b9a6b474d4240a2ec0903330a9d6a69a7bc8011d8d04d8296889d7e52409cf29cad4a94f3f860eefb001662c77212cd44f09b58c62cea18d2963cfb04ce303be055d07b253cf678c6bb238aa4c849fb4b2c32a6c992e6ce7e1777c4c80055a937bf54251bcf21a19ee0e28591822e2dc19786f631d86da2788ebc21762b560bf0d488982cecfe95610b1978d88d0f8b518918296ee77f81930afc92cde86718c956dd92bf4a105b11b06e2c78ee68aaadff555631105e23b74afc070369e1265798f4c8f29ff35b917cfa48caf674bfd2f6ddd35b249d4b1925191e57c3f18815f601ea05ec9f7fc66862fe5d7698f965b10217a2c03e3ce9b1e32c3b4dc269a455ed639ec1863f8ad0bdeba7a8ca1ad39bc4e51f7ab473e1ac92449f10e137fdf655de3b37001bbd93a1cb9ca3d0ed5f3ffa9bd17d3ff61e95b49371b8ff36c19a6012e3198498420d49d4dec6c4414f7da9d2af1d608d6f78a0460ee5d856d2931f2d25bb935784ac036cce3ec372a51a69cca90a937d8e7d20e99a618ffd271c719ee765656ccf74bacd01be6ee19f5f3fb5b778d48006cddd72595f3a2bb4a57a073a6dcda2c00152a03223acd97c954297fe765f2320d81932b88f8a5793c5a48181f46767c25a3301405103a0b5b28ff18c7de55c80bcadec42e9988d2a14c8bb0d7da21de7630c1463c48f9c0d6c9fd6f1514960f4f72c3b55f08311628900bb28dc0331fc36205cf7d4d990375bd1e93bacd1e0b3d29e2f57a7ff97caade7b9dbaa5e3227d6080f549c4705b158afdc57f585d38dc68c43b324688fab7aac39a6bc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he940adaed4400fc764d2fdd199385564ec0516b69dfc31313ac61327065a596972469d7ab72af15d59178f2f9952655406a25c518ef24db803998ea862acaf8030c1fdde09380fdee7a195e00bae2a9bcf1bccc4d521567bbd374eb889e199fdd4f9694d06fe9df2d23e830f80543cb12a42e9f86559b6029f34d168079c0a56b4559ba53b618a64ccc73f805aec9afc479b53e8ed309d99ba0a6eacf41f8948a2ce1127eb036382a8dd8ac9231123a0a8a07dfe87a8b04a79a0984c20d442d0ec09e1baabea0682a71066a572b5af04f385a79377d28c89630248b53d1aabfeadf61a917d1fc8760af81f42b962801412268138053b42c27e00ff43d666c5a26654e539487026bd8d408c991b7d4dcfb29b381032f2cd1a373bc00791bd1424f15bea34bf0c49910bc29fb8cccc4c61b0fa381e43d040733c8c747a830c21d2df0fdbcf0421ff2b02772cd21a7bbec59429c58d25a7c2c73756425e328fd31ad3b0757e972a8a3cfe284eeadaec68451d8be5aba7ab4a67862e2dee0eb770ae377dafaf27d1df7421c4f1c8e716a605682508fea75755b8563d59397d390879f60e417d0b21fa02d27935dfe63bf90b1d2a81760fb485d97802122bdbd3cbffbf8dc5adf8177da1cd717da244cfc73b022e04fbf9245bd71b5fd8bbad90571e2bf1a05837a399b184ec0468de1bb7e7f7daf32e7398a37726f62611dc9f389a7f86ec6470e612f5280c76a4638ed512132714adcab4b24a579ddb8cadd69f08d83c474a999c9e8f008726830b19b27aa7ae37e599d7d575f8242f3f86ae7030a861dac54c6eb9c2329a4e158fcd7e6ccd41e3c81955772f10e1f4294b08cd921170daa92215af4e34e4b2771bcb48a3bd9485517f020f16c7127a5109b65d2b486a591cc43222688b570ecd309e673253dc1a1cd6c71790c95310390022eb6d0a698549e7d905821d75ec44f92c66a0945f3b99e699c580ec0a2076ce8b97dd228dada882474ff5b69ad5077cad902a3fc69bd03c20f38170e6e7d1e97f406b4d9f535ba20fff01a100f4ad1c6a17a88d0d7b0ea920271999d8bff3e3be1f4bc1af3b7519e33e09a29d04cc850d1895cade79ba2f8d2025a22a596c75219328922b3be8167a102d17a6f4caab658aca551c9c6bfd144832f01902adfafa867f953ca0987f15b64a01bc51a29ce21e98846d098016262afd30fb5a1de3b77f828b531bf7ac699093068ceae96a5fd2c3b5004d8840bdce0b61d10a578afbe91415d8b9e9b6eaedb48fcd768dbff9e25d09528aec45e825d1387d84801c086a49bd62d7fd097414a4b376c34c92d12b0f1762fa8eb87a4c7fa8a2c146f5cb30d2939d18c1b28e8ded2d173fec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb3ce826322d1253e91fc0950eb2324ec557e4a703a275c9330a0ceba447a4b490e74efebd82f53b88272c8f61db0b493386712b4b6a7bbff9d9f7a8efeef56a162b7c47aa53ce2333f9eb66d4691478ad2b41d997c328ded0a316f7b9205d4d13dfaae9106f0478d138ddd461939229d2cdcc5d66f75bfe9abdac2f038fbcd39eaed55c9b2c310f7973e09d42d838f1c688594b0ff9d3195487deefaef14b178834b2e389bfb1c583974cce5ea4fd9ca90ca5db71397b5de5d3886b1b0b67d3eae4f3415746f6cd2f581f243f29375c8b2da58b5ed29fe8048528e4c3d09f7eaa85e2737fb2dfff16b34104f4195a0d0c4911f6aeda102420b2a6b1fb468ec1731d4a0215545cdb060f5aeab6a63bd11199d442e6f12930d2cfbd45f7e4b3b16c1e09f006c55645b2b1b5dfe295e2d51cb79385d7197ce736cd3e0ba356eddd82dffc1af9d79cd9a82b5a178e9309803c3e77f6825c00cafaa3ee1598408da8cfc43692b03a23e65286b3669ebb6281278947a3ad6d2875bdb94542ddfc91ef7f810584a585e19bbebc67d2195a6fb6154c2f7c7299d9d34b5abacb4714339e7eecefec1ea553d7cee68c984afd6afd2e958f7c306e203b79a1a6fa6ce3272dd14e2125d7a4830087c8a001c71c8cd822873d6ab5743c5de2d1114e0c556bb22438f37d42cea37a5bf0b4a62121665fb62b7958c70ee11e34c70f3c14a6830600671b891e14a7e36bf72c47bf8a65a035d7c5cf079da56fa906cbfeec8ccb226dc1e9330a5e8ecd57d30ffe7b22a4c95b7dc7da10ab78d1d6f7006b9eaa50c45def7538d9281bb7411f0fb38910b9f76767539cecc31c9b81b55218683ce4fa99ed82f1a4cfe19beda4b7bfc6bf853e85d2ebff4af09eba58cd812e83d35145e12711d7335b1f7d86d1ac671d12be06957c83de1bf1119b0591e464de6a154dca94c48ada78f86d8accc0ad17cbba6cc77d407fbec3c449ef76db1d72dc8367d152db47a93fa730949e971e2654f7dd776ee4cdc89b2937c820f816fe30234c5c1ee6c29694f007bf3bcda2f7c1acbcc541b0b234b45ed540e2a31c2929c858be51cebc3db180ba660b054e6485a3a2958d392ba9c055faf6e4b36d39d34c3063708aab545ba0c2d4e085b7be7eb6af524b929d5c1a179dd3815e1f8ba2ac57fe484226867492926291e2e1d68990138450d7b199d17b025fa58ab51d7e848c0655dd0f7b4bb2b4fac94c28d824bcb7146506c8693a6bd6cf3c924647ab18caa9109a45f40c4fcb53448ce0c04343d494789d4eafd74c3c0e1e1e146d289ccb5cdf65495086b97e9ede3b44019d0755b4e35a078adf2fa358a0244e79697af7558432c10664572aae37d15ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb3a4f45750fa2ec5145b5eb1b0f07f2142c20886989e9437adab3b1acec9f8e7255f3d47cb67a33eef248143068bcca91fee2e79b3d46283c95a1023c54291b687e41f445982f6ebc8bd35041dfa4dd9a1704ea38bf05a6e3bcf0f31774ed63f9a008b5fda72b74038fdccc96e1f9e950c33cb2edc5b66d3039bd0e3eeccad7d0494f2998f577e48bb378a78e55834a213a351901f1aeabc7bc4938f4f0245e65ef133b852432408be8343fac0b646a7f51131a5a2cccdc1f119fe67eafba2a59904226ba2dc9f5e0c6182239a96cf1b19dc019eb48ee7f6396293d54b288bac395c8e1d90ca81205c5d4bd6078d20fa88c6e341653fef579fefb88fa1b4eef42f4930cc6a8fe9121401c8020c3d21733474c73fdcc50d9054aa981f95374eaeace2d0d90ffb8122e91d3f8fcc262ce7c8900b658364de345f77973edbe8ab969706f7d85c93e6bbcb9717820725eb70619559e38f368d304cd7d2b526c70a6c5f141ba9c93f2cf87d2aed943c4de52949cc5f6d904f5f0f9846b22218db469d552a6658215cee664afbba62b3798213cdce52ae6aafef5183a7e8f914bcac82feeb91bb6ebe3f2e65fcaf844cb4ecf474f89a2a2f7ad1e0b14cb90953d231eb283043ff071c62ec9cc338a93bdaff75ed12c0d3e8d5b3b04f0a8fd2c95737edca0f5f51f0f5c59bba04dc2f4fa9cacf6840d858f76a1f314659f455f770c96450c7d9645af88aa63455cabd36a6806d8b753c511c6eb25269fd4bc28886fd4cdb38d09526748755c8e86884777aed7eb209eb6b3b6488622a2484218e6c84fc36e665bf9f05bd260cc0efff045a51963efc14dc810c812f408c2d9bc1879e6a09852259baf9d0b8259e9945163880970fbd145bca2d45a58ec616346a7c4e8826666b231a90bab762de2ef86b7edfc37212c4beee9159e659b6a7261d43e661068e0d87232776167a4bd03a4eeac3fcf401837e38334c1840f67b5d2544ac4afa83737b45d3dcd3105b2416e4aed482bd60aa3667ce8c6e21f34fcbbcf74c9fe3f4d45c8b63b9374d4179c6a5e9803ef7c2c26cd4ec62a34560e05828ad0903620592b772f4740c01f61d02269c09efb38c86e158e5d15c9092a649bc04a69edcafe8b2470ed01ccc85cdfdadb3f6ae7f072908e0b872f3d195fbfbe2cf1eb42823ad6c5fdff61cfcbce6b40693297817951b13a4e131b22f4d7b0741c88f536e93ecba754737818dc9b6a4f6d086ed4b80b2eac9799b95a9b8de16f5fccf66e341a27b4da2c57e948f1e149e068b65f1104ef5c9d012413d6c2a5528555c17f2a434b4f4cdfd0a74fcf0bfe750933563e3c9d0a79b9c2c61f6ba7d955e6d84bb2f736d39f31710a9bbc949;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'haa273122b6543af148a68d27287091ef06991763de54768dbb3d0edee2863458caa64a8861eb8621ba0a6c9868ed590650a3a67965e6ae017a5e51de20b67557888f2f2fc309133939efbe84f156644bbe82a88a1e4d7884eab9367a87b52881fc8f5566a6ba411728f2dfb10536b13ee1105cd3d04f7b759c4572ef60bfe0255c49ef0c78836037c35fc2c7044f6a93dac4fd71e24a42a9958531e270230c202d9deb54daa45c0af4a54a0bcfce45d104edbff52cd4126d12164d1778ec76db09afea506c2b845f414916281ff32779fb48de93db4bc9d1306bc1eb4e5fe74e27c5dc5e2c78064116ceb90cb5f79698b77740fe93f17edda3d1982796d91e02344107cf44a0f95de43415706d382c3f42e4610f59657ea34b7a462e20f376d27af591a5e6005ed6fe2a0708916ccc9686daa3457ff625a6692616c6e9bf6c3224a64bf762e2dfca8b50b7a5080f976c0ccf9106960278b8bb26195096082176f22e2bde1e0fbfa93c2b1fed6dc8b9170351924cf7fb6fa6f7e270af11311be215c6b1611ae8bedd528113077c439a1efb2f59998abccc2cc99ea3ee7220451c6fb7d91d951cd41ab6c96194c1d41685e67c76bb4f136705b53625b7c0a25cf56501b6682f5625981fb0cf2e316136bb48ea09982a5fdd30a0f996d4ce4881507f61ffbe9d65474f40cf4ebb898e10497fd63bcb6592a4c7fc5f2c1621788e8b74fd1e51b82fa75abc213531f88dfa2252cdff635b7da3e0e36ddc60f152db8aa347747477613e05028959ea91fa77b2cd1178fdce64d75c70966342442dfaf96bad1ad51bef20bf197069b43f2f15d9b47021cd28ce8389a14647db2fc54f325ab5a17ff0306959c5aa7508599bacdba8644e7f1a73a05c8bc4f53a1b8cc718c837947a6f9e7d02a20554d57e79dadcb08a12d3fce82c538acb49876b333eedbf8aaedd255ccc67660cd3c14854361fb1540ee2c33a21d0ddf5de31246b54e718f66d0f39e5995d29b7f0122335ae13fc40d3ffa7400704b87a1a12408eb664403d653bf6c901aad793e97cebad5db2dd206aca493dada716f73b5f367b2a98af791929048badff877bceae00f7bb1898431ad7f997a758683c28fe75a65b56f85f6d1ee0552a7aaa70cc3d8091f2b837d612b374f12a21e6546438a4512f6cd901fe1a185128c6361063751f0a580649ba70bad0949fba97e085ef72073d1e7882ebbede8a0bdc1e3353889bd8ab8ddc58cae3b7476b776653a05c54e52408cf31d19893dc2c00044d5b6a325baaeb6f184c8d266a410f26fc1b0e38719491c80bb5753d7a72e3313554935131c081132fc9c71561ff1fcd2c6ea21618c106946369998393a496b84335e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h55d6826068e1dba104921068d5ceaf053313d6d218aa821dab34c68faffa8255a2a921c15515ba21caa1743d7a66c34766351f5cb11b261c746d32581c670eea4712ed5a3b9cc625d582e92394ab18359e4dd27d2c444855766447ebebc2d5b2785a75208ef07ecedb44b3b4b9ceebeb7a6b322ca5ea92d06417d6cc424e32e6d60cb99883756ce41843513c787d13f012bef4abb8e163a4c7ea03127e4952d8d361cf2ce70c4f649b0b57b88fc867845daa24c00a849f1749e6874ef16fc2292ea303e8953068abb4a7a0a0994dbf217449635f83141e460d97b02d10d5e910c26cefc415ec87125c9ee76f96e666992f13dd6a9b476c1d02393054b06491b7fe897b76e59aebc31f6cd34a68514fe805089d53a3d8c8dc46e05418597a7ef87802fd1ed1d65e4011a7ef425b3e7bee8428d6ad7a218bd5d4bb9bd38e59780cc519d7a90faa4494f72cca668b47c37787c85a62c7ea273eb368c3dbf76bcec92eecb024b614206344b4fe399a9b2038cdf3d58ac572dad436f80ee02e1b0450573280aac0fa5e5aab316411eb3d3a5dde587f16bc307655d64f79a0709e9e260fbdfa22df57ab214cd9632d11d008b14db6a68ae4275040a83cd55ef39fabe657e3ba58a9c8167e352442a96341ddcdbcbaf98a06d52109bda02b22c36071187a9a7b4f4eb875bd421a31cd36ac50060fff9b2e9249d93e1f9abe7e065c1f1989f76da1b372ca360c5b0a62788b747caff74a51dee9b8160ba31955ea90e9d01ae5bcd3cf073a2e517e92c879d8b5d88f3ea89dc6a07fdc86c915b0e16df33114ecb58ad01f20cbbed10fd98166e5898ba1b48b3696ae045b0b811343ea4c96218828a1e8cbf9bf331197f1c5113feac96d1b4a6eeb69c5ef155ecaf0312f6fd32be376b2047993de81a0f1281265592670106a4ffb01bee7d6d841c4d7774f9a79078b6c7764c11f8839ed7845eb616d94ec550157fb6199f4bb319138a208f33dda937dc6f5babdc3593f7698ce385eee6a0d3c2d86f0e7a93dd45c793156ce3cf6d1085d28c7871a8e75f1b579b2c20bf98705558de9aae5de6d051693848a8ae23422b38031d18306d8f6c6ae7b46bb826be8e3df674a72f5724799b041eb264749b97878e874f43d879128b7aa2a6c003ce5ab1a32279423bbed5f104bd6d5590ec9606458c9ffb13c04f411016eea764b0f574b08c7653952c72dd7e25056180cd6e19b749eb8bc8e9da16de4a21eafa54039e5e6d57a5a44022f8c774e7a504ac3984629d7deb8dabc56846640fb82f8947c7a13f49c084aaa5e71b957c572ac8b67038038622da944c95a8482407ff8d0fca6b8fb5be22338967771e54ef90b18a315589246c022;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha07fffcc6ac8821d9fc49b6e5733054f0be84a6f3c51f36e26032f6d642172865a054400a2c1c61cf4ff073016ec7358ae9a98d6449b08f92f85453bb1da789fcdbee467988b8234055287e35e4a671cc5d48c837ce649bf546e0637e4acc37e48738cafe3550e2600a0aa7dfade056a277a9c62f4bf1658aa9e2af2c8277fe2fc46394587cdceaf8a4cd00115fc70825b164ec992ed8c02b4f3b94aa6da51476ce44bb4e5cb4aca12e153c4fe43302153b5f51d38ba328a0a8e9f7700e6f40823b37c5182927161ff3a4f677245e1d2d4c6beb540f06f2d0c3701262a63cbb924a6afdd3a5f82e9a5b62f0514566fa989c35e8f5f42794cc184f40fdd1a71b840b188b9805eeb0883d65daf9011ceec3f17761c966d3642481d69eec17f0fd1bdd4bfab973ed55226105dcb145ed4b651e81eef895c6d024e7c1eb8f7208525a9fdb46d60cccad2e7f0cb576baa3723cfe3946e52789ffa2ce27ceb821293c4d1061be1fafecd05eeb0ebb0c4e63f6fe87dc8169c64c2389ed94ebd54152c30e1481954be6d81d4a6b543937a859223697078ddcc66fe65099320058ba8bb293b878e0f48902f3fab7af852fc37e7539e8ded15cfc0a0f36ccfe543858c4e7a87084e578b0f2f7d82d71cadc3b5650c34a3ac1fd51f3b97d3e71302bc7705fe562895a81282589b8fa7ec83570b443094ee596b01a1f2c7310d1f48a4d55b62e2f30677ed1be6ded9cbd3050cdcc2591498e7888f1c85375a11120e000036fb37ad9d1e8637db8c4b27a967c2182cb06d9963db65e5fc7f98cfb43f6015e9d26ba762f057363c3b918b47da1fa1b139653ffdf7a3d0f166942f9ff854655af4c72ec1fdec8348fd0dd3eaef6ef3b6efce530360b6025ba476627bee89df2b0388d501850539619ac021f828aba349034d5454f8e659889b056bb7f978d71cba1344648d3a113cdbd81bf473160e86ba4c00aa264490c363f396df5d563d21c7abc9423bd18c3078970054f084479204ac3b724e947bcf46edef4dd266be619eef70f3c9ba6f9c4be05df736cb3a9988f740719a9d7fd1a76f670c8f9d997405e679c8325d9170ee7612b6d3073f07a6d256f3914445f0f4e1ce6a1c7e82eb1b704b4b2dba11d6a945b2e1b48e8ed7eed4b65be99846a24e6a2038cadf6ce7690c76348ad5ada2fcede0af59aa1dad76476f55a6b1bbb35ccab350ef584e75b2d5c5ebac235194d7ab071ab06bb1fda2901ddd7d48fb154fcbb8bfe6e4325b346a76fd1c349f20be49528722af0ac8abf6d860acbd3b9baf44d6927461c0b9fba9b7127762dbd128c19a142007c1ee445b2c7936bede7b971e9dd83291a581f1f3ac038c0b46559b22d3c3f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h34d96c0c44535efcb9a360b391d69e83023d270f8034ef0687c0b902f6067794e7295e4ac98f46b0c719d34699ec7296599b99f900e5808efa4a89c7e75b5611caf72ca234c8e2cb59c90ba222c7b84b5b52454dff23ee29e7e4f52bc94783ee6a7c002d4350baf5dfc8bb555ae1074182046e9d052a73d05ea1f3ffb38dfc41eb5d012e9014661d37c2a42dce8dbc995b0649f034252b9916a7e43c0d14e664556f150e21ce2328ea2e22b9860c2b2d65ee8cb4be098e9d181d4869c7a29670a6ff0ab230972dc8a360869a1205a3ad4194a5111e8dc8e9d6323d00d2f725dbbf7eb3823efe4aed30c929f7eae08277768c59095ff05d4d4e6acb4c2acc7dfe707e59bcfc06e3fd8d3f0be2190a55f2bdff65bb6c9d0a3c67b0f02e0a470f96eaa5c6908a7cdfa229777e350cfab8fccaec5ebaf914773e6f41444d5d02cf6d283eccbfde1f2bff24acf43be6ff8f966057a132f5fb3d88747c44380aee1f79a1129a7db2e46552a87e3444f488f4189b6b1217f028842a076837df2a27fe81c85f92031a610c896e70e06591e094affdc841f51a23553fd0c3999f16658d7d4edb0874efa43e437f6586f85d67991301c9ed1b372bd109219f9c83f3190c6b2215610bd3a9282eca5a264b19cadfa445ba81f99476bbe97e508913eef6bfd671cb4b9717b1122a6244616e9d81c7c45aea16ddf5cbac0b184cc1f159e4b6e8210e9c157a6ff2798ea38bfd33bb014f13a676296751c0f8bd3153a501741c54d014182ade7dd92f1432b92b6aa9b72da1b155e4fe9e213abf82825a262a2d5ef5889002361d4a4e79d3d56bb98eea6019aa3121b0b89b3333e3989b6640f9273726d1c0181732ec7522c4129821bafdba59d11989d51ba1fe9970da4d89d2a350d575dbaf1f08f1b649ceac75e8f766c37fcc9515f12ee2f11e9ca16ad8c861c611c2b06ff9fc56821c1275252c9974e105770c87a5533ec25e26a1905ff92086daff3c0d6f4aa3673ad4c69179a6ae2462a2690aa8710838a27236f2521762adca772d3b015c8f54ab4dd29a5efb955dd388492fdd58667c90b35c2211d9aaec57960ead94cf2dbac810cb1b09b57bd1161a199002654f3102996b4f1582afc0993b911d4401bfdecb45ef3cf3417be1c8615ff43062757c91c7ee0e5f73a6c7e4131ae4e0199d3b8f3185616cec9c065fb3f70a04bd6a9beee12d88e6ec9b3b41ed49a3597cda7d8023a9a78ad2d2ac6ea1dfaa422ecd90a1bf719a985b1409e155046a3dba039afa0c777a7098187785caf09f9a092f303c51bd76f1cad35abcc7d1d8bc30da2ee1d5249e542f28177b191e91d6daa882826c24b61a793432371b53872c1f9c4567475f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3add3f56e40f97eae5cb2dca4dfa23178b77655131acfc0c994d631f9196dac810bbd15fb2a2ea99ef9af6e4f6a447d5359bc031dea5c52650f5365e3486561722a9e2f70940ca2c69b61c54352f7250329784ab192169b8d23f550100dd468a2d97753c93814125cdf6fda400532e0176634aac6d558bdd95a234f376d8845df29dc98c6f319b7a918428b23e7b7b476bb37d9377e014e91ff2ca65a2d8e97746acb271385e02e7c62144b120ee35b9de653133a16e879f23b372cc4da90cb8fa602077f6120883ce3399195b4dcd1c69610118ad2b8955d5012d335894756b31977de5563d2b4bd64453687c596429ceef8178a66d73ccaae5e99a9b6d801f7665ac42fc3a69e9b06daf012a82eed3d9ef15f557035025b04642993fd429287f04d456aba1353f724bae04c98ac22ef2a6287ab9155ca1d0b2ccb4a0429eeb9749db775afcf3350b56359a31cb56056ddc766b042d62d7bd9945b5858365006517a4283c5d87b0e9e391c512d52c612b14c2d6101e61665dbb5b7bf8fc01d19313d036c2aff7e336fe15152fa3b9e223cd482ddbfa5dbd396b14cab0bd6d161857e94006a61f0224fdb26444a01c30a87282d7e48735a2d68742ead4f65a60d48fde29d7c40d71e19fd18906d905b1d427cd30c899642dc6080595f07f6d889ac6296f9d3a9997051302ab52c80a434ca170395746145ded4e1df09dbc4b55641b2d3f2b6154e1bdffa3a400c1ee5911738642130cdaa748b0ea8f8f326190766b824ea9a90d3102b8b3d5db08fc4c9bbd471d076879e95c777879927b19ed1b4cdec929754e24ce2c6729862ae694bb4db4e4cf22aa95bf36606baa3c6dd3cb688fb71321da19d9b61331648ae2ce3b9e22f5c2d9f675d8b279aa2250fd70e7f16cf3efc3f3444f46a4a891f417798845932b76c194505d6319360a487e7958ec3efab6a9ed4b69134f7d24c915fc81ae86f1238c9902cacac6578b2d98a4d92970bbc9dbc7971a40d81bf984497e4642f5b38b12e7f840bdeac049d62a405c9c8dc040a2ba826dfebaf906a07691b97b6a86778ed6679d0b65f9b1f4215464ceb61eddf224bb7fbb78dd3daab099d9a2515fbd2a827a85c805ca104a50ba59a4934413c8bb47f4f0013988db886877dfc20dfdc57023dc1f7dbd5fd0064c0f50d2b5f3fd6465076222e8e601f3f8afd9c665c8f521ed4d75b32b0857487a160eb062a5f12aa8639393c31b47622692adc4d6becf4bd001f038ea892c7d96cb91922e565ecb4b2573ec18e78bfb31d76238b0921cfb6956a07ec379d328813794f48083bf91a3bcfabfa955899a2b5072d82f563e7bb2841f836142e9ab7c54e8d4d09aed5363cb8b89e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h72cc8e5cd7fce828dc62a8fa9fd15e2bd32797c427b624d3fb6ba11cca17789196b0862c531c2c6f436479d82ad3754f9e998e13830cc0c4e890aec78dd8cc8140f2ab70918288139b881a6511791d4586157e5efea580cee6c41d88d6df8a2d78e9e6cb04ad3fef7e42f686721a16e096a8a50c784f0f6127b776dc4b75b60efda958edd9204e5e7e0aa4ad84eedf5e7834312d91355d9ea4fd651ff333b894b15bf8f5eb4d8876081a1f221570cba6f2dc1e8c53442261b00f48339637b1894f31a2189ab7dcc6edf050e57a3612c6a3b2fa1256e71d896623f8ce1638e1cd0fd2c5dacd180c18a4f736a08754936471f04b61b9e3c8b09694d2928552a286af01b1402122ef40d51b569af84edf00a28b7c997a8a43301dfe05a8672b5fd2b9434b5e821395b4731ef5d507c05bcd828b7fd050ef116474f8d2c9c94cd250d58cb3cf388f662ae37fc6ae78d3938e0d831628097a549a3f308fef85be0441c1edf4fb70a344be3172ce903b4b5a06a4f6a5e8b7b823a209f1aacbd6a3e5a3838a3e9eef0b6a82a64e0d38388bbfbb8cd7049e580e429024a04db3829fd1d7ac52b8e0fc86405018cf5eb9622e655e08cba11382b24c26646dc7e3785ccfbbd92074b0875aa6880b287744c1bb9ece9d4ab8736e2b4565257ed5ff89a0842fbd84aeb190dc9edadce6090b0675bd39e97774d841658d2d8888895a3ce2a64324fc6a9898f3f362c1ccef0b0264d1408b7f704e04d1c36ef12be5ef5da2e3afb8df558c9e920a5332661ddee1e775d1fdd4a3badca516408027a3465371f5fc7cf9bc2d4d9d01f16299f41691c2172c7fe56b7e52b16a6b12a890d5416ed883dcc52b805d8ab100a5c781feb64f5546bb54ebd95c869bc9fbb8932c06119a16ff051915cbd33cc713951b9ea669fb831a2fede3ae8c7081dad0136124733a239a6708601efcbf643ed4d75b66702019f16964e62e40a444ffbed17d60eee0b3326c3c487c1e3e6854aa55f6d94cf39d8529d7930ed31a869b496e99f93020b5103b9e951d49f2b24fe34da02264f73f54e0d6d8a30fba633536807da503e164203c063625ad4fee638b20f16cd091b7847966d8a2fad39f18862e69adcb441cd39a24532288d5e851e291b98e78b3095e2f57de9d271a35ba71aa108aff30c31ff2481375f7b354df672cfc6a3ad3f8986a7ef93abf747830bd341fab90626dc6b6d16e6684c19c7634aa5a1ac44b10d14cac9b791aad7f94416484b9ab4cb9e6abe6c3d42ce3c1c0e25edceac89c7379c9ac069375891bc16eb9b0b8e8c9f0739328ea8f0e799546bfb509d4c4a181d9c46654dfd2c089f03a946de871b5a63042d98523bea5e2f4a09c8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h254316e474c83b76e6e897cb9534938a335077355fd0677772c6a934f3995c45294fd49e079386f00577104a2bc55d18321bce6928073307373c0a290dc42d570d7d2ebb3b76cfd74f30d2302dcc3d681f3bf22c41b44cc1931923f68426c94596b8b23012a0236466c7c94948e2728dea78a42b31fbbb5941afa47cf271af35a832983910bd8b56ea617f50d8aee6a8f315d5094142451fd084374a2fe4f27c499dd5b0d6a159b6940d4404a5efe85f0726025a45c210db8e46e5f850b7dea66fb38a9afcb27892fb644912bf098d61897cc8b75023b1994748e48472a2b41f7c3e195caad0dacea3931b3c1fd0f58cf08ae6c5c579cd24f1a50a6707bf9bb426b351e8e6a5d7a1164131b7d9e2ba53abd0340e7ed55761b4ed2156fe08e03f98f37150296c45c9f7b1c10a5f5a8695ed322a6fccf6f444df77d0ff5fe10e4508360642edcea352739613a468b3095bd90ef93c2e1b5726103238e7ebe2d89e99e94ecafc6ca4fe9bd601bee26b6a5a828e4c3ba09ed5e0e5d91681b0279bc8992ac25f6a0a0b0a0350391979b64b088f4f64aebd7d89f26026deacabfd8a5eb1e44a395ba9bf527ded3cd5ad4490a9462d2030a42fb0272ea21f997ea0114367c6e98ef690e11e9e23e2727a661cdd4744031742b174b66b6cd4591e08b051544d11144f781341998da19523e5f982f02df48c4db870214e2d063faebd0f425d0d1da2bf1f7df16aec561d72416d106d7fcea8da0f22ce87d29cb91813a988ac81ea641eb7b5aea06e7ab263db6ac9935b8c4714ce0caad83793ebe4bb55b64afcc0a1da7f4e0eea8a5a7d38abf3de178f31d3a6e28b0decd7165e17a8dfdadbb86921919df409d621ebd4c4ba40307c45a9d00c87895973e2939b862ea787438c4de437437363a86a190a03475c9849d9410d3211758aad9cfbc297294bc06992d7aa44ed1162be64c45917d5242b38e0948f9ab5bac5a86294432d7df6d97d231f6ab90bf8d1caebc73bac8bf65485392030b96d3071b8a47a692928d354110f5e5a7ed82fe63dc0e290da0bb620cf0a98b321dea6d93976b3cc8cc4a7c4cf538eee6995593864ba29e6f58f095f851d5eb9521945a9d4bee18ec337e01808fa68e4d7d7efa7da515ccdf4b1e03ec3fe7c676532c91c3ce02e3cd3244865bd323eed6db780bbd50de3ee421f5495fc1dac11946a357fcadc1b4a871175a8d30acc69036154c8bab6a02f76fe8652f91b397671053c588660f5edeb7d33241fcab64daa4fb5207a64ee3c88a9d38ddf67c6ed4069efdf9c33c3be0dd5e3728bda79472075e85fe99e839cb3ec55f475d3bf011442fecdd033d120c378a3e7c57e49b10360ce77b9065bf0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h930fa768fc4a591a02c8e3ec6120d60de55088eb5066fb930559587002476cf9bd1528c6aa4269e41207a80ef792ffa4d6cb745054bb06c8cd073c4f563143ca5e08b06318c4cfa3398af0e62bd00c6c65e67858934bff0f80371dfb385dcecfb694deb74e951688fdf41808aa0dddbcebd3fdc5e2d9bb8511966a221656f3d11697070e7d85d499cf379bcd78d092829c4c8de3e12c57ef0837ab182d8548452e401467d0f54743cce5b236befe5c6b1add606ad6228029592801ae8bb80729103b5ec8b8e0ca5063185ad5348a44d469d3c1637faf4296201da269c5997564db62911385c31323cbe4e4beef8b2de04c4837577fb9b2885912c591621d996c4f4a05ff9f6dfb640edefa8cff408f728292d1dc323de1093b01efc4a45960c2e908bbe74c03374e8808be293fbe1914b07b1dcd501226761b031a71850e646d4b30bc2fbcb1e31dfbc76f750b642c3cc15c6cc85d3d2c8593cc9d7b2344843f37cffac6842f34a87a77e0e9d8ca9b91407e23f7e5999ac9d93a3ceec304cb6f3c19b576ece55dc2b214bf2dc4d4228c624eacd742499c4747b1f0ca856810a2ddbf68a4682913e4a1169617fd50e171dc4404d1b26be79d91df99f459af4b2f76f4288afd213c433d44d95898d247f332334283c008b5647e67815659b4aec9f0af924ebb93d82e27bb345dd0d0ca8c9e7c9c26266811d06faefd417031c668a978e789e10971812b57a7bc7a3b7597cad2b183abd7934b207ab5d00d8d736debb182c53c037a444948d52e96954a44f884954af7247f6ae775ee0ecd1e732b138372ef2ff36d31a9ff42a7f48544c00dea3312c4210ba724d25f0c8d78b039e16f55449f67b8939e2724bfad9da47da0e997b3654e92a00fad8d21beb8202d8d7206c70272f9931d4adbc79fe23b9afb69b4c71e107414d09cc6f6faea7ad3a02a409c5ad58195e26946e20a898d19e63609cc3582ce0c07cb7fbe7665556861e78261ae2c9b32eb7046903c64c80f28266355ee31d4ef1e5b4a81f029e03925356e9a3255b3c80f8f9d03f80fe766abe585c4e013cd27779a01b7fcae2b3beacefae097a6716f79b9276f7357728998b5ef2341595bc73b460c67096e0fcf70770035f586dc05833b0f1ba51343939e962b2cba6fdc4f5ec07d2a15fea838190aff32a17b0fe043f089ff26d4f14b8d3aa80375f0915084bdcc56066015d0c4d410443ba4dd13509cdd9562be203f7e6a94f331c99ed3fa70fafd0a7743c742c269ba1852af131860a431d2b7ad1131384499cd17282fce6b4743d45c1508adc714bf10420c39a7ac487448ee64af4ceb9d1dcac4d2834a9beb75de739f17cf3ee20e1c5ecbf8612896d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h27a0e4123280bf112bdb525ee255e823e3bdc7b37565e9dd746a0a03e794d5591283352cd41e1d809ec32eed954591fedf2e83ad3b97e68c9ef5cbf2c0f7532b086893b10800d38875923450537bb3ace9a034bebfb781e2877984279dad1df69c8db6dc13a7ed3da5374f8e5afbafe6449a3952ea20137f343ca14503cc4b7b16a7f81c6bf708114029c94fe32b145e708cce82eea6ef7cc169854053cf6cf7410c53837ffca92a851e33e523f869653bbb7710bf7415b0cb62b60e5a6fab47f5483b737368bc239aa94f97753a19b149976543f752c89c6cb7a63c53cf68e23706a046643e261fcda8951bfcf16a33aba575b5925841abb6f72253b3ccfd22b951a75f73e9bfb2ebfe192eb73549888c3267c3665d24de0e7418abd785e982bdd54840e4c088e27447abfe441dce86bbe635eb332b5047c3dafc50939e761f768a7aa5875e396db2011c3c8af23089efc16ef7e5ade54359edc74b286da7667fbb915a93e66ca085212e1b78c70416c5e0bd7c15bcba03eb8bb21fe67513745f01f8ca13929e17fd55f34ec0728307c3e30c8b9b1ad2af8f1fc5cfac66c1038884720b6377a3c0a8225560d0abb3a7b8f7a674f2bffb5f1b69e5ba6c2d4cd3e228767107ad52c91f5161aa3e8f69e9f578801b3253a71720746fbd57c586dc1edf80bc50859e97a69fe8317995f05fcdbddd3ac1e55b3d4512e0ebbaba1d0c5eec8825259e58441591c9ff30bcd79c9e9763b4a873d87386ee74fbb297caec75f5d49bf2c7c3ef450aebf749bff3b3cf02189fdd1e742558ea1aeb46c0357cd788163067bc857b496bff356b1542f57390b4514b4ebcec2e808688610141ac6e00dec345e888df28634e414e80ef2ced8d530368a70b3944a6a43a42c19f0bbb3ce1d87054e0e6b2db7bb06721f62233884fd26b57bd9422f313cd8bd93c83a7f41fcc41cffff9a2b2b45b41b7c17da91fb54f8b213420d83e0556d1c0d24fabb1b7efb4446cca11cc927dbe45eece2bd959990a86152b3d3b6adf732c6481133cdaf53ef94ac12b6b7ee715c414175f59ff422752b49908ba800d598149fb611ba0e66da426d0dff0b2fb4cf7aef7193b2fdf40ffe9dc0a947110b01214ade537df95597ecc58997dfb3858e7524a3bf52517ac4a8db22e6671a5e424f12eb01881320085b78304bd000fd57eef86850e02b1ef8d8f6af08ba4b843eee068f8dc95f67032f09c39f67c2d23d77bde72be6923a9ae19e555fc7d174f3e84362134bf0e5130cf674d237e80b93f7a328b62653d874392da57532e957452d8b12a55d364cc800da853ed92276c95139f38816929221c76b5ae83ca2a7fc19a6f547d280b9e198a172b9d9ba4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h52f4975c1dd2b77c680cfa0c21cdc891933852203ebc1fccc4f67d2f5fe3971f9e0064d46309968bfbe43a953ea1a375f7f58b56c1ebb59dae06734f13c561fe48ffcab1a579607cda8a63f681716fb7ea6e50f305466c7e3a758734fadfefbb19322c9b18be739fad28f8381a7fdf5b9fa1858bca4a4d572f1d9a27518dff2af33ec004ff391f6a0b7bd93889f760f703829c6bb09f3f4e9704e5321c1cdaf00a2d61bf02c40165dd2fbb6798903e597d19b91f7a2bd864421a40b42e11e4ec3c07ae57925eafb41472d19379555a32163a24c8d52a2853b3db788f2e7602ade89a3444978eda5715fb4336b51c512970c50f7eeb3066fba6f64cd00aff9662909376a6c58ff920121ed176ff50b54e1973e88f794dd94c84b33885154127ad3735f9aa46a947752c53f522d89de6fc5b1cb763076c3bb539220a790c90d8803babf28f24473185dfe1a709c4ab2b2b61220830492e8c0337086fcffc8e46c8e760606f67aeb7a98d70345ba999e5b9c9eb0ddb2758e96f3d83b74579acc7f4421b2ac00bd08df7abc373f9e3a4256fc54f5944c1a05a3d32c160c195202d2bc6ee2d9bd16be00214cd5e4101b9bc39f1d7ba157f298a9abcc35789b13727871eca8a441ab77b0674d0963f32b1b9999d003fe755e09ab83d02cb6df803b4a3d43c71965fd3860ecf51183b69c4012024680dc75c69e74cdf35bc2861473530e06dbcfc45ff5bac931610e61fccabc8277b329972d2ed30db225f5f14054958937fded5c18e6bdde93a82d1d777d473abfc9005cb9d6843941f0568222d34feb27b67c369b0dcec34959b68a3004b6aa61135184dc8399386eb0719c5f6c76d48bd7855972d902e16cb70b62178aeb46c8ef8d4b6e0144ddb7c21e3319775ff230e6829923f13182d214c8ef4855ae9a5eac37cd5076e75b5b0ea80ad178c13119a751f1b0bc7f0bb7f56c903b0755fb8922a410611c94d696839711d35ca2cf6e0ab32acafd1a3590df0d0f6afe774016990aa8ddadaeb05cbbb7b071611faac0293b5a90bf6b0b7d91d82352f4728a372789e3f6b8b4ab61f5eb70f8c4b0e465cb1d6b834ada3e5a13ae3476c8c3c72be4ffff939a79146b351b593553c7ec171b0e9f85eaeaa762f0e50fbdb49ee1e39747a1a865995f38b2ad09dd3655e81b8cc77ac5a3af8b0166eea6b07951a8dfb7670f745b0b663a2e53d2404c7930fae9f0d95f18ba42a70cbb98f3bff8269a7197b4a59ab3e448ab511345c594f68c0c805c3ecfe644a760b4f03b5cc8753721c7c49709e41c9671a7ba746c55264219e223b67c9c58f8822fbaec26ff225eff172145b760a51b86b6952252bf7ff14bf8e026d0bfc5ec2312a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9bc0c5938e2b9fc50a046969557fa8bfdc27253df3fe5120860ec1e432a2ee05a3d61db3ac6dbd8830782129ce8e98738b25ebdf8807479e55c2176e03f16a8048a46bccd1b7e8ee891fab2b71961cd70368253ab3da5964bea013153cf6215927569a2b819285b0b15724cf818bee5274b4ef8e0cf95c4a5988dc1377f84d1f7dc3f7c17cda26e9cabc2e7ad92e7fe572c690f9f97dae51c7d594addb501a978234b25f09fc67418416f2b4b2e2b9b7fafe38f0970850bb59525c270e743552554c7daca027b68c0e0e3df8dedf2d159d4d83a331a7938cc793d8bd928b8dc6bcc969e37bb616a4e608736ef18a71aaed4abdf530ad69f713da35d499c7925a3850f43159ec3a2215c066fa10940ca2a7a4c52ca2f391bcc031817c4915b278483a8a510eaf45851a9348f76cff128821d8988f6aa7281c8ba46f7a272063d0e08520a3b4db494e20a787e49d9297e862a02f80b945bd4a378e061d7ce40cfde7b5e032f0c3a17f01673a97e59a39850a2e277a79a26fbbef406231ef6dac64d5cbc279a2d72e3679cca04ab60cd8dbd3c9de3833d43d169d8e305eac70273ca9460b2799037b7fbde3bea608e3009cbb9f6081e68981c549932ba4a58ff76dafb814e7d55c66bbd82b13b9a848b92c9f5dea14c6a12d9bc2c11a61ea3ea047796081d9d568955cbc03c954d6e3d7cf00ce1f78b56b2950b003d6311171ae776de795d70dabd33d4c617d9d8e86e705ba57c6a3bf0fce38d365ec1080d9630553cc264a6dec8698fcc92b330402d29c8fd375bf5adad28e773def4f8da8083edfc2e31bbc5894daa0e41f283c6ab7094505f11cbdb12911814c139e519254cfc42207eec863098e7c6dbf31867a9a5a261f3b330c9c958695c9033a53bb43b6158cce0ec9ef61ccdfd84717da5cb7a745389dbb4f0225630e25f626261b7b33c475c696daae0064422e41367324fb24c4474bc4c6ab199a80975dde05b4ed5c7c76d019ea04ea91cb106c4b090063d17f1722cd6690c7db5bb8de2234b13832aec27134601e123cb6434018f1b576a5a167e634855501fe2af9294a1145d223dbc78ad877949de90fa82b81312189883de3972fcc4a848d5b0acc0753a68a59c57283cfdc2296b22f758fc34106bef81d018b5d216c73faf4daf8427ae5bbd92f2841959c048c77dc669b7394bfbad9716d39506b7b15d0a239637ecf2445810343a493c48a2458600ffb778e6f708f048aeb8ed4c62b4177347ca138a3d63513056757d2d1269b883b55a5bc16c1616577805f3117c44fabf9088662fb9f328d6e9c3293e326e115fe16f4b110f2a5ceead4d851034eb2b4711caeaeefe4de551693b4f25e886d2164e36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h35c358e318f05157cb7d7bb853d08f0bbe959b25bda6465ceab5c6c21513496f6493dc603ed7ba9938754227502c2691710dfa6f9f93518ab92009032819e781b195f4f6b3448c3511ad99db3262db18c544cec4b06dbe09df99266c16b316593cb38c33683e121849c80cb170365a04c1762b2ccae5bed5723a9f3288073764d4646e7c5b72c6fab8d5dcb3a659839a4e031ffb8eabb023b3969eba403046d9dffa6cc2a919b2fdad02dcb7278bfcec08af4752b89dae0ac859c1a20fa48a50558598aa656f3c9a38e561b526a7c46be73f0c064bdaeb80d048d633824e1dfcc60ba335e7a0bfa24e42b198db1f4462357e15d979dd84ae6a60083b1e1514dd2e109c9684932e43572320cb15f807bb0f047b9c7df05ae4a85261e21f09e53239efa62d771666a5e895bbdd2e69e7308d76cbe4c28414466256de61ef9940ec7b4c3e673c4c2cead3d521ff0944661408592ceb8b7d779000b111febecf5cfc20e7f5962486bf0af7a09da1586f4c785cd36f013c674be66bc24191e9ffe8cff028a636d0c15b8f4b8c71c61a9eb41a8d1e27266f13721543b86051ce05fe5e68e45ccda5f57714c0da734500adfbe3872d21f589e27fe0362768437fa29e0529969832ee31db005e2c0a88daa035da566a73f2b1bc3a3619a20e200be47307701d1dd6503a64ef83677172caec527cc356e6c0831ac9681aea786381d88d5fbc0b438ac7210fc6e8408d0010b5ec804c5b6b3c18de406490de023d7f20871822e45637efa43abf75ecf886f478e3a6304f67b4156a18b2125e7d981304285adca5f677ff038867dc3309215925a568a98789e73b3396bda25e64fffe3b28660db430bbfc2b6ef0704bfab5a07ce487b7514f9073bfc42d7c439796a4af1ce830c97fb3f6a49cd5a787f8be991924bcd77fc6f9b4f14deba30b07bd9c54290aa5a2d7e7fc3713f4b831285da929853d63761b22fb1fc92b16c41dd9b3af1b4409ae9b583f725fed852ab04bbd786309f1230a41bfa449e76f233139ab5eecfcc9a13eabe462f9669ad6ee8dd74c00c078cb815a728e269f6d2edb08fe42116e8347f56cbc17414a7c38e56c4996f7428b447b4ac682737bb50f31fdb495ae7fa371d76664e8fe79a22276b0c50cba6fd52a4f9b98f27ce8395e72e1b52821d39cac3b39a5c30977eb6407705a309606dda3e4074642739d966c0e95b75bedd3338da95756ee68bbc5343695a1a4cd7aed22a8e64d8c5eccb5fd5ef8ad972f2437c9192d51bee5a515f4fdb65205ccc20b79a6537aca2eb7dea771418981b8be1907ff74a41ceee730ba199a691d0483e4e5229914faba9601faab6603f7886131f27c5df2e75b133d9ded05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h77b7c4203809f2a6a4567bb2fdd25e32f9acecb8648ddbd552bfe2260489280957e0f4f40481cb974dc690f95d675ded30b36e11788da9e1ae300944ad71617d81620e5e5172cb53e0639aaa9e1b74d0d697d71b772d9867deb58a3046291bbd37e97f4011aac87999ae9f521bd19d8f5fe70618122e2a339e18e1cb1610d0cf585fa730b0c4e7f7331a71b91f2105bf89a4c1e7a736407be3d94ddb6ff227f6ad7e270c9d77913fad93e704b506fb4fec243591cb6561da8c5e20fc84236909a607fb89460e913b8bad74dc2fded476ce44ddfe3b39c5f11f221ba47d5cdedb78cd5117b886092b544a1d6d91eca5d641c1d2f05bb3400478b461e829f23fbbf3eb933396b04f662a70fc303912270523ed5bccf0ca38bb00193f90ad2b44ff4bb19f0bbafe17fb98f9eda8c8d7f18a44e6ae7ac7c4ae29e559596862840ac46a290ce47512b0e1e8fd63685efd3fa5084909bff206f7fb4a3c6a1a18e5f18e11a4b1f8c9b68bbca733b5aee3dd14c64d40e0a6bf3692a47e9a2a2fc3c3e8d5444bcf421c8727c770f0c44a481ce66f4209b4268e694b18b797677966988598fd9b8addf15758784474f8875772fa76590c048c0e35730a1b7fee92f2bbd1448756fbd09bea96f8002fb6b976fb24431dfbf7e57859899479a0d92c4a74fae7e78f3d1cc95704e320ec9be3490a9d6730e04293b01b1e68a6235f1e920f3a8c3359a4ec79570db974c81cf0e460ed4c8afc796b1a3f7f9e275c983abb1d85544622dee01363e58e328bf8626533e31d4816e68d0e5fba112fbbc955f9bae9882c24789d655066327da3e688c17ab065a90e59d8dc9b069d49a5218c5627f0c5edc8db34e826a7cf2cc649ba3757bc53dd2bcc142950edd075a288b61aee075f4dfa28c35870fe20bc8eac3696962269685958fde45eae1e956d7ab908975c722e5cea427883a94c72a1d7aa77c73da5255f588bc339d196ccf82ce960b28ef7e654a72312b6bc5348ca06621f972d4eb3e61715ebc1b672ddf1f720dd9a0331472f8f6004fbcadfa8b93c5d429da48e09d62181321710d0347e344cd7eb953d415a39e2d393c1ebd7d48e566aa29bcf6dfbbed897cc67de073a46032046a9fb75ff573f0663b6b927b0799050074ee4b2b1898e98b51b4ce12c190ac15030d6ad3f6ae25ceb4b7372c0f31da85070641c0385d6771387b926cffee7f01a7d2c791c05a06b367a713fa58b81f2c64bcbc887364860084d31606b7eb2e7213937c246382f12e1559437597224700f360144c2d5f642ed33463841229f29f890b2db369429cc1babfaab2d621566a3252ec2bee3f438fa884047228106623791e119b1b6d1411f0a592a0867fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf8d9ec0967a131995e71909ed4f5984abf8bb153f2780d77741d1071878e5cc3215dc2d9712f5895122f8be00b4af439c253d4f24e8a2ae6b7e28ea65e2395bca5e0c4189e67756e7773b4a649c4ced9e5d0820a9f3fe33d2ab5d189fb4fc073dda2b3a435fa85f3983c35bf9bb667a004ad5a78d9ce4fd38d9cf0fef8e81fcac3e75d839493dad5858d808cc490527fd9515997a6136f3480851cde0818a09e39bd71fac02b116850858c1948d14eee42c16d6bf632cf39e896c53c906979f459e07a4f8e22a7b6e1d18b3ec4dcb466ab87d1621358eb8a5fc31320b06b7bfb0a7f2dc5d1f468df3f78c59abd9c0d30be6e27cd127769c63716a97b3eddb6b55a73355c418c89739593716a44a962b6a2562c3b5c11d62a28a5accccce060c2d0934be2728525242c4533304b534395d6ddedcf05874d0bd5a2681f51bc586210f01b7c7c37a356deaa62adb5bcb896e30d6928991c24a4784b371bac7e7c1fcb557cd8d107ee23808d802f8a2a2161d0cee29f88279255e350e5d89587b2191eeaffcd5c681260db0ad0113342a21b6fa40a86b8cacd0e2cb8a2fe2aa077413e05d743782d40beaf48a7da1392978a5854dca34e45975fd5eb2993888d5e03586fbf9680f0f10280f220f9c760adea61ae4dff7e3bb166f7f0c7edd9d0c58388bddf9d7e475488259a1b250f14e63eb721f6f0295bf579e4377d9ee44e58af6553c1469b6127d6c655c6d5baff9ffbe32c0ffbd4c4cd675a2cc7ba7ce453eb51e537be2a6c6b23f551e9da47f5f477200f23472de4391bbbc5fac8a6a9f0c4fcbcbb5686174cf9f693c6a83fb274b66728df7884b9a4f2f4676c1caf95baac1e830fea53e4727e718601d1a899c7b96634744f08fb93ef3084495085f3e9d1d105f6f1c2f8a7f8cefb28afbae0cdbb9f323e5c74d237be5e5f8d7d16ba05f1929710dc3a79cbf22e5156e9b24987fe248c68dc995d9de4c2c2b429d51899c1c0045e273aee23cb31d573dfff9e3cd0e543ecb2f6f8129a130941e3680557e9770a14cf278e9e04aad757106089e5aad7a98a058b05358d78ebbeb2bc88c3db7d4501620aa9841ddbf517f71c9a6504e4523365746e0ee1170438245b0ae036e1117eb9c18584df7c2809199bf1d650a4d2fb1a4d2b2ea6bc2d4c7ee1df5aeba2d2bb33f04bfe22a6598103d0257f9256f8aeb18e1497a80e9d802da13b98d959778e1a5c926e8316fe23945d8df33a618e2ce09eaa34d120f14c2c35f36a72430992b1f8f9a51adacbf8ecabbe70792b68555255c588394b582d46c6cc69ce96c7fe2c4562a5bc72d58d29e0688433123cf51d800cf7ff74ace18eb2d7a5f9be3e8ecbc0c4f1c596869b51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3ea735e5d595e1f15c25f21e30431a26e2ded77f96d10abeb1e0b822b1adbb21802a2fc9aaff256593ead0475f4874226a76ebde303c29ddbb59b96a28ea6ef45cbde6acf2d35a61ed692c4826757a5324871d15597ef5889ed9049d0d86e43127480d006f0781d1d5200888d34a4a3ac62760cd11908cfe481d0087bda18e0ec6a72976794c03d0478fc1a241c6c9435f3d9b04c9d254e40f9f63b923a689e696da84bb924017ceef76d2af5c42cfc1710815d30672eb7057e35fd096c6d64faa6ff1c98d2d5ced2b7c489ee312fb9b51795018bc0f2c3ab78fd03996f3a4635fb3a19e8838f1082c9c644bd32db9e22de6bb9998e5e0b1f9d5c49684b2ac93229a7d3ded85e27675a32a86e514af315efbf394dcb756bffb18376ab2da9dcfd4bb420e7c59d9da499405eab803dad2a6a23ac750253dfde341a5f5b95bf10bf708ecd56609bb380225518e8069ae206581d888321a671562ce4a8d41302dfde61df7c28ed8a0e6a47b2444fc1011154301014928758186b8437b8dc5e1fb8873c4f9d3506db66006ad4c8ec653f57c9d160d7f46218847a413a0117e9c9a00cc512ceb58808d3348d09590a387c2117d7f53e674952fe77d6aac5e07d489318838228bf37815b868b683c32557b86e77238118b649976a303061bf61d2bec71f9831d80f43426b46365619b41970eb5ffdccce836912f5da25042722932d1e0dc200dd0332a762b88f674f70841fbe1e32673f696d23638bce00737cba49bad48f07659017f4281d3c8190146db48e63ad6cc73e4efa7a7919a8eedb2314b50925a61d272bd89489d5614bea5f6c8a638d7c022816aa7ab060ada6d8cf379de3f414748b82814b7ec70d085673bba9b7b6ac4d5d1668ca41c552672ff605216b52dd4c446bd53811a70a89759999e13a28259c25189a006a59ede92901fcababb85f7fa02ab55d0bd00d935b102404e8e91f9c410e1c8dd828b1c1b1de3948bd8d76fb53632f5851d02190ab050ebfd1080a6b1edac8265ec7fbca49cb2be8fd53d7b25fd1497e2bc205a9d533b12955b9dc2644a9908ded7bf189ea1397095ab35b60224ea8f7257f58a4f89d4bfdacdf3b4e4a7c4e87b1b57275b1b649bb4811a7bd483d3a684507173a1e3ffcc2228f1cb6e2c4281b1c82bfd89b74f9d0549402320a1d86a48400f6f3fe08263b735ee141dd3ba6261f4d755e13af10830a232f05386226b2a2feeaf30d88dedaf4d1e0e540e88f279378007a3eb2cc75ceab9a48280fb84ff4e8ae9925f07770b6a113c149fe870a17190cd945e137d806c5a1b6a48bd572a5ac53bce8a9f2d3af5fad8ec419a388c413d604d937abd3ca4f6a4c6cf0589dbd198b3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6744c866f6da75b0034ee17c003d86250c57abf91356fe36e214eb58e3f5dbf1bda56c6cdc775447129b11258439add2378f53be0e6261a54b55f0f0a912480284cd112555084c2c6fa27b89897192a059e7dfa67db1e6aaf679e874a0d6cae0d0d64235d6aa204e0d25bdd5036eb9ccc342a03650f6d39c8174e05ecc6b67bab6d9745c61a39d3474b1da3464ba731e44db2af6a8b2c4a432bf7b5961b2688fa14942199ad617cd4f07f9d5a6a5eb057ed83ca186bc31eb813b241b2b6462ebda391a6998fcb91b8693bb0866159c37b24acb6e3f5a9644563f742d99a5ab2448b5af1ea6207f657703a4570fbd7f07914ca2022b1ea7d22d9a83da98a689126676a13f999997e7e6df03227e4fe61637875cc013e7b9915d9e88c2ee44d0474ee1956b462d9dff4bcd44a441ca3fbea8327e4a4b2786b78fe9df07e423375f5e3cb74c9dcb4a657815e404d24ad58ad2414fbeec23e6a1e7b5d25ed362dd899ec3aece425e8dd2a4077299022e27bf4f5d5fc36d42ce70f41a0b104fdc6cb357a838c424bcf215e768ded463e2e54672e551814986ec03209173236a257ba3cbbc031965b490f5fe982426a74e9e8f22ff9c574c13ca0be8c43e2bb2d400a3b2e1feb262e6ffaba3d35e066e22f23cca202d02e3b19bca2c645f00d4e9544883981f385c7ccedc5648892ac7b2747b2d3385cb679511df43715b79f502069a457138232218c20afe8cc3fa9b4333e15f80fff24748782b603038e4ae0b0f2c45f3d4105874a9266221eea8e95b1153fd8df99cd239da503715a36083773560f238c863803a10b8db8c5f0eed980df2c3b21ef04e0c967d27600e2c6a73b9560fab6f4e9e989e19ad22b3aa36ab77cfb27de05715eea323e07ab699a9fb17d5c22c9156b26e948869dab12d4412c86b75f95c174ac6a2247d0f0163a8a450ea722d5f3b44a36393a1b7c3837a60bcf4980e997e1af5ba352763dcc07f600d1b596fef08702f74ee256f2c1bbbeaa72171ca7013aabd657c4c6b1f4bfe6021147e745fdf1d315a29af15ef871bc57244e7b9c5b35d1e59e7dcb8cb8f12ad5848fe081364c3a491e9a5e0ab12c5a756422aa21e4ac4693344e8856378ecfd6baa592cb760a78c548f1f83aba02391b416c5138b9849e9533697cca7f1e0711b27cb8e0cf756f4df95aad7f8d23fb1b45437163434eba3a2b5652cc85952b37fea13c6c26b7c014e54aa639bdbf993b13876b4e1f2baecdfb4a12e263170db15243f9d1a0687e217dcc75f246edf3ce4464cf16ef089125e813f3fad561c41c361bf3e5945eb4491f484b35ae24d3169a8d385f1bf5233bfd70c85edc7fefbd5779fec5a82294fcf3f3c788ab8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h12050aee2489ac44533039c9a6d5602d036d7346b72a99b9aaf734799902856533db14ee0ef34df232fdeb305df3ef3ba781e428363220953f405d10793535785733ff9f1f5b1a8d79d13fee2b8848aa4861992e33f7115ab5e0183b1d45ce7b9d303efda32c715b9a4712a2c794f720509cecbcc352d52106b9f401b057b1fc2deb3c4d7fb8671556a2361a929c1b18d22474414a87b8af1d2f39d7faee862cd71bd86e38388310cd243d3835e1e5dabec8e6b5694a38e37e5e2da32870720aca11c29c84c08f6718d0b1c756da69bd1991fb2b0a0a6b4887197038a0a4e4a2a995b0b656f894c21ae5da85fe5d917354caa32683783e78245351bdfdf77ee2d1dba3351e14d38ffdc59e600262bebf6a6fac134f0f2d7942b258da619e0bfe7bd5ae6653745ec838ec2910ca57212ebbbe39c05cc4e5847feb2e4944c2cef5837f4dd744fc3b472b836fe4faffd717f5f9f6173a4c65f0dc72f688ff3fccf1b16a06b744b0630c2106376118c7cbbed016747f10cfd1d64d2d9f961c847fa5f0a18b45125b43cc270e39d2c22fe8c31714d36249282c21f6d26285b0acdf302dcc866ecfd0590b3f0eded3f60091a4e81e7e8a9c5bb373c4201ad66c0a2f2e2ab2cb9b604647e4286790cbee755aaa06472e0614f9d0de2cbbdca03de0f02b1e63eca07edc52512b60e71c4dbb4754a7359eb2d614f51c42641c468241e8a5a826c171528db7d81d242986207cd558fdc3d4b8b95899f28a43ab961fde9fb6270ad4e7b217f30a56164043752db6dcfb8fe0f403f28106963ac16f6d1fdc771adc29b6a47623de170093091c3d26f85dfbc3f8e407875e13a68fddb0c74c8d98afe86b27d853e71dfeb49e15f1cd1149465b9887a33c5ec1e3046a84913110af2f2c164a066d5e02a847cf17cfbf859ed688e595c988d3494d392350dbbc60c0a9687f93e33db59a1b50a0eaebfc99a793ab289b739e7be70d21648a659bcff237184f8c452b8816d9a1695a9b5e5af924f81b7e8d904206011dc069fb04350b876bd84c62a017a3e4da7cf7f5b6d1ae09d759c3717ff2d34e9fcadd38afb00b343ad397e76a42769b02d61de97e2020a825c7db09bc7884e6f06bad3913b0b7db09eaf343a6ded83ad71ae454a7b67f5e1bb022bef48e44d627196b3ba3c28f9e112053b092104ea75b9443931ad5fe1fcc9779baae0e7a7c77bb5284aa2d346bb757bd0db92bb3b034b3fe84adc5be7827c650cd606b88082fcb783219aa29745a365283bbaa1943b64284a5d1498d8fd8f38a92da0fa71577a5955bbf504aa75522e617be2ba7c60c71e2db595aec74d326adc3f498f7262c8f27b1a56394c12ff6432571d8bda8fc88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3d047b90ce5981f5f90f0a5b240bdd623aaff8a4da605bcdd9512dba9f26e1dfd419c928d0dd02252e4e417cb78486bf84428cfa199d447f66f0493ea1580bc1368d9dd587b8723ad154a75dc7b6eea6a0bd768fbce4e4357ee33ed19095e05e3154df522c01506b7a5ce274c7100b74319fdf6f07d2923644bbc48b9d22eed918af7bf339efe25f6fe95790ec1ae5dff06e0f6a5d180bccb00046abd7a61d8120a0140edfe7fee611739ae45ef32a1f6afeb43d76c167944e5d2acc385a26ff7cb5b14211eda984c23bc015858c705badc735b77df965120aaad7402fe9d7a4755caba7d64dd02f4caa0ac7e239d05d76dd365cdf61dc26cac787c7712f71c73ac1cbe7468001e9e8a3b0a2c24af93104c9ae12f8f1ec27b7853fba108ed74adc01aa6384a5b82bab0c2c4826f2c541b9319dcc37013393e1ee84f21b97cce9fea570f4ef4c3339c090ea29e042ef16e93e264c452cc737a103979a374ae5fa835f99d5f3375efb693a0ea457825a041d12a4b117a09de256101867cf0fb8382ce210eea9f9923f5fafe9d4f39baad194c6b89624664d731abc6649873297b92d832ac6505a41906391d511f6313aba7f16242da80416433acc17542f7fe4569ee9158bb1cc17808a9ebab73425779039a99e000c43072056ad1617ef3200b1171738d1cc76d8e7e1acfe0c0ae89fc377d6061148a237dbfa3bcb7775d213dbfb30490c08ebc2e05dc16d5a8a45534750767671a6a6177315966c19f8e67245c8bef9d793fde640f21f5567007e401abcdcf8ccf2c6d44f9b66088ffa756da5b2fde85ebe1c0bacc89684124a679419d68317a17617f4ad648aa371c4a65795e608ef83bcde59ef7564ca153c5737b89f6dc1f6b68dd867f28e4d9473895b2fb1ffa3977879de6ddeb22faeb64501c6c7e429aeeb49e3b87b0db8d56368e8961c0a06b80c91547cbb0e5f7fbf4408986908cafabe7c06dbe89525a425d747058c5758746727bd274cfa156a81e1f9b2be51b635adbd96c4e8ff5f7c1dd9b0ceb5a4afe49ac2e0b75ae964ed18cbdcfafe1f47d583a7d38898a7e0d245c6bc883a30518332b050f569614659a53a084f5c58a4a10492eab9a048d90cefd3bf0b1e6cc755f1ef387b5b2b52f4dfa06b857b37f657f2eb40fb1d73b298dca2d43f6b6eec4d38e18934d5748b024aecbc02cbc42e6d8a44edc06e578cf5250916b8e575092f2f139340ba5b50475f0082569f1b0538ac5b0d404c7c204d2deeda93715eaddac57a713814465f0b7bb043d7b32eb15364b0cc7df68558cd603e36b393de62534c6ea60d6ec7a8160c0a92577008d97f0932c18391acc0c6e2ae65734583670d1abe7541590c1a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h76a3e128f237c0c41f485f3a30b5c6d3eb0eb1e27854362a9fbf7b5f756f2f37581de2e03264d224db58b56ecd42be57d5d47117d7d7c1f0cac89a856e2622e01c3d22cdaba24fcc26904e83487021a48c04ba78fab3bd683d88faec1f3769b369b7db16d67b40f2736e50dc552e6a5e5470af12058114160677632ce4c7c981d3974f77a83b6e63158ebcf1fac9ed112dee995e1accee763fb4aace889454e92c54da79f1693ec267c4844bc71bc0eeef9bb133e0f7a2a409a65dacd6d6db866f6271eda9c721702a5ec012468a142f461030ff10c3e4e366325e536186ca4e0bb93d97a440e01453fbbb724d43344a6d4dd0a4284f46042cbec15011f52e88456e222a4f34376c8e543dcd5c8b8da1aa38bc0cd8a25037b82af3fc64d77b346557cc5f9173f790773e74a3021614451a7c2d4a93de7fc1338b626d798100a5c54ba5ccc7b50897e0c6f601cf0516865e47e339d776bb037b62709c7bc9d03a95775f71f53a1c6d477606019462c0b0910dc8bcf3d2ba0434748f248f11a6753effb79c1a499562b5b982fe225a53f61ec8c734eb504e8054aeaaf1ae4a554c9278a0d295b197563f326c6e38904752060bd528ffb9f583e9c412726280fc20fc86100b7de926f8b7eeebceace5d474a86de6b70c007b515036582f8c0e230c8278dc979298a8d2ebb19bea28b2cea15b33221c8445226db0c0fb8aec622bbf81522bd27ac224bc62877a7d4cd568c1ca2bc8409efe50f0efbfad171eef2dce3f24dc7cbc012922fdbbab083bc89e55b433168b2ce467bbcffe820e76cf29606001c8bbc2f32369d855ed5c87f9256e1c85588dd97e1cd59b12d0dc36fa426a344a50ca5bba9a1a3768d4d379be8ad2a9ebeae3ed2d84ceb57175416e6ca128436602fa7587dbd1290d0d0174e94b41054fc6dd174ca1aa8d486bf6ea91e94318b6e2328ff2cdf446fdc918b70c35e93268504d08805dda5fac4837c6e852a3c08409df2bcbdb958fd62546ff38f9951496bac2ffdd6492fd1294a169137ece6ef73316eb00b978ebbfd8255c532331063acd117ecef219b652c102d8a99692bc53aa3659b681ccee6e220811d4d440589ef61ad863bebdbdd00a05f92211d0af47de3008ebd118a52ae2f38166b5f75271f39292e171638d85ac03abd891d795f581b49fc7e89dbd85945cfd95e2e611197a435bf111f5158d0f165072d2cd1568d6f22a0118f84bf47bfae90b71c58ad724f8772c4b8e5f3e5e4b72da8c131754123ea5dc955b8837966edb6163719611de1f9f0f0465cec87766d740fbb31774e729b3924c29faea66e65d2e4c34bb8752d54589877bddc2e1532ca782706de324be3d3c4d973dc5ebcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5b569f6fe40740825722bc892670740aaf3a6ebda681f57199574e08941ad1b6d6d82720845a1de10e6891361731153bbe2bcdf2edc304aa74bafa02aa1f9cb6322d663feaa4609c56d349bb25770ad5be7bee356879dacc24f2adc422420fc77290d832d2d7b795deb05ac798a9e212a8b746d088fd1a268fa9c14026f1da61465f29c89f399ddd6bf285c8014040351fba3e29a7740bcd4521aea59eb3b69a913d347a0ae30e952acc65910e5133730d72e880e8dc40683c22275356dada4a9bc48c3a65906553b4375dde565b83e43e0b21f30ec8a4f69f0443e131210c0d8f353daa87a16e34e5eb27ca204811d0aeea10dccd766ed88e4cb8c280411dba76a2eaff516cef264f2ff95cbaec457aaf889df51dc29e4b079e1624a1ae2784b1f37e31c43da14803f65496183db4a2a9a76932f38e41c873e5c2b5622ca37426a8c5c66dd0943d5bbb4da8a2dec19c169c8289d174f8d5c7e4bfe414fb84cd39b0d60f573fbf8dff1093164aea3377ebfc561cca0d0068a25f6f9787fc8ef197ce840f31b0a09571fcd66ba496d66e6cdfd7a626a48b95a543ac49aaf0ff002209e94281da5052e8c49892d11dfed5e44ac3a07e5b4cd034688c7095115d317b2b4dcd3c35c1cdcd4e801b16521110b69f92fa1da8be8658141eb6dd816d77849c0edce48337e0b7f6c5b2eeaf62133fda9bd7482f5e514adce561ea61cbc319faf7360c050d40dba8b356b312cf46c1216910b0636c7b592be8d261f68fa0f0d9f0fe9dea2edf1f1e07b8d968a5c89b688d5d8b45afd39ce4aed2b366793a1b335534e138efb1e5bceff3869e39aa2c8f74fdc857c665f698979a39d3f6d844ca0ea4699d6e7799310ed016cb02f6cab01d337217c44faf4995f68fdb62ba13ba770dfe062acfff5c88669d4d1bbede53f0a44f3b708f39fa3f8d7e3f4080ebab576c1039f93c16a01c88851b7e17dc81237928fb4331033088c51a9bfbd2ed9cfb6251184da9546a7d5fc334fde66ad2eed01afbdc8984173c81c64568911b83844162887a98871b6aa660f2b1ff95981f62aaf07e34cccd010c8369090ae9345b69dcfaa2f7c79c0aba43d32b277ff6978c7d0b5c34c4b0b3fa0f5b30c20eaf17a513e1a2dd48b7f2a5e242136d36c17e9133a3b2b7a80ce5db4142aaeef0123c2b3bd5b3555b35482dd8814eb19e170fc69ced8fbb65b3f558e2791c0deee9a47f49a3ccf3ebd6b1485ef8f1b260dbe2aea6a8f8d5e9826e16b571835b5bc57ef2442a409525bac63e3821fa819c807a39cf621108d2449ab40e00d2293decdae0add080a16cf63e7c94cc6c45b30ef4a979238507eeae63f1bde36b4882aad9a62d680cfa7a22d7b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he703357da4e0736fd431e798514b06e7d31a07d677120ae85397691d37af682df0cc63fc93695ac81b7b9fc7b94bf3f0c508705b18f20efb090a2d8e62760b4d70d6b5ee3558f6d1d67997dfd6e80b55df06ac5a01f7020d64eed25eda81e5d3e04c90d4a75346196584b261ef865d37c65043f3a8e09d715bce1511025b038f3c663f2b335380329b7c55ca5a71b2d96888b372006e843b2374157f43fc0b6ffcbe0411a76b6da84637fc431485b31375a11300a0801ed3f02f1006d6a99d1443e4826290ab45418c7382cb5776889cb24a128b16c2c1f46d741e0fe784d959fbefd06b8b966a438df8ccd15292a750bfc1c844b8fb5eefd2d22100a22fc797516e4e466ae3d213d2b58ef0ecf998a986b3a54b5c46379f9b57c6b9f8bf3b73955d25cfb1e5027e3da848845a7945a25d7a445237a5e41337ae3a55af65727d692cf9aa22fbd5372a903e2d7ea1648adbb56310da6a57fba76faaefea10bfeb3e4f5e5e390fddcc8280172b65018fe5c3e14c2f027c81d902d26bab0160d11b39553454762303da0946f78dbab190cb8a3ae0430460be07e6035cac53f23aad7a4e99f1f4fc7b7e2d789d7e6964dd6816405c37c3c2d24c684b2bebe45efabbf6a452efcba9edf135927b77edb16d0b1e24d1b21c7e365851143a9c9938011f0a544f39538cdd434d92c12248a6eb625464cb4b213bf039cedeac453dd75c81614f9bea690b78e71ffe599ba36eac1135846ed85c06df1c12d5b5b60411ecb4acfcbe0f747c52324f2da44a04e6009cd5b63c3f1dcfa48d105d4967d723e9f32a55b2b48a3c122ed6b09980521838072b76e5ebdfc7f5c1e5fe5ccf982f513d6ceda655d7436e0d4bf87a6360003cd2bbec6868ba20116330b14aaa8fa2fa4e990326365863d161f8ceedf3cccdbf5bad46f8d67839fcffa972229c8157f8837d862e2403747b298ebc14c0e2dfedd52623b45aeb4f65df7a7756fd6ac22ea20d5cf9c54626011b91c876ecc8591a51c7a33b4727d19ff898bbe3a716813761294b23fe62b0c4d33e294ce3430422284f50725c80495fed89b0845bcc3aaba6f1756ea2a39dba94a6c72b1dea441e2f99fa366b925a6d3caa82021fe490ac2d52e17baedd653ae69a96f575be3205828ddf3a2672f1223edb18162858aca4d09f2bff0d4554d70dbe68460700088bab92766803ca7ecc4e39a574d4e18540d04f6f3f4ffdf476c8ffe07fe2bfe8e4995f2d4283b1a99b62bbee8495579374b4af3f11ec1e7f490b1e26a3ab81eae720b819777cbb6fb1dd6e86e1a2d9f2282515e506566657e26c569f6c54ae10d3330fc37d5706b2ae8a330f4a6643dc7ca8a952e8fcd40a29bfad8ab5e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4b55b28d0066965579a8fd7790c788f41eab7d7f4351430050d3a444b4beee45c3fadc80f0a9596502c1a41849d08a24795dd2fcd01d86498f287656679a54d457860f49cc72dc45492fb14024aa33aac133477aa6e954aba6d3a8d2bb1318704e1d58f5530bac360c0dec3e788404be753c493d4448074bac3ae558afe0104df49886effbc8525daec84aa3db78a156767776ca4775453056f18b3f3163c799e080ac9ee8198a4a83960414ac998e0b8086f15b5213ac3c2f9ba8d8b28f4e1bb4ccabacbd82cec1a2162ebc01ced5b2059221d6ece8c1be394ec771bcd1f522b72ea393422a9b9b7f77338e79f7e99eb57d50d7bcfc8754a036f70ecce91829247d48940737c7bce9256580bdcf50857ff11ca34b2d4bbff13090c61637f92e4bce6f708992fac407f7c0e840e5758afe9408498abc5f2860026a5eb441eb1170e0108a84e0ed1631ed21993c78bcaa03b5e3faa2664704ef9d4fde626c13d5054c244ed3acf5f2efa8c1bc6a59f79c32ff145604f2e4b6678bf03fd5c28d770cab09d5d4cd305880db36cdb3a8aad5cdd9e36ddb881abdc70711e931f340fd84f552bacc05d216ec4c16a62a7c4ce8250a455c71039d83201aa0084cf15cc315a05a296a93ab9596ea1489bcfd8ec406af3cdde323d6ce87aa9d4ea22e2df10207bb6b76ef77e51c747f78ae9487130b48e7f20179c1a3a097cac3fb7e55a8525d36ff22de1aade7d13206627700f28645019d5fb65354f82a53944c0e73af4258d9db25273a92f27b983b3d91d1be9c5cb7bb5e0bb576e5d938c8cc80ae48f77e775961ee03a81b22a42cb7f220674ad213654290030eb1739e5e2fe1c5eab9c7973b225548027dca8df993e2b394af9be5f45d165bb27440ad358bbac3379e7df954f6c62ee8c1e6d7338222b6b43c0e47a9a0bf71ea76300d52682209a95feec9e5cc53ca49434b248d087f862336c50a7f0ec79e00892ec81725666a1d20eeb43dfa2d957f5aeb24d702e188599b6621cfba36656c69c9d4296041022513400c102d063a2081710dfd7c7dd6565c19171253db035bdf0a8a6354e67433a8d0d73aa273d819010983dddf9ad27f967f44a8c2116edab033aae8b46d8a7b6ecabd9c4cc7142c95d678bf32017920fb911a0aa62265feb208cc087179da63e993ada9978c9514b4eaf357c7d295940c31206c906961a662b9b55f6f3fbfa8c85066d40795ea63f40e1dd643550e7927bda29bba142adea4e9c0d8b380d0e3153c9cf6e3d34addfd9bdcc83c9bbb6bfb873d83d9c1e49aa18d61d2192aec59b77c95b2c6327f487ea231f969c354016bb45de30cffab9a3bb10e84dbb06615dc4d924b492e058dcc86e544;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h598547db73d853de74f414c9625adb7550c0245e1b84caaa1d328ba23dbe4580c2bf3b81ae42932f4155069bcec202557fd17b311add9c1a1e2135f9451b1c3fd8a0c135d28a089abedd88ffe126185352548737d45a48c36d935bf3e0a02d7036de9873fad37e3e97fdac1fe391ac062d80b8259c81af78257a7540c347356b9decd65c078bcdbf2e15e86a8fadcc1111abdd131e2cefca723cea98d7da6953c63a8d24680ce2950f95547329beacc68288b44a929d548240362996fadf9bc94e5c5db34bd044011e9242bae87fd6299d899416cc5af0c9870105e0dd4dd552ecf18d95a1eaa37ddea979a663cd84a041d6c2ef228088c4d3879826090841724e28ab2ede976b74d6f82c08733cf6f3eb8643cb0a13bde623361af82a1339fb3f52d93d702ad2aed9fbc27c1d04e6b86dbe24b1b42a1d65917f2e32b8c9a578696f703c11f487dbed6f86c36739f359c7e56a4e9206becb0506c78cf6e52421e733de256a6f267d7ba343146665e8b4cfab0e57c41e42f8ffb4f416b5ca0b28c13cf49f2e58bf361a25aac16f424a6b08282081b765f3945ae80f52c6b57229a9accb79cbc30d742612c15ec369657fc71b6c1f300e7e948168593a5bf8ad820fda3a462e429d6ee71d1b509f0a0759979a90504fec9878c5c7f29668f3c48115c7079d723c261b8390a3ad2b5cf728536ca31308a78f87b0ca23173109b7743c85d8e60570898bfb5544f88154ca5cb393e09965a53ba123bf80d4626c6c48a26d2c1fc5998aec6c75681cb68af3aa5d78366c7e6fdb02a6ed5ee962e41ed0a115b90f8952578ca61cf983782cc956f39d7b1e0eea485e908e35c42db7dcdfefdfe82d00b2e11105c733b75f710425e11093524017bacea9bbd723466a69b96e96476e9e4d2fe88f1a70c6500c6ec854d1c5090c089776328ffe606d9d3b74055101dcdcc295853f495437d1a1673e05bf74311db34d2427aef92cc4ed5e7e225a509e6cc7d0cdacb21bb13ece9a3203a325083418b75ab31aa2690a307f03b8017f5fa152aacbc81d7435e84c3060cff644f230e8ba179a3496a8f3dc462940b86fa9dcc2144aaf24cdf0c797249ebc44d91b38b77eb8f0ba577b911d96f2be5aaafc7b522f5aa43de6f14f71c108cb3d2a16bede866a3b9fb21e4df3ad02c357e9d6621290ea5ebdf7fe13c4b025822bf848cd10ae59d30493bab1a72ad4ccecf60b2f8c538240433adb8784be1e00d6c9e37bac44193cb30a82a0d62249306d600b41746503bbc1be230144e6fb85a7661a65ba8184912590a69e231502ce47424385e67194bcfceb3559a6ae930764fc93713dc1d6022c27c2e4e52b5885cd6021b74300ea411cbb32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h29e4cf67ef4dd463087a12e5e47c9f5739fa86b7fab403128fc864f6e5b3fa7901866113b56d5230fb1a2c6532d8024f461bbecd8c9ac87e8ff3b8216228afe22c4d5ef761a240398d2c0b10a276114c1f1f239424f9abff3f3b4f30af2e75f51c73f271dfde6835a593721ea7beee40d5f9ac8c7466952cdcd2b472f19c2efd3fbf878067441335b9306e391386fa1784050a5cd98c678010362a8c4cc6f622e495ecb4563d98792c1b16962c29bd0c7912f7e174dd493e8951d9d1ac7fd2d360d218202b4e134b728c28e82122a49c83589809301a1dbc1e9a0fcc873b7b59fa8f7ae112536a680096f5e07d67925d7a5e53bd23ea1fcbebab968162b5ec3e1a325ce3f751422cbd34cc39ead99bc0d11da152333117f3ead638b7e79091df5a812984fb125a2a207a16db0b2c326aa42462dced289baa3e9b0822fbaabb072e54fb435f082101077f85187bcca856c1f7848418933acd025d315a9ec845ac754662543e9bc954edb61a7d4ce4795b0dc5f71de430f2480d837e006691c05785ab1c397767628d1ba4c8a84660b1bb5504eeaa772d75ee7459f742fc8edd2362af45cf9dc189d0cd5623121c165bafbe4b83f7077b23e8d62f63c25a297c7a7a34a70dc28e5a1658a599657aa56d56d3c00a073fc18c90b9c8fd802f00555e7e3b6b1e2274440aed8911727595fe8db6ed936ae4baf9877914ccaaaa16519b25febde272eb5196d2c50e488d7c894fdb7576bc125bee7bbd053b5879aed299f797463b77be78e42a7578a5ec108835ef3f7b8f5f8253c4e3ff84e893ea24b778136953a3a12b7f1c292b0038a87d980ba856474b94b04bcd313cb2bc364c73314f5746ac7497b8d1407ad45dbab08fcb3cce9d015776aa2cd5f160b661b6aa628d5ccec57163fc0ced56f9686f99aa050d4ec2996fcff4834912ec3aec8a966a2a7176aa79e40b026dcb3bed851bd17fa497b5ecef83468baeb1b6a0d1ae4aba168008d79bf40344ed92aefaa355c077ec6e396100e8fb0df9f51da2578d6cb0df918f4d71225bdad5edb7b1755f0fa797e89b4dec66168f85488ee134bd2e5da2a0304f37e2e8b5d7038716a495000d4765844270803ebbcb41657086c0b64802d6857b685d575bf296ac2e0b9c8d7fdc8ebab83350b749d0c7bc862e787277def1cd1888b776a4c134b269cffb8690f955b9092a559cbcdcfa653b8a2bab05d02086b983c2998d9ee8d374c491ff038e2a9062581bc5ac5492dee11a5fe9a50f451893c4ddba1c7dee4bb13112b2394242a252ecb905fd4640d90c9a31a210dbb0d9daf442fc2b0ef3b66ee441bf8f87c4afca176eca30e76bc2bebf4b439f68333e8bb2308a5186f23a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h2276f37732960cafff18dfd8caba6920eb6a75f881663f54ca09945d426a808a1fbd090513ae15ec0e5ebd9a6a3ba2077cc70f92c0f8cf8d9aa76d4bf237e373dad98212c39c3b48a8bf6494bd03d5dc3a9e7ec7d5669144e0292260eaa57d744aefb353e99435a578350aa5f271ec17de0cf061a5585797bf6a92fb8fce972336ae43626701fd3d73d772d81e2c8f02a22ab1d1d55d1e420a5d1a9d1deb484d5b07c11b3ba08516b692074d6af062bb22ba9966cb54d201c2560e7d49e1b8e1a2769456ea57072d1f3e70e978d2b37c3ec83506a50387eaf4991fd7046d87158e4a45f83334e0544a489f9390ab8953bb53b76087037667c94d916c3452d44fa1e0260f7d9c13dce926078fba4759f381674abc28a48c658b91acbd9a1cff4684f7c978be39e8aadeb8a2880e3ae1ba7581a98460d2c0804522842b190a02bcbd425ffab509a2b4c1bc1c7ce9f5744b43e22943059a1f075987c3701eb5cbee7a0b35d0fe6e2c50e5cb7685cb13aa34f39b0ca8fa01c17393f7f3a2009190277e2b1186ec946819391b199378f570e02d83987ea32a0023e7aa969265264b3d82079f6a3906da3a0c31bba5381c0f08fe11370ab9f4cb05bdc68ba16151c987d1f301f78615c82823c721408fe6924fefd372292f0fe976eacb03085a8a4611c1d1468f33e927f5d3a45e5fbec54fc7100da25551a97388182fe36805fe01dba0765660b64eb5425f1416da689130e3e7f914ada5362c5813480777e0b38267fc0f4625305d852cdc8d7ed171e30de7f4ca3087137aab5cfbd02d330c4f79cb8e86d3c2d5851100efd732b98e2192f3b122a14a22ba3e1aa81a9920e135375631f99b985754c9369f6e06cb491fed3b5905ff06080a6c501ec0a0e7df63ecc02d22f09e96f2d65106c6e34055a9a370192ea4b94e4f4163920d7727cee14f096d395790c1602680f315d95252d748db2b22c0b1b333a5cc1c351e93984168572e573df0d403d031df0d371b6474bdcc2024ba8e39a3e79420f1afc15dd30a82147aad8fab022b534d2a2961edde99e8cb838775b14ffdb5474c81fd2810f6dc608dbb9faf9365722fe542f0ceffc20c9a787073e3ede08de853b8155e8f323eb9441a7e113abf210f8b56dab2c61bc744cbb084f09a7e7910d003093922764a5bfe22c802dea66a6539e344c806bd4eaa48afb020ed5ae7b6b59684a60c16f95994fc293ba6e5896c9a64203854eaf533d09b45ef100f18e0c730756333598f944f6867be5921be9d3c931a07647121cf293021d0a3fdd96e03741ceebb0a519b7b20a84876180b4e0b502cdeff47903bb0c77072958cf5afaf79136262e04c560df221a0619f3d4fb99e88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he1938bd5c340fd79011e7e287504498f4f1246112f3f0c0c52a497c4b97d65dade604208012af63e5c4dcd109ee924a51255f8ee044654102b91b7ea365039f520440f2a2c9cedb28a75d317c042c14d4e765076615e947e9a75692a2db934aaa343b840c6d43ce213e9818b148483e071fe19f22e42ad3f1947ec178d914023b70ba744d6bef0007b7e848e7142fe72c629895f0fcc8380c319326b5d4deb8593f5a64f4f01f9b6ec8adc041d9551d472df9bd109a8aa5da843cfd3ffe712fc4fede1afdc8162efbe02346b8c7ed1ddd5587bc491c362391aa4c897edccbca389eae285072cc6a5b0dd9a6121850dfb1aa14790d3be1e56e3c9b8aa64ce5700fe217a342eecf721e4d8fe4d6f4c3faf0b1ee6a39170d174d7bdb206f7923cbd45b16ed7e5303639955c76645cda77a694ecfd9b1c9998c93ecf87e86c869ed309062d2837c42d19f5c1419896e174737e1d834c67e7283e1dccb52fef1bdc00360a30ec7be5b47ea26248174b129a044d551fece5948c21c6431bbfab42143b969c7afcc715548db7bb348649c34cedcd4558034d896aa3f5a8e50cf97dc80ffdcad8bbb8e36c337760ea56173c50f13c862f8d6e6aa692ba3347dc9b23463b5f953e7d493c829296120a483bb2bd76f5df230c48924e260e11a36050c50ecdff61086d254550bc755c7d9a65a00623d0df6321afaa629eea273c313dee14c7560fab010a75fc498500486b526bbe9beb6a4cf4255a078c5fed2192407a53f0d25848512eaab99377fad2187ab7ed5bb2fda5922a11ee8a80c0b2e0e0e9606ea7b7c84ae46f81bb53a0581ae50f4cd44c68e0441c9b27aa749831622f76cd04f879b25718031b194675cd25f86b86fdb08dd27e34d196d2a25119b5e027983435433726dddd4b957b88c10149f024ccc27ed36cea00c908a5e26b703ca4314e22e7d46b51bf1a950931b2babb5e0519aa0d6b08d15680bbf9a842f38cf70e41a7ff0c9f9b37c560e9ab81840ab5cdbccab0f241300f586d94f74989c02a5e5e2630afca7d85892df16b5de37b3f459a3db5cfe285821f8b2c03d2f9bb3380c56b906abbe2e6fa703b73e1d6f3fb8014aad457076df4d996e52d68cf83237d90a534207aed800af03d166dbba7ec9a195731e24f91e7bd2244834d297130ebcb9cb157509c251c5bf8c10755e8d0801cc83d5bbc8a07614de56e5b1f662a034ec03b99756624b3e787599e520a2580656cee4c78088524a84b90d0d4de949366d293d9d3a13f7ff3c1cb2633c086ec08610f131ef917f0ea2e12da11252fd583af44ae1bc7a7c3ada08dcb83f8211dff649a9d7c67110377327cf349b82ed3726a977ec87bd97a1fd82ee59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd67e06fbc37bcfa75b827b1397a4206b761f93837e8a384b130250ffeb3428033099bb1102e1cbe2aee1ef844c744185a1765acebefd584e17b4d4440be8e151abb7f0eae5db2c9d3a1ec1200457f50dc2c19a5fdef2258e555541bddee734d925b2fb2a5f0843049e9dcbe035ea7cc8d35d72b9eeb63845aed5d56092ce1e8f985905314844668eb769add3d6b9c77536f1e241e6cb2c31c61b7d5702500c0545aa0000363f53a70bc3415205dbac49fce3b41f53f1a0c3799f4228bbbae174a87ea573f39a35b01e4c288e3e0f3417310e6c646073ef291432e982d3cce55dcfbf8a86e37351ecf2fd2571e7874a2dcd5d8b31e8a9b3d17258036651c8ce5de2c47adda7aca871f55882f71279eb37b3186536dd2c39e09c976ef379004ad7b8c629c35f58ba4abfaee7ca2bb1f6f7a626da584debcfc19d3f88b6b073f0c287e1ce5d0934587d3506909a2d45ead13e85b9a40ad413303313b540e7e462deea0ff2894a881cc0407524219beeb97bc10d339aa4bb1a76b4f04cc77eea14ffc6b1dcf498006e02209e8cedb3f0410469ad77923577715c9d6856aedf4efd6349972f70308f629a8160989c60032106000097d3e2ddbb6bad9914aff098d9ebf92a10ace191f9bdf330b64b4f6ae7e7812db0baeda08c2f15317c6a8ee734a26378314d036c998f3c1b33794936f94363769e88a856bf935e79bea3cef6d00bc5e0357b9dc515ab9acad96b5b7af7a14aacc33663bc12f31fe87ca7ff5aff7c3131c608c0036e71d869a16123ef0b37636d95ca9c7a934788169abb31204f40e69a7126b20bde55dff5c58d9c602d122676548c662353aed5162c017ca4f4b5aca20fe0cbb6b3c4811488ec256fd6059eb4f6d02838342b97d658d1e942d680370bbcbaded5adfda64b546adeabe6e8595f24c8b80af7d4677adeae30e7c0a5f2f8b00e25cedf4a6b1575459edc949d133d55ce9f91fb633863ae6960ed179a41a961367e4261cf435987acb4642c75a94de0b4abe0c599b005c1afa43537fbc543320bcec19aa7036aa58b1e35e58bc7eb6c6499b3fdcf5cc01adc1bb4958f68ea545bc9184159e635d2972a2c47ca6e1c8302344c21a2029faf43017a5d15f413ad275dbe8fff3c92325a8d496241e036e34be70cedf17a732c2d6661fbba812fbe74f8e74a59ae6fb07002534f83e48ac3c007e01b58a8af90a48213f9f9208d5cbed5f439cb5c0223f0f2bce5b213810cd7bb9d90e7f80223833280a8fa339a7b7f25c3ab4e277053f66691703490dc8a926323e4dee11c924309e01906d69673bd6e78392bec7eb14e35e5ee62c2b72d1e2909d93473cbae84520ad7f5bba5812c80309bd074199ee6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he1afa807570060783ad81f48323e9cf60af78dbe80b85667b41131ef8b5a4136852d00bdd2d3810640706814b06ec01ab43f778ee78783fb0d6d58d016d706748f7afdc3278124b5a362b9ebe2a83e89882d091860bdff9e6cd1f33ec2d844895d9580fdb139650779b11596dcbb4ef295d59d9f8e1b9a968f881b10e813f6730f4d39b7a900f56e97e86dcf8cd9eb132cd67fb1fcb7a96e2bc7b11b9e503af73909c6f1675c03ada62c902af79e3ba90351451f02fff63c105372a44391397b0e0bcfa8b8e47be9868a1f9e281fd6a6880c6a005b0827fb8ccbe2d81404466db14252a07dc3ac43f1ebc864fe500b55ab256cb731614a1d1fbfa6f2ab756b1fdb3339c85b6b700b709b9951bc9c0bdcc90def0280b756c5a83aad59c459c86e3c00f5859d33f8e32c4e9822b5326a649e5cdf0223b854b4effde828423639256dc8e18171953e6f296e0a48b4374192532919d0e202bdb19d7a20712e7d1496042bac738a7ba0f7bec70c2240997a3fbd83e287fcc20100ef71eeb3541e4c201c4e86f2f81fb7e668a5b945c91239d7aa88091b93ca465f5e4e73a779c33975134ae395a53e72aee1eff3ea61f35156caec69b0e1329890abe93bb02e0423bd64c4695a7f879d68fdb8b2e99503ecd883bee4fb0480b4a514a02c08e28c9e9b57c03a25247672dd556543af73aa32bdeb7501bd267290902936487c07aae49fd3188c91b12a52780b6155d761cde3f3cefa5ded44e12f1a8ab8caf0d2ba018df89c86dd786ba81e9d7d3a7036ceddd84a604e737e9fd5942aa419e1856fd0ed5daea01482799b058a6b44613f79950b768ad307ae5bc6e96f90e1cc5148bbad1faf6378a364785b876f37072cafac9adc9999cabd82b5f2be9341ad9be7f6ae0bea33ca93c40bca2c47de05e2a1a56273e5a989bb116745fb6b8b222b4f8fe85d3272ef640083153ffb69137198921addcd8dead34e31c88070ccc07bd70d846a7b9616933a7d508ec686e9f3151615185d790b3b63ba941dde3502627f1e27d1da16372cc26e56519a413abd926ec6cb451a1a7f183305f4fefe227fe7e0102952792b4f2ac404f8d190a981e036f882ad0f206a8d239ae0acde631f64ae0f141bf278bfdbc8d75b60611916416d065b59167c1cfd4411b61ef0ef8a351f63de9507af6551c0d9f8fb27a0c0850ce86218484f9eb8508dcbdb99209621af98f7a5561bab204f422b4a9f0d7913bdd18a254db17cf99530fa963576507d03661fef9cfe29ce32f9b0262b66822417b291265bdc2ac83e3c2dfe3a5ac6cdec1e7544fc4741f5b2534807b84ba8596473f80f742277f26e111e115358a20118b10793841bff7f2ff1d138d271;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he8485c7a61d0bc66a49703cb2b7ac447a36621548ca1372865d8b499f2904c860b852ee1aa6c1d1482222dba0e10ac4d0859cb8302128c1613859c42caed1b3b2ab22a0daebb0354325663e7d3a0affc2be0b6ae8cfa0975c65344dcc23e394418c5414d6b5810e526689d933f773681b111ac785e5c918ec3d3a88936fcb0820108cbeb987732eabe625f25a27e1d353b30338ee96c8ff58643fe0771fcbfb9516bbc41bdac13a107ee81a2dc3b003b6d0e361c4f29f92dc653a31cf3fb4c4dd70297ad9c102d605a0de1ea29a3d01fc74e4f609f144a6585df365486bcbaf6e35b84b61e0e7a83e9fbabf022f446a1d26658706bcf6c0c17084d9a03828832fb3586b5b8ece5061754c84ee9f3e62cc311953366e9de8d3e36324b50928a42562ff7a9fe0b32f3adaa1bae21f97fd9928a0c224be61a511405fc8e85aa3af572ed9c80ecd68798c0a5dbc845ad6e882971c658c6c1526d06c51f5c4c0e2f095e3533f120012bf53a0614bb6e246cc1ccfc40c389a8226c6bf09e7645ade9878c111753b933e9a89448f85d407bdae1501383d1a68a6fff145fd34137e325978c5633fa07908f4dd90e6b3e1c6659ec647d1130b7d00c4a1bdd85dc3e9fd122bf2ef683fba65321efa91f516c03c7fac04629d0a079841d1059f26222903d7fcf324ad34d233cf83b0ec8f95b6af7e047fa2692cb778bbabfab63b0b167059be467c2a2472416d69a297c0bda0e2307bd24dad74b26e925f865d8a57326c48393c6b384e4a141fefdcf7367e1057e4675cb4cd96db4cc58f3c4eb2c8c226d5029898aa94cbe46c2232e32bb35053996d930f4833e84625ecbc2a63d9e480fcdbbe4cef1efe3f67f557cf6db4af2e3fc0e25eaf21ceb5ed2e5ea60a720ba9cc1578d2b73a7f6a66ef15b97d58d5501270c340c07d33954056dc91ce8d74abba5143f87fc37b74ed6c49dfcc0f9a182369413b82eeb2e1dad5a6dab39d1cb5b6c19e8981cd36bbca661e530d2c214dcfbc372343dd643f13a0507d1d53ded73f3b9d5a7428620418c75335bdcd89b105a20422f0ea63767e6f2436e55ab21c392cbc29fd267293cb0d2d7ca3a08585f480cfc5f2c1cab313e7853f60ffdf21fd09e3ebb7cf2272c5a85cde8663e63fc3922ad6073c04ab695a65c4805619d49baf130719632978e5fb41cc021e7fc2edd357ba5f678d01b05c5d7f93ecc8af5ad01d18e5b7bf800b45de3ed874577d451a2739c867481ac7b852194c71e8944265581ca2fd8f7d09f0b9c80a339e2d998b05607d704279f571c5ae866bb9368335803a95aff448fa607b62b81bcad9692a133ecaa75880088cbf7b27c03640bef468a288ee6d24273dc375b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'head8ce36ef0071cfce0b71d8b403aa0a5d87fe3ad1d44e2b512b3427955f1c1167f7445b5d9dc175a454ed0e16bcc5d3dd66ad5566192702cbb74789ab516a42f745b09a9e54547a31bad73320fa3463e3a1a46e9701229cf46086b7542b506d0b313e77db88fc94eeeef421e0ea7f765ebaa0b988345dcdd2ce283d39f7ec3b81cffd0d73e5eb27f45ef5e2e0e88404e0f26f6f99cb798d10ff0f65d95efef2c048bd07c56e7a82d62918784867f7db4ee417c8c8cc7e260445b30c229a4706d02e03fb7bd8d85c5c52bb850db7d2c1b648ef92b6cb47a9a06a9ee8015c96b602090243914034f5f4ef72da8299ace79840c5a7c0bb9e3e80c719b7de5ac9161aa7bbf6e19f3b2ef9a9b72c829b1a874fc411e58d9c97ff7d38b027d5fda0749ea3ffc8b153503b53f3fa622de022bbd36bafcae2c4ecc08a3220444288d227a3401a89b2db0cc71c7b2e1ff96ca74d7cd2abbbc82ded52d76b061b51d55eafb5147895bc39ccb5b8740d8bff1ab88385a0f3f2365584ba211d2017ad5eb15fb18b2f8818131189965562cc3b58e1c060de78323e4f6dd921fbc2b467b010c9710f60804c2ab6230828910f69f4ea91649458d022b91aa782a12f3db6a6609ecf66556277d760b85450fb47b1b9c246e502f81f5a7513d2d9d52049db67cbb8ff748a5218f7037a64c3351eea5406473d9a56607dca60f7bba2cf1982f0f4d74c72206c43b20431a4f0fc7864e07bf6fee911aacc4d000a2899440295a377722ad3c8070dd42958a2ee5b81110ae8d87c584efe55d23230b6dbad7e199e46b132c6663633844418af4e4d0aa304d55575457331de97592c9e5245974c0d98b1623473aefb7b7cc5287a235bf95965cfdf287bec0e34954b37853a7a7e61b5b220c02f8c54dc89faaac44a7add9f44b50743062b9c0be51fb7fdd279a12313c25a737f701671c1234e4fb929a8aab8955c7dc46a726f61c76658d6694671d633ba299579cdd47a7c801b12c2ad6a4ac01ec7e12a1b4ff36869eee329f54f9cf2a07dcb6c007a953b7666b64e9e758a211533625d0ef343d79a386d7d50c5df22b26fd8ac76dbb314e21c4b91d97a1683b49a516cd89c909585e9d0442a485fdb6f944961741823ef0d851e791d8a907c954de267bf34e84594792001b9578bcf334a9207c2dc4ff948b165249708b07960f5472aab83cd42c778124667e4bef02dfcf96073406d1356b9e484fa7fc7628374cbb0a400db78174f60bfad652b0abe1e6e56fb71750b5f686c77208c7328651d83295f90dbc4398b8e98298af41dd4c283b311aded39522db4e97a56e92bffb8850d34dc5b9d9c94c2e01aabfbb58793e1553974dd0902b5d556;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8977ee64459bcff845b9d14f1b3eba732bb8d4e300427fdfcf33dc739bf0c695c3c2a0f83ef31c9ee387fe1a069c793252caef67aee22aeff50a2c808b6ab02ad9c6dd34650205895d56a07f848b432dcbd97176a201f3509073b0442b833903c9bb800f2cccb0686889b745fd55c35b799f54c8003edd32e2bc1764bae525a127a014cdef98bc33792de37d5edb1b046003adb6b57d55b0c13892e0b975969f43a900b51d251e8113475e6d9a0becddba83db4f77f5e804fbcc559621e65e332e90f806df75442a7656ed4b4c6f619af0c2adb47de671520d8e162632f98d3bd9372bab79fd63caf137da367795f7e394bd960ec7844279549960c322af39b6c8bff20aa404bbd6575747f06df71cad7a17457d36c4b7b72ee12b974d7c68e1e1eafe1cf9b86ac807025dfb19038448d8cdd1028aa6f392392b18b3ce5d4a1a8d815a9da2db3b188ad38e0f76adcafac1b37b2ce04dd5e7ce2de3d9ee0a0e0eff27e2dec63296161344c10b759600e9d2e250446853d81392cb4e38cf0220faf34f51208ba5560a8c685328c9325ad7065fb38c6a1225ac45493a2dfa397402fe3241cfd2e19f68d4a7e105f126b3fd91278c56eb122494d8710da855dde8412edd76d1043cd945a7151e46888532944f0ed51bc62442fc1ff37c55f9d676dd0950c3c271c3597b3c67a39750d31f2fcbb24eb33035de9eeeddea5e7d7fa8d1b98fa7c57e1a7996b3ff9b68f7dc8220c69cc33a84745f2b23970f8f63779f2aece6bcc6909ee6f1565368b01dd586a3745670b349a6e545c698bfa5b55e0cab9ff619667f142503e643c7c9b3ce6bca1315adfb507ffb51e3343b4fc36ff901b12cee5f48a7978262dff1bf63eac71dbdf08c3d295f90b028e42ab923a749feb8d5cccde060674cf5503525dda053355f83c2d7b3f6503462d3d7f814fe7382fefd03bfd7038a7d990f3fd1b8dff5ffebf7488c014344a649dbc1a08eedeeec465daa51b69e6b26d955026c869502be00a42aaf899e2a0f46e5b47310560936e3fb8e68fd03978deac1be080afce62b122d03d4c93ad16cf53cc5df620dfed4cb7c5fd3c3d7a5957a669c14c9c336a4e885a53df1f6504c094f552c18057d66ab172c7f1bc7d672d72b726c35ea3be13d3b2ebc1a934df735bc2b729793effb2a8e4a60977d5981fb83d8ae423e6ed58cb248969c6cc9c551ffbc4dd6909019283030507ce4e757362a32ff3b6373ea35d94ede1eb4337a6efd7bc279e8a8baf326de832d9cfd7c523deca80d4d92a8d4d77199bba2790636c2c72c313d3b3b4a827f621d07f5ce6b61b14fd5956316c503ba2d3a88a83f42c1817f17fe658519a28429f0811d4d1535ce1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hee7fdc2fc01f8663740b562f47df5cc04f0eb7cd5fb1836c838ad427ed383a4691e9848fcd42b3e6ccf22db546101a079533702f9f21d9ddfb25e3228556479936644112462780e13dea54299c8857a811ac515b6be03e2f2696d9c0a8951a977aaa2356ba97c0735d9e5b63d80a051531206cfd0610f0254fd503a5a82870c2210167f5f8cbcdc801f02663cf30a872c11316d448c2c54afca10f565900b827417d5ce2db7ed0ce91bb0eb886aaf1e6120cacc012b76cc60bdabc9f74b51acfd755731454fa85621d1ca340a0d1d529466173bdee818c97fdc4df6b9dc529af0de6efbb537bd35a550526111d1c21f0498c085b4e831da33a7051f5ead2318759ca1adca4ec079289cc83f96f05f4daa54755df23c6e2a6fceb879c72efeeb1448e26eb8f1d640bfdc02ce22e7716620d5def4c7a17b2a6821a1d06da1136ad6d6d1982142c99e1914b0bed877bc3eea5578f3ba211aac333f8d3c4fb4020000492ce7393599618ff779b50568d3d0e3407d24c9fbfc1200ccb695000a53f640a7f39ed57b7e2d860ec7ef526ad6da1354bcc5cd7b2ee54684bf433a576daad9db889adfc720e13cd2a7d3378426df74de74b5d1ec939fd06d2b79a45133250c8d9f93807fa7641efdfcafd308e49b768e6a3a33929a9319ffd276bf5bc1ab92f74ed2f37e176fe5bd93f023dc44e5164f7dfc5f02fc6d87f3916503e9e92a85fe4ac5705b6e5e0c85fdb4680b5064d11860cd38e1a2fecf43e9cebcc6256119c9a950403826fb78b8c7ed1b91843cbadb2835ef471fad7d33d393bf0635ffde09020875674b7987da55454feebc0919cee7ef2200260d4b21840565f94928438f7fdfa6891eff1c2ab59e2cb6b816a2225ff534fad78de6d375fb245a8781b96fa4751d8963d8be08895099386a1c8a26cce38afc9f7e62f163a2a16d798bb0fc8701841c107ca470f4356b2f14bffa4dff7d64cd05876fed910813efd445a6f498967189a4431e2ab1307a504ffde01ca4a15ff5d4c388ad4d49e411dc98d788036e9dfeebdf64abeb9d75f1e92d02874d149528220100bd8562cc331f1c57d05d469d5ac20cda8bd5af0c50a4e0c9ef51d46c89c9242bd54d4ab4745c60aaeb84e37cf7109155c7b2c9a3683d075cb10d417adc10f8457367350291e0474a552d7dde7e3b70aded2cba6ade53006c9850c76bfbc4ff4e0bafcea8bda48a2d11d381791fcf2048e2d56c5da89859dd68b4884164733a985e16a45e7396436ba90a99cdba337e588eca305757a57633f358179536db6e980ebcd594f45e5125ebdd3dba3754bf3fdc5ce1d2a546ac20cdab703a299db5a7b94e7036cbe5586679148c1a74b967486bf56a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he36c597496eeaa4552240f4ea314e0ad8f1f985e2668738af5fd0f9ff203198625406575d40508843005b5fe28ccb72ec930c216e839d122d9a526c02ee0ee737e644e069768300aa1f069db4ac6d3d4185c153226ebc872397cfd12290319763469f11ab61e32e4f3485dd0966fd3872c7d41f4aad56790e89f9e1f044cf31c16cf7952546f765e0485cf532be9cd453e6283105048d752afcfa707b7971fff98506567c8f1f7a3b90b2efe70cca0043048df636eb1da4c5c0037f186a85feaf3bdce67ffe4b0917cb667655d01f3e377e4cc73bff0e726eb928f7ad248e8856910c270e340dc02478fbd2f44b5d6bc3e171ce079f9349b2e1c4f522b0e546a99ef236562682d5fbbb22b49147ee4ff9cd98d3309fa77a881288c8b589f5079e6864754bc7d030cf6826515f35ccacc5acabc40463dcf5c0fb063e9c1e065667ca51ce92e3a0486c2770a1031146775659cf9de15e2dd47baf07ab806e5bd24e2ac26b7c87deac2186e08dd71e81bafb9032049ac714b8eb7671683465cf84460ca89bc8f4d9aaf23ec0183fa13009e529ffd147ba7bb6005de4faa078c89104eacebf73559124ab041fb67c61dddf4470047d418053fe519db9e538d33830a163f381267581481f142d5ae1af3350016cf79b00b43de03c4b01d29b4f0d2730a8733d9606ea0fd3c02ae5ce7510c4bc249b9e7fded5768fd76d9514a8217ed109ae03ac8856aa6b5c38205500c1bf925eff5704339c1c174b2ae23b37958f89dc751c73beebff5510f45feeee269a731c7080cd44a2af7a61333a6573f43f76acccfb0d25bc68a397a99fa0252486d9d3eac18cdb003efc2f3da1d1966bfb32390af1ac5f0819633a66cb76abb0f7696e27cddbc686232fb74f5892761dce1e911b490c7de44dccff1d64e4658100fc0c53b428e1b639fec3321b83f3478e717a76094268936bd78d313c95017fa654ce9dc8829e1ee181c1665872f710f1ebd592e13a0be804861ad1efb361738e4802bbd28d41f5f8c3e02e8bc35b8e847df44d1996a0c971bf35e44cfacc5a1b48b1aee8993b2b00b81592e7a2c2bdb5befa618a28abf6e2e434d41202b95cac8e0d0fd3067ca5b8684a3fccbedab7712bcf535c5999c037611322e5929f25e9a17cdbfa5efdfac764c9480eb3d62a1fa111c33ee9ff855c07629f7eadc6cfbc2c16b807c0c4adeb380abb6574f730d9b19784dfadd2e4dac3134ee834b8daaea630648e6d2e346bd2256a0dc5c81445b9912848627e69b8ec6b70c3458785bfcdc39a1e672c0e1c413e931950d17942c7c6038096a8b8e86c81ee8a924b07ab82f5b6bd7103279d29593159c39b45ffd946cc477a3c46ef5acc1a87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he8c4ce95e625823a93ecf7b198f2e416b9c047d0cbda282ed6f17c1064fa28671382df98614423de55688fac94598ba0e34b32c9db17b4b281035dedfc404aa8ba67f975b3ca415c0376aa8fedbb6778c359896ea89b41f16f587cbff45a05b7e8ce669d70cf45cccc1b9a2bbe27c25f6e8a1a58ceac6c8735f8f7f82148db96f93774e8f59f2dbebeccebade8e08ae806aa319d0c86028f5a82d4efdb90e755933e9af63ec89b6b042e2d62a302b30cccb098e2ecdf6866fa72b86ab94dbbc5bf18aadbec36acddac5930936cf47af245a1a30628bf904ef633dc7716144a57996936edd361c151edf5dc90ee0c62fc4a9d2bc62d6ca6f808578368a880c3d6ac0b71d65efac7e6c41d59de93a8cfeefdaaee6ca895abf4383ff87f7b408a5bb32d5058f90bcb8945bbea9641d157d41792342d0e38eef660cb9b9cc19083d54cd6c0a5eec0a1f72484efe5ff58e4a71ad56b48dd0cae6d1e375e5a6c539a35ff5b32ed79890373006b8105e38083a855d7e8f6cde9e97ff43f2c8eaf5c086b875859eee54413de5ec9cdcfed6bcd87fd59fdd726c2869702c663507fe602fb6ab31347787184b2dce925e6fdc7ecf4fcafcf24772b8ef27969ee61a5f0ae1fcbd2ee7b6f6af1454babc674f362ab6d2a3d75ead547ebb921c60ff26486f2c8c88d42e4c82cfab6e5ea6ec14553475fea6bfa3b4e3020684a3bc1a45a39372c8168dbd218a9bb6b6f7f41e86f69b57e540e7fa84c8e871d1f30f8ea7a88e22963009a36a4056b0c3916f15bd3b9639ad2430aad3f0c9487f27f7363907a5cb1416f145051a3ec281d82989cd24193d83efbb5b2e1df48a9a020e2500a618d43a5dbcb1202a03322692761ac3cd85c10d553064dff1135ea020b191bc509ba6aa3a38b0c1f9d4ee52a8fd6902d962bdb1f2f6ce27575524097e78433f7a1f2eac47d701aa966f8730acc867cec97c79dc883236d3be7c9f1449abee0450165b09e9a8db82d465d3261e66a8907ce0f326f758f08546cc7017bd9a558a05748f7ff278b84402d7dd8b19951466f3a61d1c586169ad0c3fcae17da4d45238394d7c5691547d10083aa9de5e455ff98ec923960bf2fb1ac97d285b41f224e4d0baf4ba1e4e59c54eb979fae29953c8a6912d985bc2f794063ad37d24329de028985efc41c713939343461fce56b6724fecfe386611bad0c95fb0794dc8514513bb64c9d3e9a0da7ffd43831a3f3c1048d3ede93e26067634e7a9e6a69b4c5490d22b0abb843822b26f4e888ff3549a9298658f241d32ee0f743f4675cc0cc4ebac7f392acd9db60411eed84c82f88f0bd5f4e0ceb441a0eaa9fa76c75fda83321290692afa325a4279c532eae10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h67f61fdf7a01dc640b9734065dfd50a8007c75a4825f306c528bc4c1fb450a07503199d7bfa7f63c6e78770c4fe51e2bbf214f856930bee0cc35af0f93ecbafb22a3c56f3069f94bbd273f11436c381b6f447cca331a0aec96077679ee70fd902a816def60db9b09d91c5286de44b88d690df720f90df5eae2f7f21c7972dac6072f68a79fc0266a790744fd456a4a19bbff4b30550a2cd9521c10e9d0717ebb58b76ad350fe6707ac9ed17cb0e6b25b1dc20a2fd950e8c693613ae8035c6db0a8faccc7b189a3abbdb59473cfbb0eb98356c458baaa443fd056e3f4d2e74f0a8d3871879ec767d49efd9d300d7bfc29996ad7fb67440ef6c3546a4ed9b6fc92fed6a1280cbb0ce1d63364a5aa06e52125aa78744fa7042e62712ef30dfb28f75517ee25d316244c40e7fe8602f52c9caf6f52cb31a72fb00441815d05db8fdebd7eca33d3bbd212f7986e4f7e68c2046cf5896d1ecb30e2bc516730b44712b0c38c64c96ce630f8556a71ecf4419453cb6a3d9150d898b3f524612242e1a6ac0758a39e50a567a557d4dd6c5f431299786a1496fca2d740238e48b4a7616b6f609f85abea608c4ec10737544b152f3a63a8f5cb63ccf9b4462a7eca82e7e4dea5a422bdb9744da405ea03e3ebdf12ad5f7a30fae3f23a1c6dabe4823a338ee2f149c6101757d0ab09f4a7ce0eeb893ee142477e1ab251da932298925d4f1f140340bfbbee126d46a4a7f5488f29c37fe33005f2647a4eb79693c0797701aa58f55ad962651f36c0e063a56ce29109da62839a7aeb915bca070c5b9f90a82966eee13c7c7559424b90e972fb63ffa71a67ade6279176e3e234ccedc4ec3f7774efda14736f7e787e3d715f88e5c534df28d6f08869d26c4b5372baa4bbfc832f76cdc0ad759c05596de3039d74c661925d2a4cff5a3e069e5c5b8b51a37fa709597a0145f82063b1be8da1e85d206d1270ae0f701cbc3665b0911f0a7ea1b52cbea439029fd80dda98634b4dc71e14a68064b35c984a4a44c6237005198ae2373deafcb08996bf3e16e7585e2ab4785c77d01c107eebe81b412a66fd334c4a9ebf82f72e15d50ffff556ae908d43fb79dfe87aab8905fe2608c62c85065046305dc967b7b231341319b3258d58f9705cae821f993ffaa0652413e85898e6d94910b49c5074a08b3a7bdadd65050c57735c06396ca7ffab6f1b58071399462a90dfc01e3910e847456b3d59a73afe0cc944c5c46b63f345278be5783b7ecd5efe86593f6febe7e9b0ca5ec895906b1b378ba8e04e28eb2535d2ae625c12334a786533c4208a44f0fdf475cefc1e75653b1a82a55e0d03a68136c1578794bf9bda79945026d3a4295a05dbda05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6d6956bc9c540d34c7e971a36c4e5c93c70b3d937d1cb319e8da39e122d7a96cecaa924ea879d8f52b150728084dba7089d31f6a99c6f8e1245aa245248441b570a364fe4856f8476c75926b74e51a69321acccda2f9068d343055e99ddb19e3cc7998333e311babc5b9b24e1866bcf832c1c56d6a1da5be1f9be7ec01871450003271ccfc39ca89ddb5d3dadc944ea147bae39fb7a3d2483362f7764c26ead83ca9c6762532aee7cde325e2bc291b8d03ed89831171e7c4a53f52888e60588ce43d5b399e43575609da5727c4ab2f548b14cb6afff0c371f5bedb75df24f457b95c84e66a93e5b1db1012fcc67317d32221c903f3c36c6c6740049534e1a5d98ea91b18d543da0e4bf9ef440928b5c92d94461d7f8a387200f6313abf265876bd0336b360f3cecf72ce50b93092bf35152ad83a872d05be96520e2aba90bc44856c3a19b18ee36d9595043eeb7ca1faf643484f3e8ccd85d0fa3725246474f5cb4a7c951ad5c6250dfa5e7344ff52eed1e924efb99bd7d2026391d26a660742581b1a302215700e9683bb19370a6288b14077b57d89f409c13ccc1f151c61da3c698693573e391896029504171da2b15d5663d19dedca19dff6b52ecb05e0a951aba4c0775ae5dabb25fbd41d1acb102437700c4cfd3b9f6fb281959f7ca6d308307fd4ed4eb696777b8edf1b63931ed3e629fe1f0b433ddb1a9efb8eeb60a92079655ee6a90032494130da33df7558cbd2b303e6c73fd7e66576cfd375ec0c3b8439d135a6909c576272718824f72685b6dce79d943a2acbdef99d20f9e101a0924badc3acdda693959e08c015685d635e37a9aeb649ff27eb58030116a4841f2d09a2c2cfd1ce905fb5b6de99132d5553a88f561a353bddb0c49a0d19cf81b59d08710319794c032b6e14a2c3a616c9f1d08d05a820db0fd43b00c2c1f45b766b4efdebc1b40bd9eb40af987b55c0aed8ac0215312a17c8d8897753fff4ea26ac9fbb7da4cae933dd2bea509f1bdf290294606db2ad04193c36c01d9aaf8548be73fcd11535af97a6e6128a3f915343db595d866b5f97f950cccdc0e57fa99ba4aaa20550833f60540c5840c1b3a5f5816de7dd43e78db4031634196d113584d9b25b201356651a3aa433f24e39844c5a8e065c56e7de16551c09ab1bbb2815195a2f2b1b4e32e11205482056d0b1a7e3c86f338b8756bba20149869114d124e255db96b8f9f97e86c32b07fab4e0fad04c543f9f826b8c8b18af2aee6b57b33f9947e34e4296892120aa836c6440b77abaa2ef4a920b0bca5246b71c520302eabfed69581dcd0d7e4c17e8682aec9d6bf30bdf6df6fdb7c7b38bb36a43280abb65dbd69dc22dba2b58d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3f68646a0eab9c5880d63df8fe19b9a632be38aa8f9fd376d11d4d533dd69caa3ee6a1179e78cd7f684db08607106834d6eaa2b2d3949fdd4b4909e9f26e0707aeb07f5203cfcc91f4fcdc22a1c00eb53410099e90250e2090c5fd20c58f92339ffcb8677e4e2ecffdad880383ca11e4ab5c494df96e5fd1993797b6f1b83d998a51d5abb77e597d9fe2db0e9d830b6e1244bc0e720c1a2935bb806efff20b305f702cac889325690308816753a20b683b07cc7ebc7be00a290877666a3cad4d9b3b212f4ef69bf79d9b9bbe7e6ff34547e4ea5ccbcd82c81cc1b9d0f0c5211ecc56cfa05501f4dd4179f3c342de7c27da971eeae6a6e5903f6a9157aa446eb6de1566c57988491eec47cba703822553f23657cf44c58ae04eda0427cd6ae41b7c42dc29ebc06987404b12ffd948f510b6edda19639452276b3ddc472e1bdc95c45a25a677642a04316217b402929e19cb490bd0e6f92b0ab9f0fa232ad212ed3d60f9c45be4b57b21f639ebff2acabac385fdb70feb4009a587435cfd36fc558f618618cef59228e8853ec5424630afa423c1116cfc02303228bc012317f0a3f2ba00d5d949d9d774e5ad6b6974bc489a45b1cf3d803227ded27871def0982ddc495b36231a0f7ddfd1c46fd13eac41135f9fd34be033a1e233eb79ade924dd6898230e2d07d36a4dd4e9f739607a9b6c108ea787f1b1eb850fe163f2272409c2d7dac79ff0401fac8de14a9e2f31c4e2d3e65b0b73940751bb1e2b84bcb0fad3a8f1a95f2fc04c0b4f93a69f9bd091b11a939d60d6f408c62a0c736333231bc68fe0b125628f20488572ac62c598604332b2323f6666518b87f4c4fdd34ae2289d5b3aa6e45618fae79fae52d4cd58005a597be792c5e4f8e9d5075abd7d38c64b695076505ffc98b00ef68d212465a188430df5b7378783173e2bbe35796079c2e02363fb574ba1fd2f527cfef09abcee29b261429b0ada230e1919e61cf411e7859256db814a6cd40d7cfbf7eac0a7d99e3e50c1a880b5abf4a39e795b35ae8b5977345a9f7c6d5824ede2a9c6b080a2fb0788614c1450f2291672289149e5d05bf0c972c4135ec2726b00276dd59a74ebdc3418841752e76642d1797c1552b1e2fa50453621b72907b90fe07748a7be0f5ad09e5eff26faf74de3b8ca959ad66f5f576014642bb8e7defda23cca8064a9b941c0065d43ed1babdfa9ee9bb36542ef9ddeefa0ef8a9fccadad994aef44de1541773522464f4461d2cd645e69d2985da52c4d4d5c147bcff6e7842ef0f3233944ea4542c89798c506525f7070e6b6cb5ad498c13d002859336151fdb25479b1628894869b2ba5c3eb95c3a842fe70e35eeed0ab400717fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf158ef416fe09da509ad0ca79f3a442c2dcccb47acfe19e03f62b1636bf8597a51fd5f214844186316d122370947af23535bce191a172f95cc58dfff65474a1c327a59efb93bde2663097ac13cf1a4bf7556272039f5b6307d61da5f7eca8c2ad195524fb534fe273fe65a35190427ebe79ae53d666422719b7a1c3ade7808325d35f4fb142cfab11c4589b7728640735025c8c79fd406f0b9b6fa764b09d929fe17b09a314a5d9ecd32d4b4bb534cfd044fb733af5ee1d0076eb7c8c9690e8aa5801b455b926022fac5df874f8286f88007430af1f2cb2f6dec6ec7822d0355f5ba15e1974b30ec1702d6a6771f878a81811c7e7be3481a3ab8c3e3438b0bfb07cd323ee2d7c6970baeaa6e353138b49aa4fc0ff46d8b46c8cdfe3b41713309e63ea6055ad707e3c019d2fb3478477f9b7a0a621251d3d8158a82330ce3fa6ed42b3da56cf6188b78fcf9d9b5ba7325914df096b04e53133ad279c7604d5e8fa2e7c59df6ae21a3131e5273f48c63c933520f41ada0d89d33d055d6d62e57bc40dc1004167f518c4462ea0c216e64c8fe15cc953acb1ecc79027c613ed3dfa55bb1cbe5e86783323562b40e848d572d469df5ca969b3a416213622e17d057b16bcf71219ff0161da62684c4552abc2ce50cdebe6e1e06468d11b3147a3408f01c754f84db5e51ea618c37f42d689cda3be92e8d3c10dc7e3ce6066836da4288eaa08adba6c383dfa365859ed91664f05bce867452d185beea5d75a9b373a16e9d4bf82fc147b19c71d2c5266fee1f015e3bbf07c535759dc33d6ab7ce68bbc31b8580aa266ab773cd3e06dcf8ee462c1e127e60f3138060a5c3c78b566f778544defa3ee2c1bb7816d624cdce7e7da94bb408533dcba271941677491438923cc99b570f45bc2149e6447c56a4528342a1e1649a4b179775a6bd6529bfe82a23c790b21647090dbc3be11c1007afc30a3cd5de7f573fb75f8d57a3dc62a70bfc73d202f8de586ed5add3ba29f2b7171c18ead13227bcd78a976b95e5660cf796e9eb828b4073f49a75fcbb22da410962dd8ac91f1f4079b6d8dbb8f8c0192775c033ada4738aacb01451b8a093c7e32789227dffbdfb6b2e8ddbb4380d59ccf8594e1bfb6c8c83e9327f0a0f7f4a47ec4e8c3d4419422e945bc3bea1451e86f6c761f3f5303611c4a8b5fbecf91b4d03f9b68b69a27be32d270b40c30cbdb616f1220f431a7f14b5384ffecbde497eddafd205d6ba6140270e03b4de99645e78aa3daffee90272739625163a2afc4c2ea7446c0bb27b79b659f4841ce704e58f807d63045400fa1d43c3340b6e5d12534f3f946fb1d9d51bacf9435572967657bce30618c316c2773db23150;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd54a11120b539f0924d40d66e1ed0a6fa20098835851fee5302cecdd35b4774f1ec5992dbd806d07389d445d2fd4daa2dd13f05c3c6084c06ba56162d02a41ba8a3b42d2e984f1f140a8e1e78b2b994d8f4b7586b9fd6ef4fe12a61257a6e6c5904e42d595ad279d42ebf6b548f715539259b67bb3dcba4ffb36aa2890207e16f264dde2b1e2e7a9bf71352e47e6992cfe15aa94d716d9fd0c277b20f341b496359292fa8931091a93cc00e7d39c5a4f6652ff60d16643667b85021897aa76e3cb36bbf48cc56cad6f76609bc28fed18e3334ada6497c1bc97f7b2fea90da84db7c8257110de9b6ad61a2eadef386f5218efa7fcdbc8437bd06cded4c676f77a1500783c58adcaa5d02b0a9d6207504e165e86d7cc754e0c5c1be139af473dd4dc02846a39a4afdaddc64f91c77f0d6845a1373d1936c3ca0e127730a3483437d179bfbfd628bcdcf4efb2b23182ff72d64024711807df45200b512052060ef088b165060567f787571037116f79ffc6a3ccfb99ee072cb6c72f05f2a35342f5e8f600509611919bddbb6ee277ff589cb396603597e947e4babecbf4ae68286426acc2d1fd92222786facf778bb0aae60095d31d003762127922a6260cb6631ff16e6db453877834bbc1842212e7f5171d7bef68ca1c5af80d98e3a666fef178560ab4a25894c18ee484122b430769d7f6ab94cf013f5c2fba7b343b98428bd502231419742196128372bc034e7d2c4c857401a0da963f6e909592300c3f902b85cb1c070e7f02b47886576bab801a60badc87b198906acfbfdbec519c5bef86e2ec6746b1ec0954da1c2c0775dc123a32230b071474727f5ffceb7f0d5c8d8a21071153688540310de99277ae39ca7661442fd011b24053abd6f04be8c471b89d1f14b9c04908c854ff2c071727a66d20a727223075441be4bac5f390a4d34839f21543deaa03170c2187037c25657d36a34af45e716b9d6aed409b0ab7792881a2e357668261127af06aea1fd8733145b8bb297de2f57f6e6b7ad7bb7fce8ede19e04d1cab4b385590e4d82988c067bd93df5f8b463becd933f839dfeeeb87350585175b965c981078d52d072b61c176e3e04519b68d7298e8ee9ae48cb79c72154d7e9a92f8ab1e5845fe63482b78ec8abf6b4b426284da09525357d79bc45d0f28491c3d0ef65542b6c6e8a18479eccf89e407b796c827987f37808defdc21f4c0ae754d344cec76661a3711d2001194f99b3237b7c4a0524eec7abb40e5d8e71abab72341475b7ba0b86c1122eea278726b6e9ab5f619ff819127b7eadc8c8515b4737f721e1890ebf360249bf7ad33c522cd17f34a87a741b8ddeaf10376b32fc2b32bd6cc3ad76c1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc8365a31c7a3061dfeab484f51c17fa918a4c68d3bd23faeb09da5c460d7b8947edc0f85e7956ccde1be6b1ce853612c67116eca6d406f479547083783f6ad2b21406b92e610dd49932308f1e1aca5cd840d398cd0ada4f7c7d1ba0d64bec1df9fc45acab117ad64101757f14c59ff066a1a8b7aac16a7a552e8e4f3be90d3ec5c65e14cab30a2a0b8d0a352946065a1816462ee01ce3b4b35696dd0c6aebd7071f7c6f2ff2c570bad54a08b29bf518ef395375a05036d607e21df4229766b673b0906964717308609121a56d5b249f0b32f922e047fd6701dedcdf0540e4e84818e8a156511200eb2184b79086c409ce5b2c1af3fab5e4c79980a387a1e4d101bd20ee33cb43d89e7d90a8ff7fde1f17df5e359ea81934cd71a1d74573fb7edfe06ba179359e403c9f826cea95089df5dab5e5d8f9d99a2f92be2daf06b1215d68b90d03cd6de45f9cdb6215a88e459ddff7f9e9e7dbb4e0d3ac4c03af776ad5168c3461cb7dff6d8e39f5269b8b79739aac09c286f7a231d04f51b7bd01b30b52e9b40b50b63ee820fbb1bea7deee29208f73bfad851ce18578fee8caa23b42bab19626d4280ead5b743237dd9faf4c517d688b9c971895484b16f2ce760a6dc77962c06a7d5cfda427e87f1bd4920fb4eb2d659a1f12649c71d5f069734f448ce593502ee150cc7e1e06ead97f1b8e7af1c6622371903c92aaee4eb71977ce2e88fe3c28d92c81087d5a0691aed15918c5065cb0c2470b921ded0d566562d67497957bbc8da9fdac3b15e5adbb981c1b6144058e6290381606ee918da8a21e0dfd73c424e5d8de7c04c760092cf32723d083a59ca7737cdd11d10e11887c1d65cc9731c9dd6cdf5fd9edee986d1f01151cafc0be1704ea20130cea780002b4c34cd3bbd05442e4c7ec2edabf90247867a1ccdca974630d1e1f6943cc292774e025a5ccd978f90cc702b5012dfdbbc3c5ae53df156f374146b379bc2383feb11e111e86e4198068a2d83f92fa1a8111932be08bb220c1f2bd0168933a1bd4a28e7193059c49e1f230a299ec528a34c635338a0543274083f71e83ae470c283a3eec4295944096f55c3c9982f6d2062acb0b2ce460de58abd40f416176d19dd345ecbfefb3b8f679b3d42ad1adc6f55e1afd7e29a3b745579a6479748dfb279d89f228dbdba77742624fbfa9024adbf3ccc5fc28f68fcda0e093e1f4d61c218cf03cb3579c504eca70998ae088236ea233628efcfb508b6e9230501f22a301fc43427f2e4038a88cad15fa1cace259f9f3e578d4c16200fc0de63c7a1a7d630f4da0d21a3bce22d26c0cd647f49aac558b865aa30091845b5202879ab36914183ea111fb155f661c1c1561b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4936bc849451792616271d21b3440c638d507482dcc0d8b3bc0f91f1491a40bcdc4736ddb97902350e2ae94f09842dc44917fc89b5ecc7f3c7700d914df776b05701c0e4c2ec45c719684dee0d66dd7a5f4625bd39b140011859eddac82e2e7e6587dc44fa391f8a7b58365a72479f7ea2ce1e101a9086eff121eddcdf1aa4c7c01b6b69b1f1faa894e8d6e9ead42100f33ed41aa0c1c6114e00c85534b523c431c1fd4b1467a134cdb8a29657adbcfd695308aecfb5c6f22193054e825c1138a68b11821e314afc0a24fd25878a6c13178f0118bed66c964d6d9cf4c4578be5a0e6d7dc5b8dc88e4f606366c504bec6cf752db0ba73869d6e2757e6d9c06fa3b2e0d254e87fc6761cb568a971b1e8034b6e1f12344514d95bdc39fb70d5709655c470e77c5cbf2deeb60f12f66c6e2fbd0286af2e8fea82a35e0eea6868216caf901705517e6ce141da06d489be8b1c077643311678fac5d0203000929f0369f2a0016fda9f25b07ea4bdb20c3b0044ab226d3655a86c6783e10cdc1d0d61a4608b7ebc89e4190193db52a62c457521285811dba7025adf12888cfda3f2be531ba62185aff87c556646e88061efddcda55c3ee5e76bfb6780a2267e42e15484ae32b270da6a38c21b06918b5370dcd9e9a8aed517a9267cc6b4476cc1c8bfc1bce7a59ededdd898b058b26d2781119a65fb241a74a6ac1c36e4b27645d7f1b35bd5e86b4adc46b577f1f1b5809beb72ed4c63d049d425e53f4bd9a92c955fed8afabaf34f42f7322a71af96f3701c71d60f4cc19ee74b26c56f33883fcca8c75edca0fec5b159d2b47efeb6a22f628e1e5b98b98d70f515ee0074d500ab2a07c747cbf1845147c8901341e30288f88547cec1e5a1f8e948cd59d3c62be02c1b9ebfa534e683d2a75a5b54e1ed1b191e8f6eddebe894ee5edd35445e3ea911fd172c462a6044aa33b9846c7a568aa1e5aad528e88c09f045b278a9b9c7c2a9f5f0bb2650412d8aaed50eb042ab2a1d3c3d54c30644b7033be4a645de72f8326cd1636126f79f9a2c9119f75c5096eec871596a76f8338cf9e6d09ace1d5c3fa5c0272089fac905495af4eaab7580fb6b4baa375d66fa1e68ff60c642d96df935868587f66d7c9995ad0187949bb863a38f65784d546919b7d8c1d9fd30f7d351a831e31a25d8582c277356140d5513a470a0fbd9b7423af6315399419216f6e84d72b5dd79a6c6bf3102be93a6ded8001f3d764f5a31ed258b74e5ff0b0e7cdbbd3e577b880c18178c80f0d36c80357b99b44cec21c0f88dcc4ab2ccfc3f85d0bfcdd573c4aa642418b9298ebd7b3b937538439b2e8d9a31f0b03ec9b27561fe99140ecad685bf94c494dfe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'haa49a60aab214f8d4862fcf147be980b2461bf537477b1697204182a4df64c9819f4da1af9845c430af46a74e44f15d5136daf5d6a8e210aac767f687497cad592bdd5819fa2e968c583cb07428bf03a21a48d02e4ba82d41a69142d76a90fc4f6efc9e653e9decb7031153a2fd2e76797aa435c6a68fc1e7df91c336eaed0001afbf6406d6e0638ff51fe734c5184ab9794f728851fd137c9880e92214a7b08e26262de9d6c3e1ba28dd2d47d0ab992eb3642014839764898caa027d5342d2a2d99ee1b3baee3e5c1d9529da6fd640cbd2626c757c58699c5c7d7dae2f8da8daebaf23480df28ef346850302bcfc511d7834c1900133a04f6f59ace138f2bb8038cdff4cb88e372034f600acf50bf5ee767db55a2037e5ebe263ef9fe0364fa5e4c414d33ea7a070d0025ba4a2ead4c93eb81271ddaf57577e02dd86e6c3223cc15983e3b5155d8d7a7f43ea0b55bc50d537dc84e1eeabf9fb36e2ce4b00a7ba6f6d1070d42bad466ad37401f24b86d831764239ae2ce6c1ed5df779452a21c766a36ae146fb2b34e9352b823fd06179487be4c8a5cc992d776f35995a32d358f7bb9478048265fef25c42cbd70be9335248ee80a11530a4a40f69c157bee6143d39ec3c4193023c5963a57313c4e2ef32277cb4701407b65da866a35a1d05b90c6477d253004fa36e5f79a0df2622001c6bc4beec3a91ba3fab235b33df6a80766c9d721f64f6b1e0af5f55d22dea9bcf17861f6362f870bc7149bf746f02da64b752d629480788ae96619b384c2954dc8d3c516711e27f519210559361d9caec433d40bcd8b0e00467d62bd38219c08d312b5794a3c859ee3c512bc4997f4bd03d414bf408c8eca5213e18a96d7495cc5680513cc279a3c4fa8af38e1220dc44842a5755f554f53d3a901a30905d6718dc3033536121a59dfd415b30fab20d3a148a0a8e4cdf9edcb87e0cf0148b69a7ed369e55ece752647bb736210ca773b37452e34de9ba296a7ae93c14771bff9ca9e310984947d86322b5d80b15c13a0f6202aea320300d39d8b0ae1c7c4023fcee2dad085692c9cdcab03c9c3a52475ecabe6739085e5a4c6d0675dd3b3443da155641eae3cb8f6847c23664202d9c922fcdba64b4ce8854045e7cf60eee25af6bf5730382d463ea097f0bb60d3a974597056d423a341cf1940fd54acf89e634cbc852993b93b8224e5082712c7ed90abef2612741e1bdc54d97561d65f498902a49b76e8dfaed54e2b8692262e17d4701bfe770f8f8106d1a026b634f296af454afb7dc9973e2adf7baa9e7952780dda30dcd8d91b189f8c6841ccc17f2800d716a8e73b7648bd04dea535c96af353cd3de1787a420dd7361a8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h31b766b1ce74ea8aa752565dd9e47e39a861d4381424937274565ae51883600bef60e66a2deeea8e9d39255183b729f44fce29ceb40f43d0537db8d64a3c69a58c193c49d83145039d6113a20dcc02db4c5661ab06c0a7e365002290e13efab08f184db95a70f0033dbda0727cc613afc4fa77b276af95598bff4b89740c816597dee0f835b60a94dfef9a569f5d21002a6e607fcaeffae78876aec1183d908370a4dfe96915fa124d23bf2a1d335dbaa2c80deaee3d9b05c2365ffd1aac0d1db0fba9dc68582b671aa5a3d642d330f96c5f9a32a7e83e5dc36d2bb38f5b7354f115d2c3835dbc05ed6aa765e0f36e55a778399ad92bfc0de4810f1adfcf0e10a78fc385d633fc0be0c46770056092f1602a09f0bbbc154664c8c1ec57031e92a428ccb20d120167e947c22778c2b1a67bfcbdab09c8e37c1f5f5d3aafdc9dbb7fdf177d9aa3b7719cca6f108dac53b69ad3f6ee230f27e36a6929c4aa571d33d4946bdab564e230d7f8149fe33d0ce877d561864e0d1e1aa3a40fe8a8e859d780eddff4cd3cbeb0dc27692c2886fe9d42b693e19fd5ee444f1d8fc2015822634a644805d291e35655eb43d49e957de2878e5057107233a33186b4e4b4b58c20095eb0e3c1ce82bffe21d15a7f99c53d46bf974de00674b1bb8ba3c807cda118a11683d5b5ebbdd6c224d4569cb270881364aa383281f8baae97c8bd738d5553ec02713e88b0dadf770b46e89bf098a1bd4ffcef9fb7312407885f327918c533d226f35eee1dd6fb272b3a7ed1791544c210d0a78e658c317d5a48613dc5894547f370c95b8b7a16c38aadfb1e80e20d31e7be55941d229c6a409ba4f9fec66f0decf5f77cf086633f432fb8cd373212045b4b3b51fd352d619b7b1be7d696706ee3564365b2842c0c695b0d0ebeb5ba59aa248368622d4760f116f41bb421c963f5aa4ae2f2a9d18c31f6260f79643bb1b7517afe0add5ac0788eda38e99a978a0f7e3f1194ac67ae181f38baf3e02ffb84331e5624dd628a528eda0c0af02f98ca37c51e4b6b5317d6a6c7e4f6eb96e014dbf1be1e75fb4c31366c967df41b0bcdb90e27b3f39d866b5040414f479ec82c55965488171638289e88c6438405f36c7025ce6c46d4a3330db8ed3b672790da1bc1cdb46de7e34104fe3265300e1878ee368ea3de7692192d91fcd71d0d48ea4e62dbf8a92b1ad45fa5efa784d27cf1da6410c86c552557da0efcb8254d7e65d0b4f1ebdc0d28406fc7f650253f2fda64aebcb2062e0ee2aba1c8897c3ef4af002ec2bc8ee375ddfe5e3d3bfe7202bfc6f918d83082a093f54c89abb4337131beee466f96281d9851814bbed1f0957c515062e56796f12b053e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha9d967da2472e83bf5d3a805089f964a8ae8db402604035fa5eddaa274dfe97fb6384496117df7ba2fdb28043834715d1c5ba2d9d021762c778db657f0e721ea03398a839a3def561a9c69c16cf170b26646d725bdf1f49c61a199b84fe8d6eedc8c6a90dc3f12d647490babf3ee8e7888bf7f33c35b35a07d4fb25c21ef64feab7464b01a97da30230e9a75814a3698f30fa21b9e474cffd2c28f908d53765adc1727138e6c4adfff2b3292d28d662151d5af3dfdac877ed86322ae1e32b447f96516290526d1b5c2ee1a29b79dfaeaf8c100fa2b656735b859087e2d040f511d06a0ce829f0ff3a8570b0c3296d933fd858bc5aa8a659f2b92425588689b0a5d3f00ab263c341f6fafb870da8a1182ab60b2014c7da488871a4bc7b55bbdca538aed9090b099024c5a7d8f9bef3c0d70c715bf8e7afecb43435767dd41c5f194cefe81ea6d4aa9606e5846258d4edc7d0a8383198ceb8399b9a655dc029a8175bff00ffce8da22d5dde62599f1b9dd6b497668d08b9c51715682c010bb43c9147eccc849b864e4401845b3ff910437879b67cf4e9fde5cd789a9cf96522221e8d81df9f546c4096191cd46a4d558789037b8a5c541da328249eb13fd4fb0bd35a984d18b26f8d6035662289a0ff45e34d1e13d02256919e1c0a32a1d5c6a6f9b0722d04731fac6bb38b7a72040c5e3d19fb699f3a11ab86297e0e4b8a764418d370e90eb8f80bbe34aa13854cbd420b6506bbfa4314d2b0cd43f130990c913928864b7ff13b9ae90e1a846ed693fb9231ed2f1dce49c337fcda0828cbee30e30f770d5c71d895cf9fa882c1a35aef21aafcb889c3d19592691fdd350de086321bceb68ca64d32260a9da1715873ab783e74b9f55c9d204eed67195690822317c2e74ef4c2bb87b6fc9cc77047c14a3b8b30a3dd023df9f2658ce98626d6244ffbb79f740500c12efe4d09ad198e87a0b21840cce6c90dd34266516af0d085462da076e47b30780cdf63680f40cb4fe2aae9a8141b311c648728e10cea96f2af61d17d196f4df7a5b52babfcfe5ef97ab729494ca56689cd9e57204bef8fbf36f09b8ecd5bfb664c1c818369e12d5bace7bef7a1287739b687fc8db1aaa4cb1581e7920c36151e26c4bf7798880bf8a9d122bdfc94d820d2c7cc8458412c40625c4f8eb2deed4d9e32f0095224b45befe734e64babb4a2f90e5780e8c4cc574415be5b3fbc39f1983b505dcfdf89c0611522654f864a1fb4a7991d8bba6a71fa7b2fd0a9711c1dca6234f3daa429963562692f229908e30efed795cdf4684443c65343c639a122f2c916a905715d7ac25647236863f34881e24f1b42e0f009d65978048077a9395878a70e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hed8519968ae4d691a76ed96a7475c03d2152959070614618045acbcc438179dc7bd8116ab24b26885e64800a0e41626e5f934cd78ff6ef393729cfbd8869c052afefb1f3f7262a231cea0a3b036dc8d7be4e9bd832d1ac51c5292af45c3afd606bb7f8277dbf8c4af69105a850376b7d8a41f6c3e7269d3251c5383a3558c4cf563c52cec711ba5b12fdfc90e9f4f70e25eb5d0fc652246b3def44beba19147dea0ae9c9d824e8e42600ad9133aff40479494f58f285efcbdd849beb288de08ba6d480af716bd24582005a35ab9e70019976844b9c97604ea640a78952d26524f364e015bcfebf978e138bb8cff2f2c9b40c506e59f6dbbb51eda0742ab0a392ef01c2c8a52bcf8cc651aa0fb3f2c9d4df827699114b78a38ad5409c55b2a493fc59a08d1d00dcdba1098c79c404f1536aee8778d76ebb532c715e8bc2e6108010450e5c36e479b8518cf14995e01b8eaf8c3932cde6f03f726566f51fd0df974a11868de0f1a2e29dbc1b09ab0ae15e112b69fbe603cfcc9098621c118dda00be6168a7cc641e00ae346de5b2020f20d47b5884a55d990e63e8af4a9d0c95cbf3a7406e3748fb759e46c1973650ca35c82f014a7bd38eb06943784281c56bc5a838bb0f9d00673c4c1a7365acadbf3c47a71efbe57d13b208c08eb7eab7619ba86fcb943491ae7f5faec2b9efc364e88e286e083db10f9626ec46b0134aed316a1877fa8b8862d9fa9b1ca41bfb17b232ad3861a0a71a1519a25444e96422ee08f2b36479322fd879723cb5f6623ad6681d66d5c09f1ef198b04627ea7774d26a6ed5de4d42212d6cffd6f629890acb7d578876e69040aab7caa32c955901cef0965f6c599c72be53201768124332bb378f66052f74c056bf2e8ea272b3a7d53fd84d98fde3c459def45d0da2c093695f71adfb956f66377a952c33cfe7d619d79417607a74614912d85b4fe8df1bafb75594e54b77bb980ce4887a5fddf8e5262aca1d43b7a297b8ccabd1fbbf8e0036defa15fc9c7d12a86f162ed41d0ccab57dfc28144b9eabcd96b4185e65ae9c696dde3aacaa0d964b8964a12847e24f7212d128b5e50ad72fef71dfd0ad810ae6b8b165b93a4cb555d1238805c792be28c0bbd5af02ad4bb5445c48ebf7ddca57940ae17eb7e5318aa7471d06fe692cefa8d6c6a8e43bdb06ff54295647ee7268c248138ce5bbc758eb86c878030c62081dff7d30d7f59dbfb8ddb142e24ab2c87333a2e331ee7006ceb9064923325c4773b59b00a554a007a3ba2368262804cc2af109d9c8b83425caf5c1ce35af0d7196cbfd96ed85fcd9e9191dce88276d7d3fc88f700600e8cd32787ebfca4f57753bd4d58d43262a37fb3765;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb44aba9226a83fb5842f73f208c1ebcd4b608189b7db290d68f39e4dec6e48c917cf8fe095ce77f7999497449fbde670bac5d563c9a44625a61fce6bb4db079e45f0ab198abca0b3645a0926138900255567049b00cb74e4b563387695057fb3da43e6f8130d33f7438891941fa63a547b40eed0713f5cc30f7f3f42453707b43a1f59688f4a8859cf2f4b95d84758d1625b05fc6bcdbd20a9e52b250ef8d2e47233484f85934caa025b864586deb824cc101aeb88e53748e415d8244490deb11c512ac219f3d9e051825df1f4accef5987b9bac3a9fa29cea2742fe170a2ee5d329df146d5b2ae57e78a9a6ca8b87a3ffa9ea883c283d614297a9dee34d074a31ea225919d8955411a3554ee89681d54b27cf017023bd071024c716c805f5600699e594193c8d0d8ded18569e06422bca16368757f2985d88d255b3a5bbf9e000fbe5677af982af6d66ad8db53e53a269f356f05e48867e73847a245f2b195d0c89f8551b63a6aa5fa07d6de9d820aa42c10965b42e97208b1ecdf5c1283d15904f28ce8b2f1b83dfad59fbe6edb9baaa258124e93549396a025ccd566c370216d4ceadd462c8d8dc2c255e18afb2310dc26851932e2e762f4e65778dde4c2d84082f70b1fa10b0448e0a1a7969d2d3d13ee69b8740b6dee3dacee264a6091c0f5e444d00fc9b74a760b015bb6d753a01bb7b2de6a1cd3754c89d081c439624490f2af3ac5e5e47ba06de1706ceefbfd0eddf682fb3d18070a1600e3f8d237c98166cfbb216400612bf974da8edc8729c11550d76adb1691133f7296cd837eeadd2d47e4102c84c780677e8dcdf0532144b32d7f9215b6bf3495c9dc003bece299068a5b2740c89a952b0d7ffdcc38e84571459098557bb51afda99ccd088f271e893682b9bda4b4d15bdbd54f3fa545a2e94a60b213e8c423ff70f1368d288005793c37556b302f1c75412840bc84b69729ecca2fa60103198b00dcbbcedcc4ec5521c833997cb9a140b505a4fa6f4ef7bceedd8604b009732a67269647ffb908079da4baf950993b9456fc529ba226203a8e41f7021d608d931fa239ba649af6aee057204f84ce462d4b250b75645215c2d88a8eaee7a31299e3d14acd2bfa1337cf1379b4090ca6b2905d75ae44622601964e76fb60762f41e8d3b9b5c95b762966ab7e4b1d8ae26ae8ee9d26581d531321b6affcf6d326134603323265187e8bcd98dcc9a70739437130ac22b4c66285340d1ba65c0cc341184246d18a63283009f64c3707410d409f7469f87bc2deae4803e9cf5dd494f27d3f30f28fc01bb8e7cd843108a47e9a7a4d5a0fcd570c58d1ea8a8bf75d25043affb214d0e82fff7a215934ac6197e8b51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h27a3cf5654ee2c9040f173edb63c418b4b28b95e3f8b9016e65e7c6ce0c46acf759ebf8431355af46ec7b38891e736bb784f2596f876c04d39b1acede07f85013549b14cd72dfa097dba2b3c4a993944719336f880e4637d73527651b68032955b2f2adb2b1a819b57e2f81d27dcd8fcfca563612c25ef203dc0e285048ee4e4df829f4bc85005bc78b268cbeda714da80c244661f7502e685411dfdebe6f2532ee81df7fa6de00c8efa8c4b83e94fceec990550821a9adef0e4279e11577b9e7516f4546038519b351c0c6ad7a38f8813ad1e6fd9fe8d69c2757171e647a9aac2a1dbe291bbea9cc5757050a993ded502dbb812d822d1be515cb97b96985c6f088b641258f9b03479a6e3f0f437e285c714b2a99cb1100bb646c353b6383a26c8dc926006c0b061f4b350a4934c25f6111edabcdb70f6e3d16eb9fafda3192af8d5d71c75b2619c0ad66b884c680af507ace99ae01458e701ea7937e475b69d935e23323c33ae1fcaaae351d4e952a5341826f99ff6183c91f112b596a34278e0a95343b7c868f7f8d8f444ec362c3cfcef83e1ce9d400bd07a34548f64abfec79302570963fa6b623faf501f6b1a0f81eb48d43769041c8609281613bf68ce4e437ea06d20e81cd6b103f4f25fe704dc78eb3318c6c13bc316747de39651b8324d71a74408261a1f5eef8f576a75525c94579a0b1974c9685ee547559fa6ee0e5dd3d7b2959beeeed8b3ff665066d92eb115bb1d83cf307395dc502e7db870a57e5a044e181a20714714835d62b20526c2e98390e82c0a7c3a087c663de8bd7212b0e49ae7a2000bf7b007bd7cb3aaab7d0092e4685edd3fed95de0770ae2b074f947e70fc8e191b0ae35d809cccaae9d6df974a82c5015d6898be511f6db320ef4ce979316b572e8b7aa2c8ef0c139aa2fcf68fe90d367584473ff03c1dc775c258c80dfa6a9e8bf40d739fe14ab6d2f6980e47ddce4ec996904f4caec1d3d4d7b649c400238857625b5ec0ccab1bf8d9eac7aaf215ce5653597139a43e678eb7d44209d22e5c7d47c5c9b0ee89220da1a8ea42a1690e936fd9de68bf98b3e3140944b18f00dda9c1ab9e85b48571218b2cb7892025a0c75d950af957d92258898bb088bedb13dcc2bba04d01036e7b3373cc430013d7d1db6b9f155ece63090b2a4be0a689384cdbfcdd116d2a1742e86c8125b208245d69a889192a89a450dffb169e54081f8ddc1e56dbc40c9a5cb58e7a75b69331fe6f5744ca25b480c0d1c9973682286fb1ddfc47960f3bb017cef0ece6198f48e487790083204608417015f51889365f7b0dd005b9b6d219e5f71e7c5ed43cbda8fda4039824499c335519a73fd76a1bdf637d25;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h49511fe2e04a15bc45d1cbab8c387cc827956f78c3903994e4cd82c91d7ec31760cb77a936d4e3c35aeb49b7ffbc0083c6a9958fed4ec5a1162b2939a3edc20ea3dec1b780c19a473bdbaa56092ef3f920fc7fdb320b942aca4bf1e3a88af45c7d660e76221404ab3bca8b32c904242ec9c07538d75685e02e41e71508afe624240262de18252eb4c54bc0167d9ae78031669f8d3665154c86eda730aebfa92631f85f1b907d1fd936f0da4caf69daa6f8cebf4ea5e612efc74d42abb1d04c23c9fd3d1f5b8341b9a755a60bef97392659643f7a471ddd9d2ac66871c10fe650d87087177747615751e40899ebbd1615708960736b8d1b66abedf75ea2462265053b273839e2d5ededd9fa8ca253091175be18955c066e9caba39128ebf3fc465c86840bc01f315f979d4907b5a7aac79cf9a54ea5d580cf6f4ab9292e67f4a29776c5100f30b85ba5897f8f5a2f2328286c8571b802997f1153adc56c364d483297e6a4e788c21231abf71b446f1083b1804950a6544aae2585b55ad3a1ef50e87e862204fb1a1a7227fb386e2cf1509a0337e3a2637031cc9f3088bf1159617a169e7b5053d05a4c826c3bb44b0aef4bc93fc664a2ea47a5fb4534e86f0d31b54508d795b9d82d7c962fd32cfcc00ddce08457e661aee8e40f995026332a3806adf47671c75c1e9c764930e3998543b0600d71980cb7f652675e764676dd1738a96895b55d9f2effa41651356d506a0fd600d78daa391868bc3ed2742180f4378079c141bbf178fcc584668ade412ea5fafe8a871f6d82c5315d84c6ac7ad4f11b3a539684e74dc96d7ec57625a2e6d08f8a61794f95f299db2d4fd7170c1f6a7a26aa595245c60b431b870f7568737cc722dd9863011e1263f0740c00a84aa086e138c893c3c161d88af7166c2d4d89596b3cec8c9622fe0ab11b2ab8034557ad62977fbe9b1c81749037c9cba77a722893744fc1ade0bbbd8d964c7f25cd3618d7c44150e10647074a5f7be461ef9fac39004e219c7ab921e15509adb99e31c4bcaec72097a183a57f30835266b6972fe01fc382218af5f9bd99d7c78f2510b1badbd72330f1207c9a7eb7acde852a216d27ff3f03f170b06eabea7037f58ccdbdbb20b53afc480ecc05600cb6aeeeffbca4ff06e1e7a7ce09dae7a1a6184917beaf0fcfa079a36ee646690440d2a312350ba41bbd7e35f6d87c43951f3d3727b5dd2af4643d0949b14c442ffe7396a81a908ad7da9d2431c9c65ba120993c5571ec68728c5e8a930b018cf55c7fa23daea0b8f443d5cc09099ee997f130b7cff6f1c661b6f335975d4ba47afdd77890e9cf5d736b9350729295d728f717fbaae336befff919221709b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6b0a77a3f28b93e4116cab1a6999284ad68ac9b744bcde7de29113cc3086f2d75d2f2ca091d2fa3c82fbaad4478088249e20bdd9034465f17961a3f32b54a970cd4f92fdd2e06fd1f5ca85066581f4b03df2f2f520be64c306492b721df5573c515e11e52958f3240d97e6173536aac084418968e99033a79616a8580b29c39f53544b8dac9b8cbacd01108e69cd1ddde6852f34c1411d2d60fb230a606882feb8c6707ad1376c95edb3cb4fff0f6989de40246b932740f035e1fe745ed34403da3ccb074388d90b02463638d4f9d87f1959c87c4ae4342c3e56c2131d6ecb5b34e2beb6ff523431534d94ca89494cd5a3968e977cae197ce4d9ac1dda7957812c9ee50b56efb09298fc95b1303d34d04c56904123f00216fa5f43cf78918b50a91fd4ce126701d65437800a075bb203b00086dca324930c94dc7416621f4e0b56082101bb614237e12541d0efb2598fe074e924b393907513edfa0101631a37744eeda401b42756aebf69d030d851873e7e2be8b9fbb341fd1fa953341ef2e591480d40ea71458c38fec59f524c949d6ad49965230f74692a6ae8611602660fb084dda7aaeec3ca8e8a1325c2ad73e4fd787d1a0987eff2be86e20f7d9b7b25c57d1167bd3a2950dd50ce2b7482dfaa75455097268ae880cbe69840ad69aee70623850c0b0654a894ea8f613c61ab593c3757dbd10a6434519cb8a0173f25e28041e3b4fa0bfadf56906763ccadaeafb8a54a8a137e546370e2e065eefe03e830fbfbf8431fee1b113d62c2a19ef183f368c878e57b3c8d3fd19f7b3b74c3dbaa71c26344fcaae2600a6d503930bf5122cb7692fc4679f093c82154859ae7e5b3e6f6c4de05c77e82676ab598b0137c3ff0980924fd98b239c2a5511c52104663b836e15288fc2ef2d9ceda8eaf210234db5f693b925336296686ae90d26181d4872f82880e6950eab89c46e7b8548e8424fef4c34041dc6600ee45e5c5f60f7373c596801a9b57153bb28547d1d30720bd0172e08e2a4508273f8097ef64e313655359d623214efb6f90cf99bbaa0006b4253017d7bdd3570b2e1ad65fb59e51899da83779a9dd8d3381f74352135f45e58cc1312f10c8d731ad6a369245b9daf4eac62dfd95bb6b1650bd7f9cf8a86d4c0ae95951f7230a1e891899b295e968efc1b1ad3314cac6a3328783c556b2384abb7e423c732c1c6b1912de53036bbfb585bae5b0c01727db1bf9945e1d7c35bb40681999cf69f251f1e2fd411e0c42330eb5bc4ba63330f4d2b5e0e2002706f0e3974313d2d6255b5eda0b86d91a1b319547f9eb1d0a6657b05ad34dbb2191e66148b193bd5b40af6c12cc99fa4dfb762ad283b32a2dd80ea4bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h991c4d83fcd6cf81d15bc7abbbbe6fe2913efaae443e234e088e1289655029c529536b8c4096c2c9baeec3eb1372e5797ff1d5d040c7b02a48112b66d74fa506565ece6807b07f976acef8bc138d8780abd711c7b3c5e25b0ed3cbacfe29d794ec731586feca0495d1024bba08881401f25e51f1b6de4bd3df38642e2c7d20f17cfd35e6128443b172fb196e1f8f2a6bce538189feb9f8585a78a17a473443983836f1a56db7b637971b25d48ff30ec1e09be5a06e6a711ef7de8f4dfca93039056795ff7164dbe772ac050a5b721bf75c2bfe5c3a005ab6c9484f1a68d12dfa318baba51d4e4eeaa5ad4a26e6b5b8fe96a853d76429f0e61be82415c3c8fb7deb6ec2d1e7d7fe7046f6557c4c2d9e68076367c69ada4fd1df03a28f3521f89a15a07a9043bb4d95d6658f395765f7ce432a828d32632084270fd9a8998ab989848db3d0453df320a1204f68ddaacda29f0b61e8d1d331742b21f4361f907f10e9c2dd35600b45b7c229bb2d144a98cee7736528dff0a2bef2eb1cc268e7f356687bdc786d1d82c5e329ef50af3ff3c15e80daae7d6ced574fd100c2c4c3598723e266b92714e29c090ae7aa1b31892d3692cf11d6fd0a5e386ec73151ccb2860f841e48cdc32aa88c2beee00fba633abc4bbbe385d3eb15f9a9e5dcfa28f164d109ee2ca0000504d66bb7c3ce52d2134d75cb1db9bbb7a5485368e68297e3a2e9a5b35be70ba9b4eec69844394ac32f88d5826568c318b7dfb8e622978ca0e81aef8b4359fcf99639a3571cbf15ae24d9f7b11ff7a3ece21c1224a6a93ca43be3951698f8620f5e81e50a795c13f2d51403011836c05375fc1f85301418f3e1041dc3caf9679e6dfe2b5d33892400d7dacf00723745e9bb8ecf92a33bd122e4af90f69bb79c695a12eca76d7f11b3601ce752f94d761d11bf55b2cd5173d03c9bc7166a878fdbc5a04e13fed3ea61408d51afe9612130a52d7e9c1ed218706245cb89e46e132d3d8a16ed1383af402f5c14a33181c817c622618cab3b9554d6ec65177e6f49a785e0d33eb8a68d81db9da9c9ab29f39c1cfe374cf9747b664c2d92912da68bb89009ef64928bd20d902b6ebaa1fe2cb92deafc49d900a6099d3a716cc24191da927b7245bace28c3f3cad9ac7902eae9d3aa3ad16a20194a6779472cc9d6bf83c1808981be84514643ec04801058c05e9100ef192894e333b116889615387d9afae3ad86055925bdfbaec152afe3fbd3dc9ffcea2264421da3d24b2e1ebe67660c3b3fc7059913fe7e018137cd897b64a8cf3c0fe0127a7abaaa460e2a118283a8c7e2870d314a35f50211a16b45327123dc3c802ca590453fd6fd8f4cd43c81fdd7ab99aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd6d2592a39decad06b47c4006c4578414184d79fc7473752dd6ecf782f489643a8a40f731024d5883c99c008abb84a99122a590cbe928b9687fb49532676efab5951b321b9dfd0a4d589206957fb4a1557ea1a5fda5c2b850cde6db9514aec61e92280b9d2d463aa67d19e5e3a2cd6a4408578902e595d55b0e0d64a906546c0910c0e4512608fbfbf7900ccb41d7135afd4136f3845d2d443e3729ddbc2d44ae1bc6a4eff38ad7159710493ee5fcf480dab3db90b179e4d895854815e164fa8fd81254b0267e1809df30ec653ebc32061263f3f532cb1d829b9180b474b4fda3aa3bcb96aa05165687b45850c4ede9c7525a4389fe08debdc80066c8915752c316f0206dde4246b9516c9d0e426ccdd6842c0150ef98eb5b2c5f5fcc31798cb1e8128ec0ea1fc63b4249af39bb278bfa41f23b587bb816ca84fbaee4157bdbe11939d1db2c33451a769ee2280c2cc362f4f770c54f241682475e53d0f542da14213f5b1b22ff02f16bb214ce38a184fc15c3ec6cb32f95e0516c8d084033bad0d0878dd3a55156331d3f6ea77c8fff520c59cc9f27c346d5470600a56f8791c45bef5ee82a0ec2ac2ef2d6740642a28a60a719d183b64e8b9b111304c5ccbc04390a7e8b18c5c0b5b4c02a04e8eb00d11af7b0812133a87e279a029fcb03795e689c2ea36104ddefbea4313676eb3e31cd860ed01cfe666bb7d248ced13083e0600666528d3556f8254dd19c7aa61f83d97c847f629c82ce9052afe4edcfae168643249a666551a14165d5b5c58624dae7bcc977993864bd219e11ab4d82b2fbf99a912d88383f8f0163559556fa062389d025e3a20fe2a3a19352bfeccf9875f9ae21a583da609996f64b0448678a021b88c64010b58909979fdf15a78521a87173e100be2859d7c0d09a1c1261b2991e7db28074b3d8fed172f0ae648609c36b851b4af576370bb884f541dcec258ae2fe4261a97bedf5e2bdb6ac36f1db63cc627ea552c63000abfead534a7031f9b2445b0d24c6046c5fdeb9ff4b92e4607eeba85750825a846ac86992eb0a8b5d1a827c4acec13e9e161ddf77483385744ef87cee897bd866f70de532931555290a28bc75df57609130a328ecf1a360df91680ba48b940d1d02fd5013d6ffb0a2d5322f0ceb67b7b180554f36ab8d6427ca4d09ff2d483c4a3081de41b41a82e5c6b8a6c302f14c7e56b9912b07b043543b902ada09a91e2bcb630e52b55f7167a40e8b5fd0a52cefd54585d3913051250117f7ca24e3a7c253cfdd089edb24795626b9c0d4f17ec2ee2daee7fc8cdfee0bb6c7c3da8f429897ea30051651600554b2d6cf9e0f9f8ad6925041d10b245206d1b3918ff80eb8febae9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5c548c23cc19a89a28988eefce62c99a61fd942397f7a1ce596c35f6daac16ccd8823471a61112267806fc9c3fc5f55adcf8de3d22db2a2e0368ef114da4f4036f2013c35ecd8b0ba25fe4631bee65360c3d81d953dc8d602002317f5b3aa72c2da604f0410b266789d7dcea50baff6b4f238ced67f99e9845a2a37ca977c87cbae0e7f7e2c9d4039a74f994a60d783ecfe22a4e514dd0e8827065f127d95c980af034b4328f8ad03e79cf9d041584e446c59db565aa26c1468831bbb5a439c21be9e5fa4ff24340482ca78e4aa99ffe9ee266ff9c8d2dd0ca83e81ccb65b40642211b1b3dc720348c913582b3a1405ad8358c60b66f82bc1fc724e361e0dbd52efa3a49597b7d93efe8021849914fed1b4c403cc801cbd18c6c5fb59b2f305cf5d02f458ab42df0471698bf6bbd25f36c2b00ee6b199a7fa4b2af2fd0b638613e5306b00e6e09dd34441878339b0684f4ea71b7a9fafc7d12fe34a5442cfbe84b45610f0d885521a72d378ac6711203bf5a4451d9f6ee5919eb3803408ab70843f98b0732c35e1d3d05f10d3c825babb38495f41d06f2a99b3dae255b841cd9cbda1e6fed231fc4f7f252e8445b269de5fc31d2055b41376b038238410d2b7f3bce84487de23fad1eeafa2c5806f462ed4c9baf072f854ff0274bdf09efaad84e2b42ca8790bc0d568576fa561d9e4ec450c6fee87cdb5763defaac96fb5bd89d927d5b67f390742478760063c574bb0b7439135afc078563c106ca954613df5ea20d97b0871f558125e17b75f1a672e040d28b586c0a6c508891b0961b1afbbd84f64ce467d0f682fb4152cfa61effc212c1add0a939a41714680fb9ab3b4dad83799316b7ad898dee14ed1b4833433f5b4bdfea6fc3560eda7264a1053b80c7116474734f75b2884b54892169d30c1d62d46149352673ae2287988783fe01a51b59f18fb599a8152056ec187be6a040f7acf350d33b6192ccc6b53956edbd2b9612876006c6372ef76464a6b4d5a3d743890a7265c98536a9c2909a6a4cdfb9ff2e92b8af125f36519cda92ee05dd92f7be999d43f27c95543298fd18de6358e1e7ed2ed027b32ff472f7e890c4ea925a4b1e4249d339c455cfd4f6f8aee859e367884b048644679d571bbb8677d91275a0f5a44a6ab5f4c2fe6af30301f6f1538ded9a9185b932f21dcad70648ba8fc10ce9dd3e54aad4b389e988ae0de46a9a1a43f724665d983313b3a8afc476effd9806ef765b2c11ee4a226a5d9c536ba6428980f2eda0d961b1388b754ee7d06fc032b17c872217bbdb1fc17724b13e73c5d7114d8ffb94caa94d78a4930b12c4956d8c615def673d7664906d6bb06b5ebe43c733e0253b5c1966;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha8789a18206d6b3f0a6032fef7e930326f5a1c1211545c143a20179a99326e331a1340c799dcb613e294bda9b9051fec2f942a93f590cf6be9b0f6f5935dbd5e23e7f865ac8b62a36d6659464648f9a7fa0c6548b241e2491c941bffe383bf5a61b93b4b5d391afc9d5126046fe78ffc034362824e3aa42cc97e6ee005ad800e5ed39dd9dcb5c0e2dfd5065f6b695e3c75e174e08426d800e7eeb598869dc6a8b181a73db423223c0542e9d925e1ca1334b1b9bb0c2204982b7d67da83c192ddf8230d9d48f0db4c8e37ebc9dc46ef01e0f68905ead8961ebfda16ed770636f203da6faa1b95339e71041123460727cc9e4d9d3442c047ca54d2126c0a8c289c69c95cfc0e3a7778e6dbddb5dac3333013ba47d25d6f7e8735391656337a96d27632c425583417c5880cfbf737544860c0c163344be73baff3c32eb14445276e1b90acd579e1432738ad4804ce0975842e61f830aa453e2c1827a81ea449f37116fe164a57513b10ebe5f05a5fd5e10001f12f3705a6d9a657ccc79ca1a9460b50f4a53e50d2a3b921d00f534c0633074535ae43c688ecb0650acc811c0da5b61a0303ead2a4532f8c6a833363fc6c05d1de499255f73a18fc18b278ba4c611d114337f5bb6317582bdba47211250f99b891b3ee148178d9cb53420362fcb2fd163be36db211ec0b53b4c4ac08277c651aee3953770c255154c556ad948ded1c1b2c51cf54e34e9acdd5093c1f3d1a55c5f2f7d96f1cddbf79063bdfba401a3b356c536057d72b8623f96a6c69aefd895fc7a506ff084904d622b348f61f293422868003670ebfb2487dd0a5eb556739a3c58d987eed33a1f5567b0b6c80819314bf1d36cb24a7b5e686cbdef21e8868aefb73f9632a11825093060c216b1c11b7efa99a5cf9ba716b3ad4ba424d1fdbd8b7f15c2c16780f2db06e7e0d547b30db1a42c1c945b39584a004fa7fecf5934cf702ab071e394b128a8aa40a86941a2b61a76831ea3a0c657ee80436a4151c2522893ef594ada0d42ed348b395a0ece75c32fdb6e0f0a58c0b0a49a2d87eae90e306fa1bfd6f881cbb35c5384c9785d3019a4cf5cb8e85c6f8f841fd28926cea5bc7e2030bbefa5d48f49d9c69b17a8047a4f32f7e4d0117a8f6f6e63ff1b43be977a294ac90f5db9f4f8a7d1b528f85e3f89379451dca62c099f880ce486bd3067394f8be838ee2edfafc5fc7368d3af5d712863f3c65465042a19e58457f2afac8f5da0a0137d0825a22de156aaacae4dfac1d65b591e94d9177ab61bbf50651629883a92e0d1aa2e786e23a7127edc1f0f50612fd41a9a43891d5635457e69282f301defede141eb04d399f99cd22c040c3c277799c4eed8bed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h54cee47b998d24e1bd4debecbe92751a9691f5d280b0510ac5a3b6baa13088489920bfdeb063cfd8b8146198903d088de8923d7af5a091c808f26fa583f4f610a83dceca6c232fd7cdcf9b2f2880a7553c3f93be95899a948c48a93d187b593572c4e2b2693df2304ebc877328dddfb1251d454925b2a5422f6903e20d6cc6dcab0ee4828106bc8c3430ce2d682ea8d09c71c404f82b950117b43203988926a690a69ff886b329d4314d757df829648effbb17b70b6443593baba95ba960ef1c623e989f537da6950d4b9b5f24abab18dfde343acf7a42e0b9544d2235299b9bb9bbe9772798279c7cf792f5d064797357c7326d15d1b668ae3ad6c89637360ea1701e104be5102af0d986c22024bdea26f746ff0f88dc40aee51970458dfb56190b187bd1aa35dbfeb1029506d9acfaaacdd5723fd26cc418f954bc5a1e7851dd6e64adf8a51fc35d8212098756f0d372b1eb2345459880d1d09562ae484e4b10e3599bcd9a56ac601e79223590717ad5f1a9862626d3a69f210f72ad3ddb0a18c3e3a6e5c987907d2da436b1b875ef1a681eb87a55c371717ae8427ff76ae38f8083dcaee1b18a62f8841744c2cd7d0e52052e7e64bf95495c6e73d0ea3718541f3075a5b3ff60786bcae038e976adf5a8f89c7d09bbb1a4dd42c9b6c942e90fbb48f02cd0ed2eb0c20460529b8abac5e8b31aed88504fa895e4df06332cdd07210b1ecd37d290c2a095a3bbef5052ee48e99be66200206b068de72b5f3021adde023dc70630ffc5de2311875dd3bb3fceda1db21f76ffd21b00849d9d09ea2ae5f96c01619975966d467dbcd7f7b37960d96c2c37c864a64f8a0b3d93e55849268421a8415fe42d13651042dd176f77a488aa8c833bc5016727e7860e29ef61d46e3c8a60b4a196338238c0dcdbd01d6f567d2f98223c3b177dfca56a8129dfffbba7238c9d426b6b90399902ad4b5d0c60fea58d18c94882aa522f6d22666716210ffa93844ca675d3b6179def52380a26daded977b6e94ccbf9a45519f8fd6b70f40c18cc641f382cde64eacb9b3b017848723f0178300970e2cdd39f6e0fdbf24718e707f466fe2fc8cabd7b1c9960a10f2a18a27f3492a9bf455203436b836912d9e6a6c12545e0f98b1406cfccd53b31238a491525d6b97a6a015b100ffbf18177e6aa244a01042e30b260a6ef47f04cddf6d36b3bd14a1772f57edfcd95839e57ffe42d1fea2bce9d5f51edd8f97749b1af17007debc312382ef935d65f53acc591b47ee008d705b46e845b1e4962d364e02197101be5029bc30733d579633c101c210d4dd4b3b555b641f10689e4559911949935c053b2cf2b140024fa6134ad8937ec90c0ff27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1556530176b9a6652693c2cab605af287437186bbd1167991ef582b20faa849e543859e8eedea7428ccfe002472fa2093685afd93720f85f21a29544c72740692c905296b5918fa91f1ba4c3b9f46de748340dd93eb97df73dec07721650504a9ccbc1e6aae3c207dbaa483d4f1d38e6490e559904b0ba997b1ed0c909ac53087ab2c1efcd158584381af86ae972e09b9b444bf3375fb9b774f0201d0b6558803143e22c6c85e2af194cb9ff34921c946189f2c3caa08ed8b6899e20b752debe644c1305dd8db7e39029ef4c0e03faaa51d9db37acf181bd96825a76b67a351ec108b1ce9da72fa2a0983f1967e375b5949dc8a12bd9209b3ed57a2a474b8bf5fc37d319051145b99ea2fd14264bb931518503c24b5ae11d7a7da209d3ec2e27827ae16bfb82249bf57760e7d5d104d600f768fb4eab5429fd562b0ab54866850a6423988c681a50523359a2408fb1c8192f2944a610f55ecac82d9ddb74ba2c2efb9558dce22a7ab5358eb0aec1b6488dc9f07c5ed3364c4d55a9e8195b5e4755b0a60debc096443520d8e17fe2071738693585b73232f31e8344a78ebf8de289907f5babdf4bfc26fc7d73e46a796e84d9bb6cdf0ea93b9e23cff1528d72c54770145161f5e7657c7a2ad6d01a6160b034952843d54959907a0dfc2a7cf869c6e62dfb7817853bdeb0645c7aaad72f745b762bff34102388f95c0fffd08e3cab776e5a8c7cc4f16bb9e50442ba353de19741d85210f335254b99fab6f9dd516dc623472ddd7e7397d792d243a0ce647851955488ddf7f297329e3a3d48a68e25f61472b79e605deb24cb17d60a6f2b1f16a8055e15b254840a7e33d05487ab2d18c963c0237510dca152f35c527c9e89d7b44b393dcc358fd729fa8718016c247d09f4730f0c02ea37c50ab635dc0580c6c24f153b9b3801d4b63c19585ea38a2801d17a52b3c2e169499c969179af7497253fafe2e889496e0c0c78fb7efa0b77e25a7238f28814225c41b4afe40429ff342f080bc5928107bd5597412c772e2a92cff6b17889b6b83a49ef4c98144cded843e73d0f179422f0b886cab8919ef2011be243d5b539081edd76431d387b3a1f0bd1432933dd3566c81ada0f30abd4d0a671ea3f3c716f578b21abb6a5ebff745db5d4db9876316d0d8e744cc34e637ca4f5c9e712c5df10b83ec44922106b3cba7feec443fc959308c33a9bcbe52d074307fd36216355eccd1289cb9e1f768a44d86f608fd0a25decbe2eb88b0894f4d61b9995ede45dfdb5b4841e343af3ea77f2464166358df7fa8d2c19e18b202524118bacca7dbb78542bf284794dbf8fef3ab1f74cef85e7e4160b994419ab9e36d9569843773e95cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3f6571db7cc1818c12e439aa6dcc2e685098d990914eec7cfeba743a8a8aea74e4128741b7d41cf32afad28fb57881665334658aad155364a6c4934729f7761f7bb7f9fbad00c41c8e48dd6cef79fae47e327a45fb6674833111b9dfbdd47d205eb1753d8b292bccc6ae5d3ecd7c142bc207a1316573fa76a0fe4361c5d5ad78363aa70d7e2e1e056d3975bc1a09d45e4a6e79dd46fe30a1bc6164aa88a9178e710fde9534b9b3a9db4fc4e1321c5e0458ab68fd1fb4c19eece2fd44993d0d2978b2098e73b40c46f4d303def6c77236d5c5ac78cf88d0c17259796814fc3ddcd48282050fa1f81e1e2021b2434b83a642691aba71b34c4c7c4313796f0504affe876744ed11a1d4f26b23d145918b4da99374b0989087d6c5e20f3f9ec4ec768474c0c5f78d7106399ba15dc94af1fbe1c591f1db85754de0b649e7310dd6af168334bca1bd899c334609a06f260a79f764c6dbfd6b9951e4e8a462cba74f2bfca669ee0de076e29385d00ce6bbd421b2f5818873734261ddb92a3d7379cc8955bcf51976cac5a4684cda87c054d70e15dead8f8b10bff16907aa6d32b5b318e9db653c6aeb3a1aa94aa91684d9a342b666a44b20fde5eda02f0b911def724e9512fa0631bf0b64f763200ecd0c41b97dbe092b363ee8ae6bc1816fbf0271afbe7ab9c706c809cd8bd17fbbde214e1267b4fe4d09382110a93bbe9afa889b4e8b60a2b6758dbebe7df00b2a844f1ac092bef2e136b53320853ee5961508b7699553e9d468e28f7a9eb61942b3bc892502042bf79c18ea897f86ce14b76f421baa7516cc54fe49c830da6aca0da68f124e63634069c24f6b3da06de5c8a0fa0989916f2d6e69aeadfadc5f248a77c6cd022581855cdc239951e4a5ee54b97c489622124a04c6f82c1f3b9b78c42d2b685630a2bf61ed482fbad02f2d54c26c0ea73188fdcc451c4fb5db130fefe32147bac9b01050b8a0a2c18d755c39e2802eb805662b921e68ca4a4fb2af6f862269e7dc97b95c3c4bd22fbb9ae59911b7edd819c6dd3434113cdbe659b87c792c4f7bdecbc00f50a293731c7bc780cdd3ad766206a6ecb0a1cc5c616f4de7b140ed3bff76ce0ab8d6989147c4b25b60ad53b0b5e2218cc896a1bc2b31d5e5cb8d4c2976a41977f506eed77346fe90f67a57d0bf03e01fafc15842e1b1ede4721efa6f92bcb03c470ba62d38576ac3f02434586dfdf9efe706e980af4ba2015381c1a3edb698236eb2457de624c2a79791851b396fbf1625b8c2e045bee8cdd7798914ed8a1c978c363b5fd690bdf743be20904c799c3d522a2b32c4e41ce03672efa86ba112d6d3a7d81e307392c014b11f52044b40bac212ee5e742827;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc8008db53f2d3f1104619cf5899f5b7221bc07e0e343c8dee79d96401d993288b327a7157b0ec68ed3e317ff59dfef5f41d689f5204e3bec143241a71dac4cfa8b26d945bfe130b17e9e1c972caf3b252fea70f0bc0d7d6588c46e02dfaf4c3d0e540fedf2b65405c7885e2193457f6841e8d7ea4dcfa9a65806ac8a83406ee3808fb00f9a2187c621b2ef4fb6f31c4a8b050f88f430b1585f9d7e3bcfe746c925de655f39ae5be9b8b1dc362d43551d2887329e48b011309127d4e9e1dacc5f5eceda1d59a717c117cef84910836de20bb71dc549bafd5e70da95f296591df61ec8f1f5e52376e6b95bbf8e9f560aa96ab24c2425d3b7702a6c092a08964db01bc2a97c81fd42e783a2da361a11f2c384c776089a903df93df8401b5824c5102e6b643e0a97d8d715cd0afbcba98ac33b982094094adb2635235c8f1265953ded401e563a1b4fe84d43cd09ee593f86957da5f8ce92bd70dee06289457800d38e5e2610c92124914b64718ff5b9000a438759acd16b7d7b181980d0944b5dbaef3896bae0f7a034c49c72b6574c4afb84ae1324073878d2ca26e232e0bdc2a7034631bff2a5dd00d36158ba2503e8b627250ed6cf5c758146f2176d8a9c568afe7b26dd846e1a5e5ce2ab4997474602ad2cd2ea72a1aba3b4f0e33388c41fc59e6de40636b59fdb9d2e38e0e7a7687234758af0c340f95bab3c073bfb8c78f237793da6893f87e747704ef24410fddf3f412245a75ef9f9bb983258fb7c5aa23496ae9a4886065c4508dcee1f32e94d1f28fb68e10fc082b8b2c652628fee41d1eaed35ec90c55b4315a461400da7ccf66c4a6d4aa82edaafb488271814214307620262561af15ff40b3f318735732a737a4d68e46d12e61b51fe527276ac02760b131ed72c4b330f848a161a742a0aadb65e1f27698d8d046c15ecf226ed1201459a5fed9ce16dd109f84aa754620084bef4e55c1eb04817698e4ad832c7c5b3cb404c0b80f633ea2c3ffa16cdb7875c73e05813075b0152fa75174d1205c952529dfb4936e3d60de8cf2513a5057f4c30799842ebfed826c6f11864d86657a9652c3a1f49b9bfc95024f423e71bdb4e3a703e41e59d8d0d87019dc5242cfc5af8e0a2c513bcd17ee1ef75764ba2cd49cd7c23cfa1126609380d1a8c9c66b373dffadec039f33fd5f6cdc2197e6b00e355a7b20d783830319708165210ff01d95765adecb72c8c7ad1d85ba794ff461ddc19fa11703cd7ee319b1388f63bfb02222dd120960a38b1f9fa5211b11c01e4015a1dd6238c7d993c77ae52d3c821a3a1ccebf258dae3230e5ba4b3420148d9ab9f1b5930fee55119a4af6e70a7527e26f1e0fada73105331961f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he1ca251c03d479139ab45e6fe0fdd1c16818dab1d2e9a33a8dda6a8de92a3b44ccf2846ac66945ef49f5b37dc5845ea3b5061d5f60ba6f71b95e6b76c27bc3d98bb95224018daabddff24a1732ef1740cec0ad8756d3bb171febe5aab46e42f2711a767510149f76a2436dd75efaa0d6c3f34a640887eaf43944b9be041604d29abcf21fdd6d5df4388ae398a6a862934e83b67b9a8c81a72e50bde3722405ce0599404f580a055fa029850023c20c959395446a592d6eae0d3d6c957236372b276d00d6413747293f47eb4d7cf768f61b5873fef5be7b2711ff5d6c9a65b2e98d6a6682faddf4a576871b81a86844902c335b3f644c658cbdecb257aac4f13bf00ddc12d412cd973df4505f68d3086d4de6597e4cc2a42463f223895c1b5b932752474b9e3cf717b5512de87e5862bd0750f4cfb1ae849f9d9c822d64d408889cdfed979a4cd9f455d783aec02101e83454766b66edcb404608a8916cf482791684af3b33176a6567b3ec8f2b066f8e1a185efeb4f2fdc089892956dcce00de6647d2b5c11f91000bc506838bbc9b03267b8e62052c9a34f5184e83be45f88f9eee5d4af79d75e7a0b9672787e841ec6db97961cb4574460f713cf033ec9f9c5d6c5af770a0958691be7ad87732ef58d9733d487954d32da9e57b6378e932a546b6d3d6dff76aa2973e39ad2f091c11055c14282272fef884e7410b252126af93026396eb62aebacf04a47519750b52c6a59719999cceffd3eb5f2d53f72ffc921ddba158cf2159c73a704e342fbef9d15c4203e7789b3bee2e2827afca86ea77bfb6baf8a9d10705776bd9937361648fe9abbc19c077fb84c9a7953556cc600ba32182ca6043d03f868328549d802b3e66431ddda8eda4a4f6214b67c2dda01744eeb3aeaf769f66f90029b8308006904bbcd257c5a97b71a47c954b17f56d63a9c53a6d789c2e9c2bf79723fede27046d0dae78f388f0506d87cc7ec6b6c25cbfcb837692a71c5e04ce0208985c717c07f67edee44e847d06ebe6fc47b364e35f6869fc163a4cf5927cc05a93d92033cc31897c61c0bffa8ef1902fa71f3e6d0522f4613de6fb1b6e762491f1b2a7ffd17b3b7069b7bd25ceb947a404b75a6624d4d3c5fdd4e42a67286f56bfb4324d7b0cd9a3e85e11b213b8c62c0eab5b4afb9020edd7ca9f81e3560b0b781dd087c400a1586c51e3c6df40740e6ba7c504a7b703441147ddefe01d80a136c79d01ee4133f2daabbdba27461446a9bc07364a719789ddd2f0e6fb50b30a531a84e7f305e4d416f6929f47666f032b0f6873e953fbcd436a6fbfdcda24a6e8ffd6e26d189eeab4bf1e73608d183c33a1d9f322a171dbea391369e99c0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha8b09fbe1c3fdc71fbfc63274e107752fbd983ab2e804671f297faeb7c5b47011f973821bfa6ad6a4b5c494e692d5ce301c1e2e5d3af5b82b6d0b9e0cf6fb6394ca95e4fe8ca76a24907e928f514178a5682292c76c8422de65629988f377ff8eb680e1e01d750916a75c71e7204ae7746b0cf5aeb159a084d56eca8fbc218adafe8e701bbb52af2b694baf43cfd350e001128e23de3b1b0ffe05e105a8e450acd9454f621de5fba35e5920047fa49313a2955e2d85bde717c30a45516f71cc7d2b616eaeee89f3d7ece4422f3c73d949b683367514be185c4cae41806e6a12601647e5293f572e6176903948413a04e5b22bcee42872d24cb84db6fe702eaedb93e76e50b2f39a0c42ab56a6a57a4913d869b88f7ff3f069bc145a34fa737fd5da39c6aacdbe6888eeb8a681eac748ddf21419ee64a2489b1c57b2c4d48e8485a9108e11a4e5de2f25b0c278e901284e8f25067d4f97193a88602121bcfbc2ec6e6080bc6197ca12648c89fe7c65db8d7bf96b3d579aa32b2f96c8dd18bc05520553e4f2213bd2e38aebc73d3bfdad850df83a4d36df93de4769d077a978a44d6ee6656be345cc418406f15aca4982c1e17c13557e0b3db52ab90386ffd10b5d5d74dda65a0a4c9da4c083942a19196e81471294bd7f6f7df6a31c7ccf5033212de5b87acee58f311c90bbb43eaeba5e315b9687e55bad58a35f1bb0ed8ea53a5bdad1ea1a708b67351723ef09b82741c511f32d24cdc4d23492250f4bfd6d02fa327508a5a87880ec387278704756d949f548a332a257299dee9149549a71a6a916e81c3deaba905be800dcbdab67f0d1c0c1a48ee5d753267e29a631d3d7767032142c50975d3bf08b5f3fe6ef8c25f2086397d67079e4c250fec8855b5b2be8cd8fe6e2d5b51437bbb3363671c4f0dee0ba4ecf36f4c028f4af308c7a86f8be81893cc62d074eb2c499d1d3f3805644e3eb38dda872db6b1451b4970475e52ba1cd0554e5bf2043d65774a85aeae81b1bda81294cecfe274822715decd19f1d0cd45a83460d389d050dce0347a327904c8ec1e69b8def0f5e96200941eb34c5326e7fbe4445e2ddf1e063964cd3ec5e0fc1334c948341f2e2d1123bc6383a74f2f517700a7387a0b697fd1319940d893affc47672f8d666d437c7038b53c7754fc2c86e499f58814b6e0bd4ad2b85cc41935b17dd7199dfe02ef35d9bb30e72f15b1e828451000816341d2994bd50fae4a31a32195e7ca44170e3605678ea681280b5d2d9f0fcc34e81e88b892de486b362b16ed58c9e3366418e6f23f89306220e88372a4a7aa7bf76260a505e539a0735ffba7cf53d6b3dc14115e81f378e33225abf1e13d177c29d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h742448d8569a28cbdd884a82c337a71e2c518eaba37c8098b93af2764e6dc5d2c1ffe55b86a485ee8370f63d521e0710d679897677cae71c353c96ee844473985f2226148ea15f0f60887eb1832afe7f047fee4f0ade6de1cc1f2231f823e1fd3b99f590b24f3e6622f1bcec1b47944347c0d5943ae9c5064d805785f4b8714dfafbf5c1167bd2139ec5a1d0408f06447a676b3a1293b332c52894b39bb27f833a3daf8a06bcf23d240028b819b222a72907a25c095455dc51f73027fa04b2efa3c9209c4eaa5a8e53b9b75c546b1ed0343fb1fc6cb971f53680157b704976a350b0d82effa65ca9194783c656307a0378d14c1f662f240d4d24673d89e519738d8341f7604ddd30ced5f476ea08cde860158cee1c36dcb3e950397f57231a439445c1a2e5cca3b715ded319115485e235e4c23451532f939095465c2784dd07f1ca08b0f38db7dca41bad411c4959075842abfc2d7e3a5b7b6a3766b3fa2bea6e6f7550b19a6d6f8ffbc28aa98a833f4a03e9ae3456e14fab9c13f74e8b89a0fd272b02bef02370a0b7674a6476d2ccac42bd4fc2ddebae94e76f8d3f2e1f186cc6b68fb36ec2bc474e03404c892c55e061fc8bd1d1462951c8caa653eb60d5802477288239851e3d9f2fa6db97ad76d9904344ef8af81787fc625f5e0379c497c97e65ceb793739a6113ff1151f50c130c02b6db63da4634a243f73aaf64414a9fd49269e02c45c9abaf2349d87aeea01eddf91fc09eb6b24febc87979d99f10fcd80a8118eb140c7633f93dba3112811332b4ac072918f106b9cdd74b9e2314e307bbd3d5e20eddc881013a7ee06f5490f1934bc55d37a1d2a1ab6c3f3c2a7936038615d75d8340d8e031e769f37584943ee90c41c509fa8dd24345558d3e3527d2e1297d3d396f5dc424692ce0f898fadbc91112191e80d2873c7dde56f9a7a7079616a12085259b6301bc0823f1a6926436d9feda24535f93a9f8c027744e1df2957e3b4485c2705714027bfc3451b565d84452c864b9f11e9035ba01a4522aef22d7d3e31be647b2af73d6e266c568e44bef8b8ecb85772f6ee8dd653139566c5c6433a8d4e2e155598c65712fb81d49de874a8604dfbaf211e9881fabf6dc33242704bc1b8a85be7234003cc95ec3063cd073d7c137d537cd81bed85713f2cc7f6607a270a50fc8dabfab34bc10ffb0a6daa2c9618dd7e5f9fd115abde8673963c62bbf9004a94e14073f7acde37e3bb2ec45faf31893ca337fc0fcd1ce17ec53841245e6f89dfd6ad9d24b2c1b7058eb39b065f07c9d1d7d3905fbce76584eb270185d4575547e832eb4cc0559cc12de870769f6f2916e382a6478ad6f553498f83b08e378fe536c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8c92f9420be959b6f2bd63558f8ec5e5a7fc565c6d694fed2ff12c6b09d6590b9ff1fa9e07a8355cc3434c07605c6d2d2bf0ca525cd82791e17d3b0d1f458ca4608cc6f30108e692be630a1f6512821839d21987aeeef520b091eabe47e7ddf4eb211c1b1fbdb6939ed9c6ef80c70f6169b18f192be2b67fc868a62f22c2cc9c03f91dd978b73faec1acd9089c18c984241b11261845dd739978c0bc852a99a54e749dc5b67f5970ce8a4c2d007e935d428d3e9a77f91d7dbabc43a88ede2db4f15ce9d134d26ad5a458cacefd25be647f7379a28680b5fa0a9c7f9d8847434204430886d0677cc603661c15f57b4bee8d753f937d87762e886bffe07e31b187fbf7c0fed36edcc58db0ebf98267430e9776feac4ab55b63c77287cc32d3ffe887fdf1bcd8b4a4b28e5b21d466358bf24b62b3ec754c6b1c9d0943c23626beeb38e87f984ebf6676415fb78d9a73b05a6a89c6422901ecc5a29a7a910222f456c88c513752048a567843f83875969f4effb5e00700bf5f6879ee4b991c033ffbed97475a63dfcfdd7eeaec543a76d7069a824e109ffd33cedfad6d3b67932207a0ddf5cf582c77ad7e4ddc7352ffcd27e48d9ad99b15e464bd7e23887da15d7f30bf970ed54ed6be630f3952cd2a3c54f249c8faf4164e3918ee5add3e57e4b1f9c54794ab8979e13ef536e04dd26d3dfb45df13e1df953dd9ac8f377e023c6a34a9fc222a55f785549cf317d3f99df7636b784c2267e39944451f73ce0587d65a19e2d361da5970af4a7bc0c6b2cda683bc40d486a2d496bf3b1dc74b2b92a27b6080f60f86c0a689d4b00557fd089ce734e2f0c100e0cb902a4dbe48a067f27fbdef28fc5e70961994bde1dfab151917a3d8e959b2f5f6eca64e5b9645a638b2f17483867aea9e38bc722a51e903008d50a8b9c00bf2fe33efee753de39e2ceb590da17c3a33bf2e3c6c88b2df04a5536a748e249c8f882fe4d27142ce657567030374281975c3a42f98b5f9056d6e1561c4f7523644296f9c6dbb5e7ad7ce9fd588a89009f39f61a6a12356e12af4bdb707b9eb2c363c3f96e1405f0ff663ec0cce9bad85551ef2b577cf6e915a18cfd1808105fd9aa3f68915e66a6b8e245e93ed254e7b001cfaee17143d4771cf94598049af038af0705952f86a875eae12ba1f8e24b1aca2d85f9f3188110f6a95c8fda7b8e7624168d0a86ed537fda651817382b0d717c7f0b8fe7c10802d87e5e56a208807de482fb6aeac59c1a4c7b145025c28072fd03a1b44816adc98707dcb94229252416eea6a4ecb2f4d7475e0595611fbaf5f871396829662169a6f8d841e85bbd2762f1d7aedfb29da0ec808fce4a5292e10a1d71debcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5a4a1dbd88213b3f4f337ea4fcd7da5e22a45365a8d33d21e170bae996a5d3d1cbd60db7417fafb06f9ac2867cfd02694a6a7be887934699378dad63872c8a2db1900d30f32b3c57e62e3fe58517312b52c60d167ba9715b198c2f78bb35e90db3c7ab0fec7e6cc57f467e9e2f7ff6b55146d05af6881db69b57d1400cedda3edbc1b28bc170bd5c1072a038cfe48ccb17b3854efe0fbefb2c0a9f2df2c00c660ee64b70fde36fcb4c2f89e3863dde834db2d4aeff3788c4f8c10c13a591fa37834aa5c0ad44ef51c06321d3905a1453b56f58d21fe808dd5e16df8e2c4be887d19b39cd2d7fc5be0c6f45e599225cb9d31e58bb2691ba6363c6f4828a9def757613150b399306325f6bda2583bfb175af886b0819146153800bb27139226ff941a5f95c53acc69d42e83b325a8c0a249eedd49f911fa231495411e881e573e0cf60eea212d50a598b4bc2bf133a3fdd185c4c813892d1f824b367166c59b1e24eea34e9d45ce173a7056640f79afab2a5d765f739598569c6d78fc778179c471f9d58d8e46c173e78891dbc78dadfdfb0b9fe6005cfe6e19f1ad4c6a74104f086d912f3b2c8b3ea812fecc8930650371271725c24ed4cc497ee37f720481a05f7a8c88e8ff81bfddb94c0a5c304844aa9962b5b8b275bf867f873772c321f289a8f1a9535e714a5043fe1099664df898afce9b42ba865e25d846548a8d81213ae824beb440732b67cd1559a053f96651f9e7718626e9df3b66a0c6ef3811f7e2b202c4e205feb956ed93a9f28fdef240ffea71f1a53728c7af1de0f0ddfae87f30a633d9e5675f845b1863cdd9d194a230d663847e39939b686682885c368a02df32b1d3ebe6d59363090c91d6ae3a164a3295a35c0d5e88cf5a559e0403128310bffb9aedd0e21574e4547cd0a25e1059da4cfb7c5f357d68a0153280b353f593a0d7d9e28b05851c0d768b10422adaf814608f4bb6bee2325220de4ad993c66dc7998bbc66645855fcd98d262a4a56f2dc285548a957fa2a22d6f50db780bb04f0a1c627f7d71d0f9cf925d57a489075585994a29d8aeabff9f6890e7b1c283aeb1594c41e22430dde57845f30ef686e39e282773d4d5bee41587d3a406220e44c592c47ef2c8bca6257e7cc3ea4c0207a809ff1f9204bb9b1b287a3afa4af58754f075dce4d64e349769e1c99a5177e7dcf59a57674ae34996689fb2a8f5459fb8a5e78ed231a757c81be050378bba3d16a958fa5d7b648525b087b27d84c0913b06f4f456f6fc058418bc7445839f537044527c5e5ad50cd82a4be46a43bfd2aeb7b29500849592ea8094cc82b85667f80ed42ba513060181500575b95c7fdd0d10cf3e9b58a7d8a61b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd6dc91eaf260381f55296af2a4de03e3a87b55bd8a046be99bddb167dff3e7406cccdb45bb2b2b412b88a021dc3e5c02787e08d09965f8032db532cab11776c757c0ea2a64cdfbbfc4bc4f98b9e27fd2c5ee59a99ad7f3b9d559e247a4f7cdb1c5109be12a7e614b21f092132bcfccd153d20bd6a6c95c7656847bebf0bb4c695be7f5fc3061cb372807c5cdf0e6bd5d84b6a1ca0171e99839ae2b4d47e3e16eefb3b74f17f1225863d674c4ab132b9d592bfe3e5638addbe0adcc247e84c61a95f35d18dd8bc4beaa61091639d4733d569f64331bd7273daf61645287c51e850e587ed92c7b8852fc6eed5771b8aefe6ecffc28186f6523ac41f1be3e196dce957111d0590ebb18aa8907e310ff48e3e98145a3ca36e06b20cd9b8c84cea286b35699ce01d39d06b8e986d518a3ddc545f671f202ed15ed37740426bc5d5b80d54bd17c4224063e399132023b4bb684ce0b2a42b176b15b4ab5bbdfc8ff57e561107827fa83b49a340319de8c268c429a34bfe059ae74e72ddac37dfeed326e96bf752c0e989d569b9bc1bcf5eb77a7867eb6306aa537cd3985e910739d0ecfbf41aafb92d854281f39e65fa7275d072f07bb755f902eaf81f1ee81e9597360fc0c17ba0b2527d008a2ba9bff21861a9448784f2ef835a4c4b922e3213397fadce60ab21a0b910408634f486147cf93791a4c7023e78c96bee1ece4098d06b4d9094ac8552fde3b58d339b1796cfbd78872aaca5064315ce5803273f492ab6103616fd4a12cf5c0ab4b5f3eaa67558ddbe05277aedf3ba8625b269abb99fec898a4a50ec4c63d9768f3c530578b01949dbafec4e5ea257c66c8979e47c920650458d05ba9dea59d02fae7168f6911cc18ef67149a6cdae039a0c509c9eea407372e0011fb3135ebe8dbfc5a9e0e7954a1d4004403897e2a47f7a8c9ebca7129427190ef459de959151e3e8d653a73bd83110289d065c041491433fa073940625548d8abfa98b39c76dc53b35dee350f811c6af051b72ee4c59558585435f3be4e2154339d3759ef470f40af57e73e4e66c307de3b7276715194d05e3c35d6f5f730d7dc202a8f87b08d75e7e3ee56ca3dbf424faca891f18f5f0886f4212961c0796ccefeece7f0472129f6bda49a3f02bc643ecad273ac91734a25b5caf40001cf430ef63ba2461ed792a7ecf154d4b80607b545a29367119795dd06811d9f9f2b5a06f8487eee71b5d3f9cffcde10d90601992fdc756af96e201c76cf4fbd659a8750d44c8f3bbb6d41fbca3cac70b7de3353f982f5924b30c1d8ef4fefbcaf09ab3ee77199533761b16944f9097c16f046a02f3564243d6fe427d34501269dd8f9f24a6d43b992a527f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8efe55112e1f3f77db386b89d4c553e23d77340f1e12abe629e39c90a8fed536da355a4f9277d2383dc8905898347db02fc9d4fbb7f96089a6b1f671123e69a340dde50756bd1982d445e824e10a7818432081e818eefd217a7dcaf2781986eddfddafd7d59d502c0538f38e97828269ec5b538a3c37765fac5be6d6925c1b080d85ab3dda83a823af1a236a31ff820dfa5b514ab00c8a2516bd9e8ad0f8474de14bfc5cfe3f8cfd19a5b1aeb08451e9d54b962ee7a84ea63fa6da0a3f3432a4a8ce1463d919678471bf103744ef9f68fed0123ee1aabee2cfc1e36ff90b51269fc39412212f75f8217b4f296644258e158f3e36095b84a319b4e5b5a090ccb4853ef15197b91e4b38f61c83faed2dde1a97091a0e0686516c0d69a339ca7fd646c6b8ee64ba41a0688fadffbefa53c91d244c084b1a8192112647172d2cff71d77e745b416c80b60e0fafb109ebae5c42b01e7f04433e09735f4f9a7436c1f3a512498c0ec3aef34edbebe1afd53ad6236116b3bef380fb31e02d0cecd03c3bb8569f16f65ae9d9517cbcb898d304a021fa7664dfe79d32e6409d93693e921c6ee85769ef081e5bbb4420298bec2893f7002beb7f1927517041823a39e2150ea2d357e2fb3b195c96c6c9939899c23e9adf1c55e0fc19a14f93dc124dd35fae1178b522f9f0f280c8428654a854cbe46e2d02f6914fcf8f218fa30908beca9849e896ab7096b6eccf847d752931a07b63e6b324b7bcf71b4103abe42af99d9f17d659eb389c511f0039c80b38622412cd085adf752a7d66e6546dfbaa5de5ba8ccb7024f21111577177621cc42f557fd7ad4099b066f7e3e3356b7614a9a577b3da76db6d39cf1ea627a1ca485630ba814dadcfd6075a4d7c99b1c0417b2bbed9a59ad85c57efc4caea60b1ea7c42c7f064ec0606f3ec14d2269920d25f509425d0afbbb7069622a2de623a809680b9bc03ead315616eff7e2c927f02f87f9cc9bf8551eca4f242b708f382ad59677bdc4510212b4afa02bb9e1ca0a085d5fd2832606165fa51de3f72fd052b2d76085bc17d32a10d5a5f15861f954d6f958900d1bb7b2b061148a60156b80dc39ce6e7ad8139184f382e5a6da3f0089b454612915e8b1cb9d7e065abb9ab4418121b359773268bcfaf4256f21b4d9928e20614d0f4c1b3d7debd7ec83e67557dd5f35b5a689f6a481007d74803134d79a1ff14474cfd7efc3b5b34763c46d1791fcbebaede3fbc51ee556a7ba67999589ca7c9077c7581445451f2add7fd72d44b1d1d61d42270dfd0315eb189abc56d9c449c75e10f57c9e85fff45f90804d312477d9a4eb5fa6ab1c612c8c0a70c1c62585f962466c8ca39cfa9cd25db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1a193df1bec31580c44b2d39566eb1e52fb8e75ea4d07625d3a812ede15cefa93ba44a94a5f29a44c6e02a4d8c3fc7e91db7fe7805d317cf09e1472f051a4a01f19753df04d87bd2b0f66aa878cf9e88d6650e2360261d7a925facb684150dd8c82540148c8d4d56a16ed5e6b4f88bb5217b9909d0e62cc35c7adea1aee7eb9fd1325c1f9d6f3cb0393d7705ce40c368938e6d74d87e08ba965b18f4e5502e63995cd4a550d53d6a366b864aab85794aa7df1c7e382ebe0c611572a9591855f3ea28fa54fdf11947032795c2a1ba89b02181f81e7e0de666743466c2f601253edbe105ad59ac3af504efaf54038b9863148f51f467ddc87266bc5ff191b02218d991cd06aec5f9c2d1a5e5e1e109dc32ee34807d1894ffd26ceee6eb150059903b871673b838a121c6190779d0cdc9f8fee80392040684c8f7f7cb64716a52568c0cb4dae984781432bb4e3ecfd243a83dd00b838a9dbb0d73f6d9d1a427a9067b2a24c92456da9ee7bdedf261e6d1236b72766c4fec818f223190a5a9c7fb17adee8f38c0bd0d12894264f16d8b4151f60f04d03be4a88b5723be3d190129d02b1389ef3ec99d993cdadb5d5ec3a3f1866cf969c276c0215f4a98403c4c5a3f5466ccc9fa24fecb9765ce89335a4485babd723137205d46a5f6dd7d554ffc31a9b2e4e4bfee51c13c2a9415f75a59bb5fc0fa1dac4406c07d8ab668027cb88e771b173890d7ed39292c98408a8d17f1b2b0915b18a94a7aaabcfd18e6d7440364495137e78bd3232264224b09067fd0b4748affb660d415a05c0f94a967ce89807522af1c4f2b13595118c17f231d256d8cbfeab95cfc8d62bbea08723d65e435e2b0ec36ae0e6efad4bfeffc0febd299c462fac2988c767627e6518970c3c73baabcf3deeee78b67531da34990af7216133b8e0222d722013dddf1885bf58973fc26fd44d2e5092e716373675ee869239d996e18dff36c1c688fa4ea108a7c355fee8d0a0f00217fc83d4ac15249c8e204b3c28d239719b0fe1d11f4c1848e9adeccd9398151a674ffe8a32bab43c11da3666285b59417b302a6cbea435976e5454579995c12506b4cb63977c6a752e0d1a32d88bdd3c301f5c97204f7a6b1cf0c6e2418528517ad46529dc7e59494ec01796d631f4d57fc1fedb271ae34d1340f16c7bf7bc21ad72e81395e7ac29a0c9a88c426217f74ab609f680bc00306f30e40d5ddde4358e6d162f96cb113d8d8318af9f1edbf308b13da7673a157a48a8f18aa21bba85fb2f2d69649bc9f961398fb564514feb197fff9ce1882101cf9594309c18ab038f1cc3d3a0b1a014dae9303a67873d6761808b90f6708e6c92c97c0bd0a8388b01029613;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9395dbe54c1ed3c219413e875cad51c3edadaa408bf4a4e15c150d573b8b08e1960099fd293d19c60117aa65ddc881280549fb13f8e1140cf73f6425856d3ffa1c392c46d5c059c7f26ded5e9151ba6349044278b751bc76ac5dd22098cb41d7cd305c263c504a5b3a5d5e8c7e968cd3c13fb25a704af5c95968c766b469da7051aa8849f9948e8fb2741f51a11c2309369d878f59cce064510695b2b7c21b3410a4aaff9f60822998bd2a9b1d80fab38d646b5c785db95ea5b1e60a238d8ee2d20ce1ce65c71e0c64ecf88c2821356cdc06c1df408db8d2e46380b44aa5ef493b9c94f3f0eb50eaba935491ba9fd34fd243e011bd141a6ffb58849046f5cff8d0c7c185f6781922c2591b7ef418c8e78867c36f04dd43cde8766cb3d87708f26d8cbf79a427695db3b7f927cc38585ee38969260a74c37b94868377d97ecec6ed55f8dd3c16a8cdfe4b8e6150c7f202457e7e6cc18300b65f513dc4a100bb2a618b06f2151a87e9a6a7e812f87ad2f00cd4e5ecf2d3c8ef4053abceaffc6170c531b3a25e31549a33dfa3034c64d81a3b36783e2ddb667fbff594366097b7ef00022a00e7e6eceb6c0100057563a149bbfcbee8809e2f364efc1102bf4e2508b8151058a3b5ebcca7eecf3c8954383f78d4024b2b5a845b5b29016e87ae14ae2662d1da4406474a3ea38c1be0374f0f6c659b3c4af172d47970904868f892dde50c07c5fac7cbd25119b425ce22edcc3b76cdaa0198bd617e3d10a951588227cedad4d2fd661701d45e1b21973b15ca173991f3631024d186cb7c36efb68014ea6856164d2e048cbf0d126f1d62c0ec7b4b28011a79daa9bca8be5a94c432f7d82f21fd56e080a07b31771461f5326265900a55b21e48c1b4332140affb3aaf32892680948d76d9925006a0fb304bee55e1a19a3adb562721031dc1553ea36cd7fbabe9c510125e6f4853ba6f9f7f34a5bbfce469bd9f38bdf395df4944a03d4cb110dd9819cbbe72d3c3c773f1ee320bff3877eddc92ec710ecca947ca706c9e19cf9c9c1218d8d93ad27b1cbd5bfb22efe6a3528ea12f6c6f256ef1fe656c2c55510628dac4a839013f393f16aed3e24dbefaec3ef2c32d03d632b0b1d8c119e0cc4e9a81cd84f717298ac8ec647e93f448b61a2bc108c73eff1d19f7a8fdf5fceaf3aa3ad999ee30d31b17e3ce8c42a51d79117c24f126e1ba3c29bb6d4468f7a5b9a5914cb0b88be42f681dab6a997dc33e0dcdefd85b597d5b46eca6592b264f9a0b9a7cde4c77d2a61448d0762bf973b36f6c5b5ab8929393654c2c9d47882f41491a75d80cb5f212e2c082abc76165cd5b683ed3a0bfdd08adee17e4dfb762fde24b2fe7340d4bfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h9d99ae1776dba9c61084b7e9f5e9467e36cf6d11e2462c8a23d7a016caab5e93846a5c3f8c0be2701429c12a6d6987f6aa260b2c082a3b4eba5a40ae78ac8fe28e2874ce7d07b06ba3cba580fcadcbed5ebead60a1e99ed7770ac662f22712871d0e5501d88564b0cddd992102558c11fb7f9dd8feafa5f151e688a6f5da99f830ae09cfe63feabee1f1383a567a06e14ef3a0da5d38260215b397ac697030d9bbcb6452f6fb4c69ff3557f8f4e550e5b8615c51b79ace10cc50e1fad54460c6c222a16a2a89bc18601299c2c4fbe8437e1e84a84eb8819b73cc30ea038e9729f82b02eba55e06e61e7d8e31760933f87e3124ff1360bfc30ae897a991ce8af4bf7e7606bc48045ba5aa61f8006442aced42ab9b8a1e175398c0b51fbd428c30ee50df3f79e049718b4cdbe596d6af1e7756c5d33bf43c451e6cfacfcc732d2f506c1217431458e58446bdd3bcf8b2d5d9bf57ad038158cc600f20be6bbff57e515bcc52cd99ad23467caac8e592e3506bacbcb848f038be7653c2a48234e9bd1b8813449adcf6c0169ee96ccef277fd689d9422b29d6629a2f84e553a9e4d36c3ec03ba6df30d684a4dbcfd24b93fe5abf70d64fa415c522eda79b521219bf3933bedeba086776a4b31936253e2e83c10094e7e1abda4f68eb56ab407b82a7344054a6cff51fc5cdd90120314d13f5b34cb8530750428ebed7c55508af9ae772dea4d64fecda1baef73fb164eabe8e52547a71db882b4c7edf81a09cefe0b36563624b561de73ffac781e52501b9671e19273e7ffd8e6987942a02ee2a3ed3f0b4e333e608440ab825381cb136bc99b12542ea82f4a95bb6a2b018753948b94c6cd009634da53fefe173e5d82a041002a101314774e3de15d2792ad8846193dcd91a99a4a371042819b21ee449c3b1ce8b0b19d670357c97524aa5afadb347c8ec200b2da3ff9d654e822aedf38542d1b3642685e23f6e22621269d912a468aab8047526a9209d0e8a144940f3dd21c03b33068bd05e32745596277564ab264f8b780e0b7dc9281e8bae9537dea55af6313cb2e3af6cec9a7b2b368ab41bf6ef1beb5885b0eb4d59d9691d9b9059cd2b54ae19c01b40f3545e0507fa0937a2e197050c86a3fa2792e11f442a644eaacb73bd558e4a6685ab657353001f8e5f7ee45a7da6167a989f1ceee1e1acae41dc2f29e96d6c4f608163703195e865ff0a0448a5e2400e6312158263738e3504b18e5b31c6775cd5136fe2a763ea7202805646edbb7b14ac4289c6cfdc018e67851994a905f5ab67279c4c8a7828e89bfabff503fb67cb6f4e251a627ccee5d377e03ce24a88e02d5cf65553a133d849b42026ec1a4cb6b07b84bc841;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h43b36ec65590828cc56149b75f578784ee61b32f09e9d607718495e8628b04a641fdf4f90365d0baf69a57bed3e9cf4971cb84d0823dfe5002fb316ba7b8f5782f75f6b666ec12d5c5377cfe27837740e1f36faa9706907ca5f863ddc8c1ba3fc26caad78fe69b2e9321a05b9c1e3bba13c465ce15113ba8867fefe9c38482af77fd89a9097270011e0c053be83471479f395516b1b75945cbc12410300a49bfe20c5f27e165a25024f95cdc871b227805243eed9305f2ea5a9c8a4ecacea7d37321935abf6c81257c9f13331d0d8bf7b6e8e93cf11140d3f860d6784b78288cbbc6cfe673454ac480b06214aa60a4537f46a176c543b848d2f49a5fabea8d0ba37872267c3717dafa14754a1b16bc82f47a33a3eb7ab822f01988056e3ffcda9a60ad8734d3f50b0070346c01a65f2e4c505d81d2ab180928643e6e96b35ff3b1ab03258f8314bceeab82059553c88e1c22a1d7533a3b812c419382134cb88c2ff6307130d1262a733b71bf1ef65635cc65b765d06c88d4b1d4ab8a78a743fb4a1efda4d362b745834be554042ce837fd905f3a0a74c270af4122fada3b4f61b82ac8c5eb99cd42f791d86ecd14400d6a38f96b15d0d4ef7c6e48786983b434ce844bc41140580b872c6dbf4d40dd7ae0c15714422797a247cd2da52d29ab1f8406f9e61ade678ae529844ac1292848ec10d0eb7fc7ae17f5b16eefbc16979cf9ac421daaef7096c4c4d166d719b425b102b3905e75fed3bbce044da484c6aa0c5f20be931b8c377ea4c01216245efc3e6a210b640d18fa7063afbc87d06cab186371c048bf87613759c322dc5b0ecf5618ec9dd9d8538645cb6cbbefdc118898a02e3cfa9aa724194c221ff9e82e420f12828c9a8a1446e718585df4110ec6a82ea047668b9eb7586a756d2cd2c5f0afc8b4b26bfa2dda5ecbf51273767379e747c00bf3fa711c84d57ab1f386da9eeb312760b856d70d82adc81e241e329fbb04b48398c74d562146b727169953b63b4ad0e1d738e7993412974b4cc18c161fe7452f12ebe63402e8bd3414407d847732726d2d7189a633d46f53e16b476289b1b6801c4085f7cfa24b200acb5855d739fc734a50b790240057963b7379dbe6b4e216e07ef495235a9f8558c3b91a8ecc762790aeb5bab86f57b2fc12380a7ec357862ba6f22da3c3d3e181067d853a9bc32bd7101d926f12c1fc5a9d2834538d122e1a58f0beac349edc3c753f15d7328502c5b3b3a57545c4ec8955db33f48425c0230c7d4c1dc668a0c25694ac96cb0de84a2cae4f23cbbe4df007ec13ddda59f3112d38116d1acfe50b6bacb7a4dc146003b48b9b4891f039304e01f8fd39906acde076fe34086c4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1bdf15736c96aa6d4e48b6fee8bc2d0b2468627ca5767fed727bc1ce457acb7ef158463bf6400a67bb6d6828e012779e252b3beab1545fb2d179f1ba86d205c35ff1354905cd72900eebe31bc78ef877f895e86891c9b9c1fe5abac66d4046092452f26b9ea3f317fdf325c0f6b38a936c0f6bdc1322a27c3032239df7ceb1b974aa45e883377d989e99b780d11e4ea022b2da2c85795c115367f7a3daaf00ee5e6117307bcddf230a50bc2449b6d0bd007eb71262019d50acfe9293966ddef923d66ef7e28d266d2d6a222d900510944d7a0c56ccbe476381d112fdc03216229464f3a7f1499bef00e12c120b5426bd97ebd1e631e70c71b15a586f31a108e31175c361130bb0b29478524f7f9c402c3850e40d92e586e306a39c6c8df70731d50ee251b5cd507aedb7113970665eee4cb9b2dbc21e285a4ec76fea375814ba5d8ba396369c1d06bad148a362569aa00dd6927cd4d29556ae21141b377003c437be8fc4a91ba0202cb896e2e32776532a3bacc2401a9b4cdb0dea6422f4219bfb978acfb3f2064df4e79cb0c62aa3bae7ae0f0dbbcbe7e0450b628b218783e2a02e84d745e9edd9401ef21f61ac420a100bba59db618443b6032786f32ce550cf8310e183cc9a5664f3a30ca306753795c3240987ea1a807fcc18b364ba2bee718d4a7962ca698317da4ca89b39682285a055c7b4631ab482e691a9247a187def2cfebac76c0a529a68cfe376f4483a84b34f7ecee0454d308a0284d7f82f301a32e0387d3e038b1a2db80bc4f8b5658ecf0018deb544dc09106277effcbd6baa6f677d11cf8506b3a7880c0aa15f7ce4aa06f0419199a6185a7f550c0f3d97ac67fc570a08784fb061e832a1083fe70527df7237f62384cd587c79fc5d71c41830329bcb5ddcb980c78a962556d830960404372815fe29ff5bd62aed6d576a46215adabb40e7f33d8964c6a8cc71488617c47e0b0bb7303efb825f1681d0162bc14fec7ad182345ec64dcb9307739b65146ea945edd7ed064cd0e36a52155038d4c60bf93c283ac8363ccee4a1f7116afe8fc07d5ead80cf1765377c700eb94627b9f42576e6ba188a112a0d06ac954ef78d8ccda2eacedb4b2fa0c1d5556a5245613533733723bc49e341f2f44957dc2f084c693e44e5c008adac825fe6cf5bb8fd661fb7fae8788efc8569a40b4153230dfa831865b36d82d0d5c62e4eb51da7133de8a25ea1b74b665476ca92e4c8937bea03d9d676e6ec380ea29dbe0728c0ea147c5e170f3b01fb4c4098b9b1f8ad6753ed7ce17ae82c49868b63df6229728f63435ceb66671b1d341f5993cc1b8a62b397dabe6481770e75c5b82732d51f765eb1527568ceb7b2bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h21164ffbf009ec563a8da0b3471566655618e184e9567a0cab52717461f0e6c46d2661cb0b7cbb3c66c30a68cc2adcdad54d1a01c62573ccfb14a7546f9569e7da9125526a1fdd406009850bae70589f3fdbc9870a417952c01d938cac83827df795dbed107bff1c1f2f43bff19536edd16ff8ea0fe52ef900bff413a69c35137f55b039a70356517b4de608443de825103f562d393e3fd46054bd2a4b8cbbe080f904ab0d2570de0e94ce205bbf0e68ebe322cf0ed3e5fb9844090760c84b44e4cd336aa4b4e504158388f289215860fc8689c508067a589e95a71735e4b650828ce57af93f18d841335c662b23b81c932052abf76af600059f427cfb918d83e5151864494d80057bef93b9c6332792c6869a21f9396e8c3365741d6654df881bf262d52ed274912611e35b82314027e57c42d556a2937ba7b7fd076afadad2b816644ea69a7cbcaf8839cf736e6522c13122ca3a8f581429bc7911cf1e0f9d292e8b3409f11417483a1400d5e27c8489f91ed55712349c37137a7bac7854939eafd24eecd5b9c303d34fb1ce843727c9c78b7b97780af547f87ceeefd3056042b54080da9eff57ff8af6c77f2a16a9685cc03ed8e2ea99d946f7e00e05099d060d670be8b36959d6611840d7d4fd3abe0b152e44af7943b1d4d12a50424dce3e9cc97ffd08545b035e8419d3497f64a89c1049529f0d8eb3fbd5dc287d913e7fb767bdb569b9487a9943e22b95524d5b4348f1b636b62bb9c315402217ac5369103ebd12f0b0175fe25bd44bcb4a7a1cece09b6b514296b7ff53f929ffdb21cca9551d336798cce75a826e52cf65dcfab4fedb09229a0d81d1cb2beb56103f2b2e040077afa46739989e49b68e509d58567f3ad82d991e9f395710c250a4d71bf4fff6faf2dc6e06d85436868c65ddffbb03c7c4a7e8689be2759754265f5f6226488db772e591009188261cea67ef54685e2c18c3b98f437a0b9cc78cb89552ed8045b508c32dd32f8ae373d92e8b008591a50b3de7fca67c315995027f2f37d2ee0037d04ee60013cf844dcf3568f1806181a5aa309bb3e35ff8fdfc1240ceee189b482f77e13946e2442704144dbeeca8ba223ca2602201b462709185f2ae9c994b51463e93e4e8767138a30313aa92995e5ca4c4d1513a670ab5b58f15d4719a0b1b07bf70da741b7014a94f9645e00334e1342c2894f13eef6b283564b9641838379e11c1111ff3a4c5d0a6025b9d5c7f1bee75e7f0645ed9dc2533d583c57c066229bf9c5569443b2091add6e011e48dde1184e5a58ea897630dbc3b3bc55da0e378bfc27150523e7a1ee22336e17bb7ae75a362b21ecc641dc6e08f57474fd925dcde1e39c292d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf92f9b78205ee0798248c06ad272a8ce0e44e30862cf77a64950cf6dff63b963e4a32d22df50f81a8b087dc74105a031fee3259eb051ade429e6df619d99ff40f86c4c8f6cecdf15f992ff0d19fcae2af666a3265d1894e3183c8d80d1e33132bf6fe0d008dc0d2dafdfc0d3da02ee40b744acc56bcb2e30e66fc7074fa047ab44f297389e922b70b8802254f401b4f345d98afba172f6369f6c5fef097b930a2f6a2b6ab518e23278565a3f891661a74c5ddf8ceedca6d952463682048d9b6338f81a20fabd944f35e663af38df5cc0ae6e21037f043499106ea16fda8b490a70860f74be055f6d97ae5be419c28528934ee6138fc728278e038e402f426c713cf85764f0d8fad08d6035300e468051a19fad75d6cec7098301ad6573728979175b06f9c11735845e97597d2bad95087a29a8a686dc4c9ab1032f42cfa7ce487e0028569d31fd440b017fa79ac37772d72d6a78fb5d086a050930199893092aa124bc317d8f6e259ff6a2e7b26b92d28938e7c00005c5140876dbdd99546e5cf35a7a380eab0962cc9c438a38439d920cbc01545dc08d86c0339cb3fb24b349333adff5227052abe569c5d0a3d3775745614f82859f2e22d75d9ac167027cba27823b14f06e24189dd0606ba816dc1d2969548a528fcd688523e1956f3755e82b68d283470b2f1272a0159c299b97a841bd52ed7c56ee5c76d4490278cbd24859843e4c4f18ea9c7f6ffbc1e2657653f41a58c580ed7b0197e221e71cb563446ac4022929e0587b1e95b944ce44d29a84c08c64554b1b29798ed7230ae7e61ed7e66c8232480abfdc0cf6ea4c9558bf5f3b439390b8d78d8126e12e56fe8e300b4e85981fe984226231b1b42474bcd577a495d18a34579ffe944397f1b55c6a1cd3344f03afdaf91d1767b115a8e898b82a9d35d499fde26e0ff6d8bf754ab6e6aaa577499e6416edbaee655a49979043131e3e92450b685c9ad865e74c2a450ad1bb9b1b618eee48cc879033280e6c6e8f5f058a65e33d6bec1e7b7a29a4b7712e4c644dfe91e7853b1158c12919d5690e484c5b9d6875719bc037aa24821b3c169c22765c407e875e79d0cb5573bc227e5b65c305a54601974362bc87dfcecda65aca9bad6974383322c34c455d9227a5934c58d6119d85e3db8a10fc491c12c90af2a61ca8300dcc808a3400184810396edde66efa3973d69410942ff2c23a527ded3779e3a7f6b4c33b72d8c714d34aeabf8db076b5a76df6f76aa5ec23b898efc3869e14378746251adb1d47d2ceff1e30cb414bb9c2f2e03dbf163fbe7bd34a905cd5d5689f1515c12dd75ebd4cb2eae68716da6bd3ab91f544b69084dfcf047bd747ed83a508459c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf5b478c0cc42f0b30b804c76e996b2870ac96111dc40f0bd182dd0245c9c2b37b9dfadf75a23fdcd6bb2854002990f708e0ec389f6fc341cae37fb89e218069a85ea995df22ed17bf2505a9bc654304f5d884e26cbad2ea99aa1e99e777eeda8d9bd3046d04331ffbe64610efa488d43fad16363ea1f9b6946db10687ca559b78cded24eb1ad488eb5682e13adceff262a030b0d14e852291575bd9f8b57f3876de6d7dfa3455deecb1ce02a02215a15aaa5529c0446b707a7e87783778406c4b7ff3bf02218d1deebff307a74a468cabb1113da8621330fb34f27a8ffbcdf0704ba5a1dfd6353b8a0b8504ba51110ea6703ce3cc441f1eaa1cad5b4f25ab551a3e4716220727a66c7bb8e9c33e20c4215cdee945c754c5d3f754e0caf65dbee6f613b6080294e4d44d7fda7c5a2bb126590ad4e0be4e60e2c2e27d953f479e87848abb9279adbd510c9affaf3a4d2401d4c6d8a376afacc64237d4815930506762065928cba7c7c78435a78d061d7caab4d2bc6df7a97b72f279f461e73e7e2335dd2880e1b07486206b098a5136b23ae89054b7d707ad57d4a7f462b9cb6e1deb6e38e664a4a9e848cc0b5eec19680d08998b6d80e38e2321d85d8d1a572f103b04a987fed6e3e735eb93b81233e47bd26a2472177ce3f88cd2a20a8e5111744fb5f3229b8fc9abcd0ebe0b5ae0b167bb74ea6f48f4ed15cb04aa21de39ecb64836536fed2591f82a422d76ae1d09669356fd16f261e428bb34af5f48e7a47897448990f43914e549d8bfdf67c0c52f31b80cc6de2fa47d4df9e61b27431958c303a864e77c2a7e76cd31c2f164d3fa125e665dd2765ec037bbf139f4f4bb34c2f68ef530e54816e01d5dedd4bfb9b069490120bbec65aae1fb00168e26513e3e3a05950ea66838267e81ae2efc2ccb5f5d83aa9e85ef1581c7642f5a4907ebce017b3e40c128fca1d3664536eb5d261a732f5216d7fb00496f927b63b5e11871d6f07a47c6bd32868f4e04cb9592ea680e5b647e1bb5eb68d29c30c0e26c5a50094ebbbec80c908171a3c894336152b26eed8864ce69cd39fb8fa17bdee0dd369991f8bedef744e29f63d6eaf26a870a44db09772731b02b049b3932486c267e75e56066cacf4cff861e948e4c96a81aba99862b100543a8c95d4d201fa7ea5c897d39922412b814a0e42c2cd3a519523a4315c987ea176d633fb693680407d36c5bbd9aeb89401091441daf4f09643bf57375c969236891175c0b143a3cd4ac16d4f5a5697d3a0f83088e06f07c851d250df676c9812e45d60c395119fe156e240fb62325acfa87360e785d61e6df6cc3e4f80dd3272762bbeb6aab0463af58b6dd5ac4cde69e009c1e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4d49f5c671db687bab93ab02be73a3f80aaf902f2b012b135b016d6d1ca1e1c3a7b23b6026a75fb99c013f154383ed2c599e73aa43b938e8f46b9d75f59819aed6716cd3101bffdc9d6d00832845b47644e2ae50f8458dd813ba95d246756a58167ddf93fa696cfe5f057a083241c6a32039b4657a4efe3d318dfa6aebcff8ad6f464e7ba7799d7a00b11e9f63741c856554ae870fb8a07ed07b47850a60761bca8e9bb5054edc24bae94d9c5de66c15ce5313e7eb92806f54d02be6cd650b7b50610077939b7df23337a297220d1b48df1c4823bfedeb1d21595a5ef618dba981cf05db68a0d03cf75648009e6de04a9b33fc1f07703ba88fab93f09670cd57de16d0a334f6584c02ae8098f664e6152e69df0220c9dd84ed51abfba8167e5de388c5780ee402c3d985fe5a6eca61e20b353a3a24e0d74fee51d808d14b100e85f99a032686d82cff2848bc932f6a837f7356f4ba011a65b2b88f4325aeed2bbbf1685f068f277cedd36ecf40d8bcf7f5835b25a8423edb67da1d1c076d2cac9918b2d80f9f2288322ecaae40b8b42b88560261949feced2d41119d25bdda02c053da6881d85600c78e113b0d5a8504aeddaa98a4b6e953c4d4968f8ec0e34e184f9be96809c7e826d346ed33334043913d66944ac2fb7053479f331bc72582476810a83f56a8fe32b907b21775146fc881391491023fdfe81ad4ad399600bf7fce5db662259647d450e96605d4f8ba3d69c3880745566a36bc74968ff90c75473c181dc1962cfcda2614b709d26906a818d636ca4d37c333193b7bc39b7e630740204673d504e4e5791c49ff8be1629443962966675c46be9526a69f72a99a74ddd3d3d08d4a2b0c85f690f858ca52f2416ab9971820664e56fd01e06cfcca5a3c30b0fc58f333ef58020451bdc755054492330998939f2b8ee0c86a4d2a9af764e36b460259f94719a6ab61977b0c2d6aff2f5e742c92858d31bd83dd23c9436fb78e9f9b15da17fc36f3509f60fd6ffe56e47116e8955ea6e07496f4a3d1a4af5247b0b941afc4e9d935356733eb6cccf8bf7d978291b35efd438d8aaf1754c61c8bc22c2995d5663c5a8e1dc623b0601bd857f2574795e463da38b667f0a629819640df2ed1aeaef27d8dd69c23c15b4a79187893459d81dff032d14571793c072e7a469da0bac6d6980f3845a46f424208f82ce5318a53ee3bc1d1da4ab03dc2f46c611862fa6cbdd8c3993ea360ef614c9483ccbce00da70cc141d8c239cf3b082cd26864b86e1972210ac91a230e1eff71127448b955bb95dd7ba4f7af78e1d1ca876dd5b10761ffe34f02e4d0e702d8541376074121af5ad97c686582896b2a59c108a78d44b3a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h83e6f858002934a767889538875ae34fdbbe42fdeeb2d16134918aac9caca9c1b9feb7a5f47cd29704973592113519f250d7e721978fb944c4293a9ab646dac1e778b007d22b5281ad133a837043f5ef6f71ddf775d70a96cf395bdc6909992605e657692318554196a03f8936894365d98e23a3055cc96a7c58bfd81b7b15664d7bcdc482e55b4c97d4f21f3c72385db6348fc09927e1362c12c4595940eafafb2f8b369b057d807c85085cf6b126a2d67c1bb3d5bf4c458ac241716e7a184e0f1fae096419f83ccf226e7b764edd3ab0b98ce39648c566dfbd837e3567f3de20d7a5de5821658f412aeb9a587723442ecbde8a1866ee1d72731f4819c4eceaa50fe77ce66407e8e139eb61ba3a39bd614e66ae5482046b8cb317bd0581b4959ff0c7955b82d00a1fa7da5faaf61a4489fe1214fc75361eae4187907452f69a8734d663783fdac9a6c63fb9e63ed7675e1db5d9d5cd222404bedcc43989a8e5ff1ae4452d8c6fe1bbf5ae5d0aaadcb2bd86032d2d0e29ea8a15a215332cce07c43e128ac2b03e3afb502246b3110c501df06c07795a324b352492753ee403ac1d31845070d5c84065434b8755e25b2ea8c34ad63a946cfdf3601f694f144061f570a08b1638b73eb6049d1b05a781dbe1e49df4c1f58136185741482624f7e5aebbc9f4d5c9821462f1146eecf8f315e1e463d5fd813e2ec2d4901b0202a7ff429c70ce1de7dbb4bbb295112faeb989f900e1969e22c3b2b156c8ede015b78f793716a544043822e6190b7461ac319b3bb869de83a5f0dbaca5ebc04e4901b4737903869b71e94ad297dcecf29c678b2160e72045be5a3bcdf9f077f7efa7ad14fa9bfcbdd59b22f156c61c051166cd4faa2e5c44afac16b9066d8b58e96068ac55e74ac949b8ea96af84c9378f8b98323faa7836f862a4a19a2c8a495a0bfa4c76aa3f9485b71cac0a8dd4ba273ac937c6a382f160f24819a5a3ce8460440e6337e4f2415f64b77423ac2592de6bb05b8b95cb0894780746b25214800cdc884d35cdfa0d44187900f33ae06b2eefadd11968ec41642ed72631517346ab0f17f97e7f6981ecfb8a286644a43c3f769f6493a9ab8a42a2f23dc360b4622ed12c1000ac423c3f7767571bc80ff50b4cd6e3018d1c9e2e3b75e55a514347b3a3450e871e070b98e729936d90f58b2db8450008b222b991a7c30f0a87fa1fd09d81f1d314177876bd7a2e7994afac37631c86a1752ae2d6176f84b6fa0453f2278b31970301f161a4a0e2ac3c694364d12f98aa573f50490c06e59b5551faa195dfef62d811583716c6546b7a23db252042edd68e5eccdad82cc6cfe8ca1edfaabe8bd42aeec267b6726deab36b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1e4063a9529fd5926be5701a704ce5d0b6ee2df1567ca11c177c336677c44c94ee71ea830cb329e69ec7aabb2e992e434d8e74c576b7ebc16241e925c6c304ff597643b45b1cc55d4fe24d188ade18f501d07c86a396dfa36b914fb0b7a22d63cf111e4fe42a4b4631e479ea2ada83214997aac7d58a020eee47b38a8c0475441b7849ca741b024fe9a4441e973143b40c9ff665f961bf099f219925ad152bf1a035b23f51e4e483a550e0cd5fc8801ca2bd3dccb120ae8c86c472ad3396828530b790ead228dbefcb1c6afb8554f63196a8747b3a5bbc1d597b62db8638e319943aa2de8e252b6023cbcff55873b069e6296c1f287c4fd3552594b7eddfa66eeb018df7aebb822738129c8432b24874c442fb922048e9416508c7db9c7b4bc711340f683653d48f50b64a72af74511042bb1e42df5b6f4bef9127b46581f523b5533f5080d0d0ff538722e42377ea9310e5a568cf695915344c8d9699cebca5c0f8804bf3c33ae455e863713100b20203c704a4d8f4004862f0f1f019fb109e47f0aeaf28746c3d9d7cc46a5faacabdf5d1b60e8959d671b99b3d3973d78f5ed061b1021874185a0c03fd29c8cd32e0ca6c001edd250ff2b6372f89150c95ea101d4cf127176ffcc33ee20d178df73ee023c261ce505ecbf11f0e5a58132a826fd4c1553d910442a586b7f88453432665df8067008d2bf4a389081b56e2c5d5a1e4406f3819e785451306d966ad72afd0344fb68966b385834405b2af81c6ae610e0971c34e39a447e3f040c1c95287d6285b848304ef75035f1c639853b5f215da39745e1d9959aa0863fdb54afded6365249a7c79bc03127e15479817830b1386eba24c07bb6879cd9a252515f2d02ce2a626b664d068cbc1992dc374f88d9077fe03b657b16a099771f8da9353dca421f6fcd2c85f996403588de0d874a8628f14ef24347f60647de06c74b2d62533ee841a4a2c344182bbb8c01ee5d8e9ccaa41a6836bc5ac9dc149b03402a5b53c7f27fd34e32ee296207e7998fa554e971f869e8ea7ab1ebda022d9a7f398e977dc4b6caea5bc5759929305a28fd3e1b72fc3bf114f3f621477b938df7d94a7f6872d60757199dd93042c9c13d9e2bc73229cfa68eb145e9145047e4cb2d8de8ac4e64a8df2a551c91beb48136c40a2c66a8c5197553b1f16e0e713ad71ac0c92a14ed4ec090883e46c1ec2d4d67e7a9259a27e64c58b62457c2fbd021b892c8df59ffab687cc8bae0f575c97fae79229a3d6fce1f5c33cc3dda58c37debecb89779301a0179da3959ac03a57d97c8525d11aa6b5c9182a9365a3227298bef2256e56da89acd2602070dab2b7c18516c7227278d118e7957dd3ce7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h2e5e26417667cbc4f996a13854bd6d4b654843b45fd0c77a3b2f7169fe7ec8be0ccec2d70294614e3df3f49b2627da20fb9b815f92c5e046b01152d32b604209849d3c2be378f64f1d08299c6a7be850dbfc3cb8ecc448209d9c203a5d88a5f72373235949a3c5d1d49e23f8f4703827053d0e1e4754b8c8419d950655a20ae27a4a9b42c7af701369fcf8f273a5f1ab1c4da771305ace545810824a1c02c9476158ba9fe56dc70fd32dc4f79cd33638ffe12565bb7deae03705da7552250407ffc7c2788522598e47bb4b3313fd07afd55f701ca2715b0b283760d23cd9d52d24705eff01c022102d04ca0320dcebb0ef7174facf35ff29107e0b239311647358c5600bc74a3cfda132b654b6941e742fe3d41fecaa105c2cb38a589cce97b5bc613c9be382586328b021e24e8bd27b4cb6599fec0d3f863d6012ce910ceba1079f39cdbeade124a171a9a6e087dc30f227f8193fed9af10c4a5465d6f9eef34757197759eb16a4fe62c3b6800f99f4f78b5a548efca5d06070c98b069b862d3dae4b534dedf59230236c66eda303f8188d6fe85af685b901fa5bbc8012e534938cddb8a8d36fc5e2a730410434d207b6f8c4c17d6ecd446d98b655737799ab5961df8a6da19930cf9891ef2250ca7ed2aa0248cb2e44be0b9e59c87284a6b4749501681e17e139887c7c9263cf0f2ddba6c117358037cb33eebd2d1cb5e2c5afca88e142ce5ff1c7aa0b3e2f46dc8d068c1fdcae263de643e218dc413011bc3eca2fa4bdba133bd87764ec9ff7b76987d66221e69ce2e2dd28efcfce2845a387c332f832124bfb794e1751684525c8c37ab412e30b873bddb960800cfe0b06e0e1b1c016f3b87756d2940f52620b80bf39d9aae741e42983c1d38727bd03bf7135568e9c7f5defd8a263054523247ae9b0654d0f3ac55925891f3ca2f7838650a2d3c7e95ef9f45cb8bf7d71fc44a4ba7fb1af7818890bc39b9bef73f50eb075d20cabd04f2041d2762f3904e96679d60c6ed7bfabea53d361d68719af8f3b902b41bccbe56a47c7b4c0326c5076a9330d95ad3fb2f2bafbfe31b34d7aed0b7277a1a0d581ab780a4264d4b59c4b11356dc7ce896074626749bca729aa62cf3b9c3bb783c0d4826ff15ca747b526a9ec8db404929ac8bbf72c960bebb32096367d50d6181e3000f4ca9266c8f4123e891dc4809619dd79cb5f45a41ee8fec2b307486b503d3d6a624d6b481f7318ae569783a851aab7a517b415b5ca6bed31b4911b93c28838c47921d12baf06a15291464e78b1c6cf7d0d5a0b8267a82bf43818a110e981a15be2343798c33ca4f1012eba0c7d9bb3831ec6107c0f590db0264be6d954cece076ebcd2ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb4809062509de27ae5b84ce6a7e29c6478878429db9a4446dc4e49e783b905f6d86a11e963fdf4aef17821aeb813f76f392499d072be4782657918733ee06ec9dec2543937f0e68d3d60edc668a841d50bf01888dde6a9e32fcfe8978c8e13e11fa8377410a39291270b6c811850308fafa03ab868c0ce0ad7467b6e7a9a6bbb1f4b22a04c65e525ff40e53b1c7579fe080cf2a8a8174d721358df0acb52c8e3acc078eb610cb0ed47498d6f5c379860d698a3265676fb0bad162c45f24365943d4bf8eebe6cf8ceaac6781789563799ce977b2cb40687627caa886a4fe52c8832896e5d2e7a903abcbf037ff32edebffde760e9b0aa47ffb5aeda07590fbbee22e1ee9c2b281bc6cd4fdc19140c75adc6a2d3372fef2007339050fc2de22263f63cbbfa78f7025fb87762d43b37d7232d7add308a13079851134207cf382e52a26cb1018f18b72ac5cdbd1fb615278c34baf56275a09b28d19b025c2d4cf27e01d25fe6937c2840bcd3ad9712281fb535614dbc23f22daff485d4d86101bbce731eb1e3d03ca03addafe1c3a10c50a9dee8740d42a9e1addc42ff7893335ec74d5fec2fafdae8c5f3b2a395ded971b69d1f2a6e6e23a1e95c9300b4feab080ae3d1c418fa5595804b856a825ec1f983aaf49ce553b91a1615d49de9c5ceb4e0570d23a68c58aa94b4045fbf185d541443438e62d42f283352c99d841f0646c7f8933ab2db1096b8035a42dcbc5f538befd75e72b52c6778546ed6ec1d44e0a1c24def69b7d953b210172eb3101332a0bc6f0f3514afd2806c5dba0004ca2b0741c930f4e7605a10827067d2b0422fb213b5c8e4b9e8b261daecce4e92a11d9a2b430138cf71d3dd22029811731e3d4807ec563b78ac951ebec5da3e3d857235f08dcb6489ec0096b3310c94d9cc46dac25ea53f0d336cd65625ea25aaa48ac5059f2c3eca7c104127bcc57855e540645de7fe27a59222d78f235f4faab98c364eba17a90254cf4a379ff02c657fab035e6bff125681e0f57a45dc24c9d86220bbf78a1c68dd6b959a1e4c356ba6bfd8981bbb5af3373e231519df3fcef4a7f85607c615ab1c3dcc1fcda460564f9814264a55972ccbfaf9c9225150d83096f70db2b23b5fc9aa645c250daab35ea138558c9c46eb3d2408995fdf839b7fea1f058a240e25e199ecf244bd6896093cbc266a0ecd8d0782fba27afc9f782f177888c782d3d1cb3e44c96c27b44fadeb4fb899c3dbf72bbd0bb0d62cfcae530fd822303629011bf824e948dc712647d23b04abf6e8bb421877403b2850fc61322d669557ec841c72587bcd9ad09760851c110d4001d464c61c0c26cd90275c532de5ca98da1560489146d73e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he19a80cf03a5ce7b025b2b9096dc1287c99bc0297ba6ee4443a8de8e26ba18240cf5984268d49804ff7727bff8d68f70fd2d76651713552d004cd158431db19113180dc0a9b94c0f88b27b6c5a696096b7c15525ce2db819900f15954a4969061d74cd6de7f1e36bf6319378c8501d54e7dcea7876402f39006383217fd61948e5f45f7e1e643f96ec97edcab8fc74ff410ab550b926b8762a7cbcf97d8358925f2b50a0bc612077c8765096616f1b94b5b1e964117494ab3ac58d6e87a9a9eef947e4e1a99bbe23cccc38c61c73339dfbd03e8428f2bd481a30ae992341dbcbb338b44e86d74e1fe669c1552b535074f850545983c04992581492383f48ec58f8ddf7fc791eff9456e5533cb218a6c1b84699ef8ad4dc6e9aa22f40ee46bf056176275e4f83ae62adae595b6409c16d8210c262f80995586aceacf83f311bc3dedaf1d0cbd25b0a0eb75f4f5119cad6613f287c4b0737e72deae5e2f4ef38d61139b1ca7b464c2d31179d793c7dd8a2b861d7460f616aa3866cf605349cfc604062914ee1d23eaf0e4f2f807f518dd85a923d9bc327c3ae768307bf5244081d5c33762daf45640427e7f1aa4cb42acd22bd3e0f15721b0ea242625618c8c91c8e6c35821811113ae1e272f354df020868fb80428bb30f9842891e57274d97506a56c687016c6cb6951f5742ee9166800d556852874d6efcd3b7ef4f910df3031a4fa848872cc1b5ed976bf789658a756fdd0d919fd263dd32bfa0663a4cf45a6cfed66dbd6108efa589fb4c910246ef5211328fa89f61467bd518c217b193841f74dcf14c3695652b35bc22a131bf13b2e5936356165b0d11e48c27e1f0d4cf45695d529cbdd9e8a1633e97bce1ec5418ffb32c77c9e51a8d75c4d5ccc31d769548600a957cd7ffe00c22f346bc7b90684d56a2e92d8c2a2931daf06aa2536455a6d0803395fbd1e2e8555cfe784aa1e8f7a3a0e514bf2b20c2ad4edfeaecabcfb29f1c16745e6178d6c872613eac0f531f61e106a4ac2131835b9dd0f669285e2b65aa69bf42cc51bd474c962aa22266f4aa0db7691e04d7feb4a8a43f6dcc957eb6d85fa50b41a5eae52084c962a53af8683981a7f79bb09b6830f4186ee829e0059515c1c854bdeaee1a4ceac43714f7c81e21986f93ce8e85d4d4cab84fecd5551ac3eef4ff107402be4873d103a6d8853267a7ff6dde3a7f38c231e5e9da1e7d68e253c2ca7a97eca8df58f67eb3bbac24433161a55f2394315f5d44e2706c00f914e35e1a99ae914407a910f27a9a10f69f1927aadfcc60b247f50ef883e884bd08c5d0b773a2b5298e767effa622b77421249b1d76b3e8e82821888a79373dc27bd0994abc378965;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3f429a9266dc4694fd268c597cd3927bc96a46962da78caba5c4999527bd2f6c33445f6fca2e3ed3138b6236051a9834cd1a55013c7ef8e41da7e09d662d54591c303971e7b7a09b1b5c5745495957948678e1a2d18e3cdbaebfa59bacdd57b6e2614bb8a2d15e381a6ae43c0f75bffd6e6881da914bd951a7d4e0204f199df0c10c6adfd5be0f0ac64983a59f158aa17f422734499958b9bb6737d6f25bbdad4c3356a5baa328b8944b83f25c882738b34f5a0837b7a7261ee14bfbb8fba1d2823658bb8f673c34055e8e558917053f006f51320652e865c4fbd7df2c0ae93e5cfa6e274102c0bfaf0d92145931f8d2884cbcf9b79bc30eaaa07b990e8f786dc5b31daf7fbf3b95ebf6745d59cd55d3bd3b1b695aad935bb12806c88572f68ec78cfed7947be735c9682d34dcbcd62fbd30bcac42de0f8097719a3a28af1eb6bdc17a38d35f04d2034562da485b69bc18385e45d0c74760785b7e82aaa0510f6ca2dad7e908397df0d02df57c19efce2cc2564b1d0f2452579be78957d3e0748ba9ff05e1c7776585d7df516384fdeb0029da9c118e5772e53a75f01139dce2fd1344f72d71f55516c5a16a55c2f6b8fe94180e7126533538ffb92a1718e8b672469dad173a4522dd7b7842b93ad50cebcebb2f61742a90201d93555da1a94465c7a46923e72f0d81ed455cc40fb6b282322944ff6713b675d8602cb8b14605fc3c38c64756e666077f4b297da6f645a016633094e16bc6c8f6b8d5b62b3dd0e821cad684d60ecfe76eb1b1e27e2523b6b21fcd9cec7ad470a15ab287cf5f1e623abca6bb9e9dc4af6e6f4d8afe298a1a8ff86ce6e6bbb2eb5394d747144812fd3bd9481721409466baf1c6a799a85b14f61b1c9668bd15eded7df92c28605a1dd491fc5f1b1e8fdbe499d38246e39847a49a32e632202efa61ac693a1eb6f8f05835ef918a8679312c2dfe1ad35ae5f11c52b00456d6d29e28657c63dd613a22ad6b45fb62cdb33e79604cdaf0b1f6010213bcaa8a7a5bd41cb3e78d12979f2473f47cb313e0f452ba609867b0ca081abc6ce15e6dcfda838e95431d2e1e480a92daf4cfba8c1fc37d346fd63eb5b398fedbd0ccd93f8827ac118c064121fa5aa91fcdb19c5555b2b00ef86f47b0b062af1c062abf9703fb1033679c3e0fef0f58ff5d44d5b3de7fe8de99e66a7de8b0744112c4585ffc57ede9f89e7adffcc07a4af5ea64e9426d9b9a8d2050f32df623a0f7f99eb6641c6cb5c2dced25411aa2d220edefa3ec096b156da2786a6a790ea516d78126029ebeca3c8b37447dd9231d422b9f923e5e662d1b80bdff49cd95ad709ca292ab8c8c256beb4191439edc9f65fe7d1182b5be91f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha2b380428955094830576e0dd68ec2bd67550a2e5ed3df43ee7b60b09e4972cf39513c520843370cc58865c26cee4acc59030bae0a2076d9ce8cfb840bb4d90136a9cbf9e9b9596731f90aaeb118161c555afaf9f00b49dab7ad975b62cea5157831ffc494c4a72a59b5d667f1de434d71d0228e7a2fc900fbd0501669c070e120f9ce68cf1c9843a04abbd071f5252ee2998b79f76b2298b9840b8e81387f031fabc96c5bbfabf13232fda24b5559fdd534a48dbca00f3233f3f49f78ce71c827e8b0b48c5c9d932adb312e70c8044584922f377fb2fc9f8a07621aa9a59fff1fe93ff9f471205d7ce2d0910ad95fd54452e44fc5e6e04ea2ba3f6bb686d3953e576d023975e39b6e8e557f86596e01dcc6e9a7baf1f653c5e09b92c1250da1b3c82ce6f04a710d436f94c413d7bcc0c9360df09fe8a4acc6047a2c3f34ecbedebeb8d621ce2714cf1cfd2329b92224cd15952b1b25980a285464e586063eaf907b31b972018f06ef7cc0d369bb9a81d1d94f0300d5420e838338396e48153134fa1fc553e529c04b069a19513f301236312d59a194895b353806c4fcecbc5279db3841b87680b5d3e17f73fe9063d0059f5c002cbca7feb0f0ba74bebd7dad5d6a718d8c6211a09f06607c0204533c69b31482a42841a774e05a550e01f8ca3e69ed4e25257e382ae1ab7419f33379a88075fedf9a09adc48d97c28a69efd9aeaa35261aaf37edd20714f70716efc662facd2e5ca3685213ba560c8a9aa2a64cc34448d53322acc55e1d0ccb3a2a0bd4d982339dcf22f8b6073af148e4376908d29d15e66414b68d01d2f9d4af9e899b5dc2293b28303b0e778abbe77f83ab67561e8aca0440141e5561f58b4b2221f24d774ac85f1a5f1ec38ff1a318de2b3bc08cfd305dbc716b47f5ee60ebdd71d72c7dee54125b7936e6f0075b593303f912e290129b5a2870051c5aceead02a57f436eacb733ac485eac9068e6e0ec59e4da6b68ef345c9295a4d9746290fc7840fda2c1888c724f6eedaab5997d662cb42b506eb2d6b3c1b97cc3b2cb6698a2b2b7d5e7989a281cbb0bb4a102c16fd2108cbf2b4bbc3a215a6b8ee8957d786cd8c9b5fd00841c1f1fa782867305893deb543edcd67f146bd2467feda22e2fd0e1d2daaec673d860709895d512333288b51348e7e46551af2e971e5314f9b8cf89ccfc2574d5100db20d06b069e65931cd071b1cc23369a34f93f39d55351eda2e3935f450b29bf34baa9df2698b34a9eb6932e48bfdf550458bb68b26218dbc29f031ca955f679b8db859dcd4a963ebb8d122ddf7e1bc69bea212329059e71b0fe43370928b2f26abc4c93147ca562fc2370b7ad0f82a11d78fe3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8cde5a19104209d128e42c5d2c5891fcd2ebc00334ea99b3de077e55209c40a9441b7e8e3c51aeb2ca6cf5be29bdaa82d7223376c3ab8bce7c0ef00b9a4909aeb7f1bdd040b5e21aad4b7bb34b891df96946e0e6425a257a2bac11761ca9544e840aaa7531079ec2c37f0af5fe4283651f89a16720ef61d20dc77a810987d50953b59b18afe8ef864b41c74d84b4269582e8daed1c10502eecb875778585ad5b7b399b14562d76cd421b84d7fd1ee66fdee35e6a88cc94242bd6282398c33af298a98ab0f9e054ffb4d1b9f8779c6fb8fbd90a2fea9ef746ceecb5049c829abf2793632a207aeaf2bfa6a7850c5429b3a1ae1e3663477d347b7d41c80a5aa33f8f14ad0d3ae213ba6060dbcb2e33d3145eae39243caec6a082ac4b2f67f8ee91fd1143f511d4e3d44234deca81a84b126e9ab458541bb24feb5779a549af1d149caaae1d548105fe7b4539fdc90bd92751f919bd32230ed4efb43e033815855185785da2af760d8c84fad9b9d6238d70f5f787d6cda998bc8442db3c3551fb636c46a7003ffc049b5d5d8c3b68535589d2e7a3c2b9841c331b12b40310118139bc1f1c0d41ce3a5fd65c2c8a47c7907e9a727faace07879cef66ebfa50b4117c524d781e81e639e486797a8f9cfdce955989a1be1dfe63f5b79a4bbd86cf791ae9187c5f3700fc5d280a56de862831b2a1e8a66749906d7d4f17fb660a32d88d6071987fe3fce67f73130620346155f68858cfab4e0439b62a61f873e11427fb1199293c94779ae9fef503c4071491a3078f2b344f29445af7d627ccbbd47ccfd957a1edee2fd53c4c8b478282f038c44dc7512f235337d08376d8af5d07aed3eb9aa66b7d0732dd25bd0e633dfb608d8543522ab1827fb7b3d7ffc8c64a21e32cabe147aa6d756ed4db30a1417bdf9e9d17f0f9a139413510744f539529f00e81a848d156bdb04c5543a8b1479ee6166de7d7ed3be116c93544aba407055399bade118a5513f1d3dc88ecf56ca1c1d65a96cc87bc4a98e49bcfa15b6819b18f0e3f16da650d212eb9b4c7f120717b7d48187e981c930bde7b45af8b0c007ab9ae3606cf8a13bf440314ab580ddad1fd849d9e309f8be1f231c674615a317c759804fb2b097a02bcb6a95cdc5924c929f9dfc6103e3b1a64abfd749641e86fce59963696a25b23edf5674b54e5d48f2d07c83177a26ca4f7b20d534d06435622f8517eafdf9718b0b6f440551eeef1c61c0f2c873904f8bb90c4ee91c923585902d3dfbc522b373e364a9a7676161cbae92baecaf3d1579d270ba3ebb69f1057531dff6b61731a3d1adc799ba843723a9701dd2d62d5f0f667ebc3575775fc9edd6f6568ba3ad2d7a437abc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h690d50ba737a341f97b4ef068419af4dbfdcf3d715531fc4bb2037d3abbc8534436809a99db6c80dad27ab89a325627841f0eda1a0639e58ff41a54b001a7bade769ed58c1a83f2b38753fd69e417f8ddd86e47b52fb11abc747217c7643756df20116384cc21cfe4989a73e68bf921c36203f00a8b721c1712dbd11e22d1195ad57168a02ffcbf94d136fb4618a292714701fcf7de991863565b8b96bee68586a510adfbe1d0d2232f3104553f5883e554517c222653a4bdeda7f5c65938255ce32f06e58c9afacb3031d87cd4d3621dd16086e074ff0074d015792fa3b5d84ee715614f7266082c6fb84be089c5c3c32f6aef5c99dd7e204b8dd186569d96e6e898746e4eb3f80d9be982790a34c36fabfcec371cc96fca0dfb61067b08b95d29b428985e801504aa3d5c1d002ba4a04a960ea3af91951ab0a2cc75cbd33a916889b1121da69f5d0901a26a64d5283e3b98b23ae1c813bf01ba1fa8a75072162af8bb269823c50b4eaa5efd477bbe50a4143093339762d0582413f1bf0d8992434d88d141f23d7183ff1d42183ada95ea53ad4221c72c0d13497040af7214de416df2fa5016aea4d2b996a6975c76840d3e4ddf7452f3f93f57f5d0403d37f0f83bdc673ebe6028d7c3e6017396d18741ec507f067e580febffb4384788a0ec6f3669e4860712536267b758d54627182c73aaa08416eba2c2b227dec661c57d01427e2585473898989dffd2b44d236105d6164ba2641454b27baae12dfd921042c4e3de410f68b7866bc6bed65f7e43d2abc434c881c25b69615d1931377d8f34d3e4f5ec09bdd2a509c4d83e8b2d9d1eb56350d783ef37102bb9293a4435f9e4480043e9f8cb43caef0b6983c7b1ceb1ecdd4c70ccb479f62e48ee4fc9ed1770d352ef8605c1ca02558699c330cf4a249bfd87ef6f5e7a47042a92d6de742970ec7376f11d3e5cf51b280cdeb09823e5630cb13bdc67c40c0f0a75a67751280f81df2f9e6fa83e8d819d21be9654140d8819f7dd64e4c7b61ba69a63cfc9b170c82c01ae8cf29ad5a5dcc1e3a965ec6c607fc5c6c38751f9bc500ab637f0799b59c22f271fb1b26a3253a57f36204b55a61b736e5cb562ac5df4803f00d0065cb52c3c1ad87b1d514b2e189292896f54fbdb1d4b38bb99b4aecf413ab2d1afa033301d7968fe3ae578e0fe7daf956986b89c3b5f6897484d793d9558d768a719386a7fec040939d0cba8443c82e182150bf1569c8b7234869aaaf4c648e30daa6d49ddd458413dbe7d8f62ae8004384182b327f0af3904df76a92fd752b164706b19329b0043b5f3b6fad2a81803252fa09479bd10c2aceb1cd81977d65537b80675f4d645fb3f5cacbca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hfb7768e394467780a66e46dc72bf4beb22dc94353cedd756e273025726521ae996b0c04187f3c13b62a3e93bcc48507e6e8045cae78c5d02263828e8cfbe4a6297f1c84ba66377683a0ed12b8a36d14a8654aa51caa9ba13e5dfa8fced40001fd51abbe29b59d88a97801ab5a4e33fdde58be3f5ad0a401c3d29c5e998726cf8191fe4cd82852b6c527e087951548fb9bbb752b5c7f61ea06cbc12f225c5cf08eb3a83470ed522b961a19390a4e25c10912f9e9dff76e2188b0ec8554d926608fe03feb6a4de1f36ef7e228096f7bf00f84860c82de05ebb9810ad2a5f196a78b4ac8c93627421ab1b98fc8320314280ea50a556d3bf52138aba8f00c7ae7f89cf0a97fbd3e7b4b25357798d106695b22665d4c9e2cd30f7715a1a09e700615238570a69cf73f76378a814c3bd7105549584b40f16e4a61a3b3fc453ffee0a57045198422bb6e5412568bbfc58d65d30010b268201eacc1122c8d082f00e3bf1c0f5c54fad91b3e7f40b005bb8cd5cc2a99b1c1c2f5112f99740fc3352804b24583fbebbf0c37ff4a6cdfe6891e844dbc967e6655aaa6a763b0b7fcaeee6f5d45dbf9017718fbb0476070f968bbe7c0afe176c42d8ff7574bbb02685a268f8b316d45e58fd3ada65b367b1f14e5f1a8ee5c064233e1907c7a2c41250219cb9a191a294b43fc180f2bd3d7854591398d5b3dc5b9359ed60748c638ee400913a396c30d85b643e89fe05f1b37e3ec74d1d7d9cfc19ec58794aad9082521b5ae3c3b7e11a922a2f5b0b95a1d88144589c2c427564da2ae68c89db226af62c2467ad0fcc55ae58d2850d62adfb8f388ffc12778fee504c4dfafb8fd64e7bb957b920b5bff8db7341d1fdd9e9e92707b9ed3d5b37d12132888e43c1d23d0e40a5b32707c2c840de0a7689f55f4966c587100aaf335322c4f133da59fffdb96c66b2ec990156aabcbae40b17b49989d46af11a48d86c21b864fefdb40edd2c0cd147586445c5ac029c74c7b1c0fc69801f2098bd3a1f6d1bd99986b0b7c933cfb4730ab5b419de068f4f526eabc4ffdd2199f19e5278d44efdc0a498f5d84a2856ad64f4a460e3d539a68ae5aa1a2bce770a1072a29197e597225ed5105525472d1014e8bd5629f797207a2526cc01ec8546742132e61c4d885eab9d427f40989bcb392dd3571f25e18c62b99dd4b58fe1a54901e98738357924be29f791982ab69a191c59cb6f25ce64cbf55185e3689d1eb8337b9480da691fddca948d92eeb22fd6ac2dd09d1cb85b71809f0d877a4016ac1a98eb654eaa8fa325f7c6c9057176c0715f28b7a36c74534109d74c2aa403cabe606b116d6740f56ef3f2b5fd0c00f88cb0c72a4aa764593f7c8472;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h90dce1d3f91884b77bb1f651ac2bd3b337b2991a9a14ea672578252b1e90e16dac357f8fa91e279ca7e2734aa4229048a85bf615b51639a9b8456f3e9c3a1afd2e455bd7cc9cea64a7fffc560933c9ba01a37fe3bd7a3a585a0e52ca9c5a0d6aeadcb8a0ef5a6f4986c3b3fa832fc11abfe3691aff78cd45b41b177c6351c1c974132b0bb9c12b279de1305ce3f93c9be61f19c1a9ae9bc8bb89d0d29e3e78a2e4293eb84cb5203fc6f3917f31cbc5130e7d68ed91c82eaca58f65a8142882c77e6f58058b979852f7eff8b3d04b58f464eb1be399d9954e7457f6bc8393b58e38b918c3db0177769de23fc5527ea954bde69ffaec4e57c73c774618e9959a8f449770ced00893d8e29275a4122b32fb4fee309639f9bf769c006c987cfd67f2efb800a172d45f4278d7d40bcb238819bd7b8837dc57afffb678cfc3b78ffbad1e0567dd2d15c58e87b4b496431d920516787da03e8cd9c7282fced216b2c06179f7ce1a95c86c0b9ef8f21577d6bce1fec950cccbe97a35ece5b9f0338a9559f7bb113e03af49874f518dae7cbc16cb8191f8993e3abdcce057857d4755219c03a7400f6b0f4f8eddb1cb5f5dbb5b7c2762a44fbaca8055138b473eb10578fb5ac30af616f40141e3f9a690da14816066b4f44172d04f92ce1666e25c28ed41a879bde2f1abebcf7553f41c3b42d992f502694cf84275cc269b16725311d0c7fcee261bfea3f9f01bd87e317597487491bf845bc93cd4d2e6ef963c9bf95ab6a8c4c298b902c939108a6f5130d2276428fa8bfa0abee91b820af0afd3421ec39426177108f12dc98975d2716f0a20218a858ef0f4a4f6ef5ba108f92ef0edb173e3dd61174e41aa5a361f7415e5a586518236d8e86e05acbc2710b5244ef027fdfc6be4c81ec1abef73f5e522718d1a334e4b63a59eec613f0428426087bd0d47488bc7bb18a4b5e187e2ee923c13c2809d41caf88b30627ba013484aea14b229511d7e3fa78e7164e23ef1d6f52d5357197abcd2f614cc84258def5efce54d24b3ed48f4df8b797f6f49c3fd8bc51d772fc92c93735fe359e2cd376666d28d2b3e872bb40e65fb064b578a6833bf5dce097ab6b2a895654fde0892f21b3b20eec220c6c7ad41957ed2109a6f2f51f09407c786369a04da32cd894f94c9a0275c5d79f354be5300660d3588ab786b23b2155e5ea4b71c6f9d9454a35808e00d5877dd1d94cfeec92931c08ddef72a4f12290ff4392b9e340b6415ea84eb177519efafc732093d844feecd1db1d4fe5b6937b6c0b599d852b87ea55ba3f8b615786759185b38a0ea9f4937cdf40c76d320f51b8878376163a84d2bc1932ff8d9a705883411f61cef5cada8d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h43cfd82813c066fb69bff99eac326c2217d50566ec3d36423dc8db850184a528667e99a43bd99adcd7627bd184796f93f9689169ec0e26060f22e50d3705f73eb801b00979c49df4169780be146d4fe00801241caa2eefb1e37f3fe58aa7e0ea3863c39e6b23c04228b241b4432ba2578f8c92a1f3bd140f1574d7005dbc553564867edfb90461bd311141ce4731dee68822f0a4d621a8975d69d80ae536b3e96abd3b71ee04750d2c2355c73f85bcba91d4afc4ff6e3c9b7bbe0ad9405cb87339cf3c03b3145f2ef97eabf87438c6a3809eaffd95378ca58bb20e81bd4308bff81107d4fca808f26998a68609dde0584867b1c64e13f840585254a88a00267732ff79789624010f645a513f7c77bb8c46799b18e3cc8ff095c4dc5d89fdf6312ae64dd7886927f7d97203a73fbf28d4ac51d1a19da3ed4e37b1aa1d204b6691c7fa0a32997bfb82be6ef4b86dad923f7bf94423b4eb6f5524fd471adeea4683d16566ec95ce5415a2fa3373ebe0950dded50fcdc722b4946833a9e8a545e0843e4b92b87a90625aef56178a9cdca2053b892f3edbd050a24da2634e474ee276997fe1d4719becb03e7ea402bf66904390aa7b321c2ef65f272524c6aba2cf883b1002ec267859696f7a002c2c59895422ca72797caf55b86e132f359c82b9f1aee3a857f0a33dcb811a735ccc55fcadd069490b0a94fc797021da0fc69a656377dd4543abf6b8313edb36c23bb26385b9f19ffbd5dd25e21e159250cb3bcd14c8a6309c0831759d98d382f72ab4dabb2c8399fb0ec5b36b9eff6a2896d5ca1049bd0ddd4120c508992004a7437e1f7e07494be2551134c8d2c547635e47a039b5ff8b4d6afd6e31b2be9aee84fee117a388a3d84a3775c9d7c9072fad97127933649baeafa30da9335db088fb84b10f77c37147fa265251d584e17385d6229c9b28e247cbe6642c4cfcc0137edfed1da11a5887e8fe1646dab1775a4c0f7491d8cd16a2bf438d23532bbba9f699138868ecda32100f94bc99558eb721af1933c3241f12507f325e8b438d697e4004c3343db493879f1dc5aea81f194816f4523e08f1cb20119bea54375f1a550e0a5ccd725f6fadc3eb5f69fded00fcfeb6d46283295a78095556cb943ee098b422353b212c33c362931482be1c8cae040f0e7688b02fbbe32cbb1d0e599773ada0945203575bfc846a15a19a82f588de374956e31f901a90a082a84ecf9b1ce72f2e3d0f293e3e445fad4dbf50040e1f6af6d41188fc96c9bf82cd6dab2f63aeb2f0bb20f775473e01515b3f9baf6096af423ee7752b7330525042243439928e63e2aa39e6298332648ee7e6388d197742c4b9ce0cc1f8ca02862453fa10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h518bd0ecdaa388c147a3b4182ce46a9641b4c0a07540bc09759cedd26000ba6e59e36e778910dc72d2cc5801282ddb18d64c264e2240f032421f571349c3e1d834f7633f984589af887ffc46bd7cc05c509a9765699cdbe9c46ddb54e6d56b9a052778f6f4f3d54829d93a73e66001274dc106cc9990cfeda40589d23fe5b33116fcf4c31c9919e591719d58c7de04832bdb86be8569106b9e8bdfaad8dc27ce9d923379d3911916140a435bc74046d504b5e1c31cdd6642fc98f6c4af368b7918c9bbb2c96f3653c6d800f7b6953323e82bc5df7c4f602c4ebc84d41c399a6aa34ef0ff07ae870ae904561fc39c93c0c22ad98215ac71c81ee724088d6662bf468474ae66d94799530bea024ec92261a90df6ef129c8fde9316e3ecaafc2c4029efd6fafec589511bd16b87977eda1b5b8e7a973548cf7c5949d9df26b49fa6328bab7b8d68fb90d12982d23341d1e61f903e377a61109412bdbe17c24972d51385649a79d168b1072b7fd02b9332d4e5c09b48c5f1f625606f5cbd2e117c605f3ee7bbf9d1995dc4e27b09293aa01e98971e1dbd89f9030e4add3700a7823baad8ea715d8300ec6c3de975bc8b206fe2595b345496831d0c310dd786f2ec067b9a3b88e4d431d259da0da90aff3f7e16ac6a2e6d460bdcbddca12fce4e5b4842b1d6d4f2ea060d42b465a78df91a087f2c783287e1b28f5ad6f6fed5d371af10bbb306f20a3349761232998b9ce21ff84c62b0fc5ceafa0fbef819a452947a9cebbcbc2a2be9a6d8bf6098596091401384b466c75c1d357eb4b73f9898669734914c2752c533dc2cab6fd64eb4c379b0c09df6eba824bf88eecac82a09fa5d6435351d333e117f4fd9f757a8d99e0e78b5734e386658a397590f33e208e98e90f2caef19e68c47dcf5e50325a00178d1ff598f5867eb5eab7116da5a7bb333ba269d1e2eba0a0eec48f09145e8e94e5279e59be7cdf2320d37d5c8b0b3d19a8f1ca1b85489890cf7085a184fb75ea9e3b5a6feed34d8594ec6e285bf75b762a8ab3c6550894fe389bd51e9e21ad984438bfb57962270302b1e60469bb8d10faaae3db92af0ee5489fce0e36b02d96d3fe988f7f4838c02b86a3789a7c9f84dfe643e0202d432fd9a58bffdf586621f5e21055c9b5994010040077fdfb1ec0238bee3d8b829d555e0d57dfbd4f1d700fe0900ada8c4df62d20fc272cba32f31e1a6ee4140ecb7da24a5c71f935092b783516b2603862a86929ef241de92cf75756b2d2768b71a7f1f5142ae4c32ac34d67ca17db797e70a8c68be9b6124b6aba8c8878ec2efd0b87ed48179b3e5fee42fb689444ed6e2d6c74238b1111f4c01385c78222f98ef3e49d5ea6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hfe67053ac26e000f968cca737d1d18c07c77b45860b130ff383eb932820d8889f9659562c54fc4b689c2d7d2cf0e38e38b84b2bc5cde8cfadd19d592ef0955bcede3a788ee07f5df73bc394125db12af10b4d8df0c890fbb65ca5a89a3c28122a1d386ddbf2461bde0ceb02ce2826ab4aabcc5cbb05284529cfdddf1f9a917775f176890fa7233985e9c537ab2af072d9cdb19e0c4a79a4af0e202833bc7ec8c53a144c7daf20e425501e5c4e5b6a619eff0489d3f9f5a1f85520d4250628d7385b64109ba9749bd273eb46c385e2c8fbb37b799cada0730f2f34e55d5b3dbfdd1adb630d2bc6fd6c45779d96cd6dda70a181fcc91550b2b49d5bad7ac0b649f3c8bb3a3e4ebb58eb2eb0d5123011ec378cb06b860d76a5df86f61c2c13991e4d75abb359c963dc6468726a1292c7c7f7f355f1584d73d101cfb14072d7bac2f8b5be1463f7fe7c4e5f83dc239ace26fa4f27c6dcf80947bf1344763b79ee6f2db7df8d8b1f15201248f7edba548951bef57b5dcde9eaf043ab5340526e38dcc0d916255cb81d9b932dfd6335798486f3f11545b71481f5be720056526543bde66d928b4c4966c8732949c73812c339aea723337718ab79027b6a55727c108dd88edf8e446ef40264dcb0ad76ce049e5a4b65ea6fe87d3d3dcbcdc8ee08a5a7a4568df8d607c71de08b7f83fb878f80b23b66ce8663efbbcc22c30d93c43abee8025399eda354be0e471820a129919e1f72c33a4fe675eedb9e349f703e38e7fda12f819a995f086fa991f4e6256f43df06f87c10da1ac2eb7946a019b504ffa721d9f1baec1b35630423b1f126840fc8c53c8734537c19cbd884587beb85f209305fb1c0e4385e6e18535a212bc55461708cbc2adb49947a0970c1bc13649e3d120bf0ee6f33b75ce8384944b1ce9136db3063ac7501aa5877762d27d926b96e315089fe248c908f9bf14bd7f7897dd36674e5776f5d028d4395f0eed805813258737293ab1404dacc4861f7bcdb08163cf4dba2e4ecbe573de4e4a8ae93a41f9af8b8c2a372c0ed35af31d985021fa78842e97870435a70569d1eb97429fe218ea7246449a3ee5bd35d7c61294b93f5e0ac0659025809d0c208e8f1dbbcf348e71ac6d0a035c671212298e9d163a15aaf58ddaa922086d3f5cb16fb7eeb5d4fca05228f65c2831f69355c0d83ca801c3b16f88bd065d6a30ae8a792fd1b73144002b280a17d099a30d694db6bd324e6bf653c3e8fdbc514981c0fce7c15cd62649526a82e32c14e6ff267c3d3cbe81f39800683ea01ff08f2b33a53858c8d8ef34ceb3fb086512fd857460481c07ae55e703c5176acad810ff07a84e99cc6bd86c04ceb03fea547707bed6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hbdfcd634e45550702932a0c0921d2806a6fc102514e9bee9a0eee62a2b56e26e3f9375f809de33bc25d3feaf58f8b20173ab87eff6ab3f1b90ac09f307163d9346a97c6cfcec42d96f47499d13efc4720ec20762b26f49af2e6e249572b127a3c630b000e6caf120dc5b8a6cdb52f2a02447d7706f4a943e6899dbc157e268af552235e90d3583b637757e1a76ca1d1d8a10484751a1515881759964a4c880cb54542f9c56bf12b0699c46cd00b91a15435d6028db1032693df593b1eab420b0e55cd1d5780c0ef8019b258b49b45bbafd5224d3a81e7902d28d0c555140caa25003d5cde13a2768d88244aac1fa84b477a6aa0b473dc068ed3efea63a816abf8c4cca2ea677d8bd97629ead2af7562203dd85197285ecd67fa4338d898a2afc92205e6e95ba594778cfcd258854b9be7504f2849f4fccce20532903a54e66c98feb63825ce0c8addf02658d4a590caf3ad97b447a920a1ee7cf67680076d87e11791895b872058163099688daec2acf9b0496205f5325fdea500f4fbfc532488bb3ea6c0bbf2fe851e82ca0eb1e9554207b2854e5a9252f8d0384aa1798d7711b55ad2a8e56fbc85daefa33b7dc570a671ae6c4936e5a7f5e369eebe9f6ad6d872bcfa97f802f119284381e8af15aca49f5b8591ed230f6c5532581b284c201325398d95b84c9f3560a27e2359cff93676e3ffc7440fbff16f67b84309ed3993689b532c3e87c2ba10457c1702f1ffa8acc74c6b3db097789d403c22e4ba1ff1e9ab9f0a7ceef05cd98f6d78e2085f4cafad1064f87ecd2579bad2b7eced9a49336fa6f3b2a82425152c27663f3104232997db308903c6d4c4e7421df9e3b8642cae611f2f6fbb8173d5bc5828306d3d25b950c839bcb4db45be365d27da521bdc0b7814f8ca31253c020e2330014b915b75e75c16533d672c076c41a560a00763fb5d62b6c84608cc921a6dc01369dcfd17da68511d12e854075f0eca7c60a0e1e79680fd8b93aae6d12136d5299f6bd0cfa79e886880910d221ba76bdcdd4720642672a22cac801f5c83dd66b90f074a722ab0bb6f88c3e588ca4537baec6c9ee15eb064487f72d05dd570026f63c3d3cf5e166d73daffde74b75ca003c9b1a1614c401cb35a9220339ad6d4da92370e5aa7dd54b83f1382b19939b8200f790df45558e8c677851b0c84d8335e9d53435554cdafa971550baa818be98b2af1149220c4e2d22bf73a16fa5a8dbf07b7e7f287f0fe87fc018fcc4e8df882d6a05359d8ab9376ee8f2625dfe5b3ee8b3716c0c348596337f7fbfb5f5c7ffdaa00662e3c879ad2bc2ca5aaae475eb4b7edd411393baa833873797f3eda76b3afc4c9238f62e6f1c2995bf7180;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h964a6c1c64e547cbee56bc101c8b8baf1f864acf68553a03d5c72ff97ddc158339d940c994d5ed1bbd2eab85d160b049369053473188c6e5446e576522f7579cb9d083e7a7f6bf51050e63d41b0daf273573716904d58ae60a53e8d27c684e942626b46540f7ab4bc99847c02c3f6a4e5b71ba09162a90ed9a8298a073d6f16a85acce8df76fdcb036846c0ec366c37c45be606eed10eff13f0ac97ce1ff77388aa2819769eec19a4a37b066b15a8e3bf0da33fbf9283acf090f255d3b543e65daf8db54de3c941dc5ce22091f97924e15937fbc97b8afbfdb6a605929428238b087d441232bc034fd87aa16c6c344d674a53d5f0289426e36882b0cb431638a82081f7b8b6a51e08a6151991ecfa1129526e37f5b59a7224889ac3c3eaa914967db779a2dd669717d65632c8ecf294252103b8051f280653be11bc3b885bc61ae6280a558d93f5673c901dc5e1ab8fdf11c622197f9c90fe40dc68a64f62c5eaaa40c6d83b55ebe2cef0d0da35224e39c0c4086d0bbe42c4d13e4751288410be62b24f74e0c74c4ce4ab5ef91c2b3fd9c7f7bb2969ff60bd6dd060c34ca42eb71beafe344fdd497421639bc49e8fd3250cb56d48e9785caf2b0e9f1838a6e88ed518ab36570a8fa062b0861e63b744e5c77f039b8d646f144c1aaa7049c695dce7db808e0c91a2afcab66efe393c63f2abde18631b344ef0c841293ab30ad8fa7bd7cf7fb01348b1798e1198d4e2e42fddac7d7da0eb8f1251cd73f0daeaefccbd3cdcb778e6e7081c11eaf1744f318d3ebfd23b2b2fa7c5df9bb79e565dae29c636a55b9c640c5fd408759486c44d68afaa0babf0f83b1eb65f52164c2faa2a7e2d957241eabef0aa509a5da9eef67beb921c1d51bbd77832f88b5c0e7e014f3ff542bbe238ec9525d9f09a0e71c2ffc5b7553e0852c22d6c750c8910cb5972dbeea14e3fa2f903758f8428f7d7504ffd940f6f7c71a658c2b9b3f185c0704edeab3a4aa4d7534edfcb2725674ff12168cd62c11d2b16cbf17cf3aa0f95d7a9ff5f0c3f3f06ad64e2620ec9676818f73bca3fe2310c13a6570609acc574db052704aa40e2fe404e6e305727a2dd65f063713cc9e15ab0b78c0d3737306578b926db1b1a755ff66a7f67e51a4236a9b9bdd9426ca8d681b8c6e62ae273856ed78df304ef0b45ee87c3f9f507db3af68c799025a889e7c6341380bdbdb8da7527ed6e748d35affc62d24798e00ea77f3606d757f6ce9e6496942b1403e21403e7e57f7228b2de06204199992d270bb91b5ecc4ce4859b56b6e60aaa84bb8d4dd4d2b4f784ceb5ad873a899a55a2a25226359a17f598ab2163298f2f00d62b341eedda80aab69908c479fb7bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'haf29fad7947f2e7e1881f328b95b5f057560e07a6392379a6c81b7d2a3017eeec148ae27c68a31e0abbcfe76b7f42d56bff2d446e681c1409abbb53162eafe49efe40b4c1473f1eda047e6883acedf2250fddf9e53cdf59d55659eb3bcc5b2c6bbc6a60afda0e2e17f0625e99719ccf64d4c4b1b563227d35eecdae4604ce511158dd5afad37095595fd5809ae8d79393840d9143013b268e797faa574493fc024801929ded2b2b1b479dcee6ee1c7a9ae85320bbdc7bf0d4fa68ac94ae5950e013086eabb285500eef8daa506e817de4149acc06d4b8a3a4ae48696eeea9caa20f2ad146f91e1be170e154f723ca18a85edcafa4cd95d8eb3fbac73258cdb4b87e85e52544c329fcfada75adb4ee3e7cf01cf5a37f50a497b52ae10ab0efd564b288ab1babb31d7a0f10bbb590f9a7fe51af3cc2968150f7bea19e5d41346bd81617e40502c6eabeca90ea101d17f0d710f5fdd4de906d01cbef98ae9a9b69d420d4dc231ba633f5a5da21a6f5d7d69e2005b64b63d2fd210be781476e643697a14bf12868602a3d405518319054a0015b588e29492171f6a32062e882b52eff1016cbc92238f42ed652012f650530760f769081590808618f0242fc269d687158553158fe286acc0ecd35548cb08d42ecf4b4604f4a2cd4894b9cce0b9f064462d4c640cee05f1e4a96eff079bdd25adb54649f8a6aa08ec77a9908c802bf89bb96d29bf0770d8b7cbfc78a3d7cb00c975a96b7a0ff962c6e90adc6356d89acbd6cde9e91503f01b726a4e775071ca02b7341d345140aa554369a7f63c39ab769a0c026fbfa033fa276dab0febc1cbdd0ab01f859e66b3eb8b8a9719785b371fa693c49c1236ef870abd972308bcfa6af84d21e962f92d5f11be574ae51189ad91ed11a526dbd072d552c1a8c9b080bb5490f8cafc2ed0e0796a57af04a73b613d4af329825d0a9a7bc7e59464758b1bd1a54e9699d0742389f08e584e1f46f00712e453a5c93be2b03d0da1e5783b045a8a56840ce67db4c613e775abaa987bfff7a8f4c457f18a790f2b9135f62c877b7804a1e296c7451a2910d975e3c4c81b406f378df14ac895e86acbaa11e755bc5f6649e95319a834b3638b7497543340f1086818df7c102eacefd7e2bb6b3f99f611cbef9b7aa79ff30cd874a13555f7e11aa9d8e4b578340929f60f9668770ffdf0f9befa8759e4e67f6502ead31b4ea63c95eb808c8e61f29bea77f641d43072bc921078d993ab606f1c2287c350cd8f94e535b3a6bcb65f303408c2634d4699bc2882f9f4dbc66fe1d878032b5feee79948985303b09dfe3c2bc9077f5dc681bd917f8ad15f43f038f054db94c207a1797370f1f8c4b6ca8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h7581f3b67aad88043cb223c27249cf32e416fbee438ae357d03017eb7fe91e7485bb0ffd115aa8d42e73a323418b7babcf6c3a8033224ed299aa5d469d1aeb650d2692273fb11c4888034d5af42e5b380714360c818892b00da79d930e9c6939b7d28d64fac80441aacdc51893a980a1e85fb1b1eff1d59eef97cc1e27732863e3100a34a3b80c495633331c930dcd56261980277992b2aeb4d028d8b7808ac96c6b68396c6ff050a406278cd912329b3e96db1fb0ba4f3b3f686cbf5e32bda98e0ea373b42f009a821709132169af9ade179187814864273199b707385f3cf772c05037ec362c1d32742f53135fec6e5f9b4af89aed1505deef09e24dcaebb15cb0278656d540e5d2713b8e7ce9fd6db05aebc24fda2b027ca5b271b11f3fc44b88618ddedbff125142b79d8102a36e2a2e8e6290560103c80fda80438509209d09f320ae9459fc65af755bbad86de8deb2b2653ac86d5cd1c51d8f0ae725d17f3f22359d58022291238d2749ea744778f5705c47af3c1a50e2878a66e8bef9912f78bbd5e9dda1da67d5c5cbbc302ea21d7cc28af85ff97f4b8a1d92035aafbbf28ee622df8cd585263d7bd89a32b8649d41b7aa33465f460a8d44409f7b4f9e6cb7c9e7d0a2cfd0693befc6fe0c6ccb43ac9e87577cb854888e4772616bffad9e4565f536a54cb76340337ff230f95a75f0b5c8ca3d866ed12ab0921484fba35106123f80eae84b8203b0fc4612349de053fa0954b9ca54570e4fa703238ac2e7d4255843be5f45f7d9f45e8be75acc3a109581661303192399a29584aa6ed8424df74449540f9d832c370fc441525b5c3c6f76b39590f2d50bc1ae945ae20956ee042856fa122edb90ddbda13cc3e9ce6243289f0a71130706e2cd88e96565ce5fde8dd636f3dfa8044b330742c3ac6e826a6a94417abf3eb1c4262f5155728edd231003b6c27a67d967beff3ef0510a2e05bf390c9832e1818e013a596580256dec02f54964d2c297a09b0975a2e24f791f98c38dc37b103f7e4c8eb3c0e2c663c34f49a4bff785da393ef02c5e8fce4ab200dc64e67e2794f81a4fd5317d2b6a642bf494f046f0c1284cba5f20e73a2140055b1c902b81922a8b101b8c51ed83e6ebccf822c82a73c1efa84776b28260c146ce66d7d3578719e14e2251e1bccd5c50178bce0037b031d7a26519c2e427c4a6c9690769728b0fd3e1c0c594bd467200c5d2cfbb1bd8885d094e99e4a1ea69f886b2905d39d5673e71bf62f13a30d29b1afcdd5b8e65784dfd1b8e962810b46e21b2d6d381c245ee3ff53920e2113e01a5265ff9c8d26f7f88f734dbc0364dee0b8c785141b51ab161e0218f97f448c938420c76b0ac95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he8d21594fc67da0ba52e699c0dc82275d28498c8d15f67886001bed67cc58b0de2bd36afe6cbbac166428d8eecfed7f944724427e621590ab09785ed68e8dd735e6bbe8c2d2d3f634566045488df4411c469aec9c664c21ea0dcee352cbed9ed3f9ad7e6147f7e6d437eab3d09b96e3e13eb0e340dc89fd28fb21ad086f651d6482b1586dd4cd4dda4e7fd2f2157c1f9f31aabcfc134432e7e2ccc27dcff9920d076a5bfa1fbc4592bcb58472160b27e582607cee278649232b3f5803a42c874722935835b1e600f742baa8f53facd0261cda087406e3cafd07fc219b996c21f5e16c53dda160f482d72b786d3bc9f3fa61c6341215197e668dfc6e140f427ab6e14da99bf59d4c65c9af282d2a49c14c1d28aca60956ba9f7ea5e1ea6cc98f04c06d52975ece962163d4e0b01fc6b370a4c5e7f13201c0ed455393d3ceec7dcfd50c1273a2228607d3981d3b4096e46bb294df84c144e62108fa0f564ee79b606394c99c1200bbc77330cfbc0a4988c1b0cd43352adc0ad29b08e84e907c94db40e11c623b09ddb1475341a2d5761c91a3cf6fafcc40919bd06a0a011dfa865458c49596f1de87d9292b3060c0e727ff22a84d77dc138241de46a1ed0ab07954867f95a8b08364de73db865b1b754bf0b5ba6b27f8e48fdf650b3996020c3581f08baf4a475bcd94c3596e44c716a30ab083774f0fbd69d1e7e97311a5eae3c3eb22c623fa586a45710905e0299da8019c8c2c775ee8792f56dd50e20f75fb57c935b76627e0db1909b653ad5d43881e908e68b8ec707118855e2879e214ac871c2ae81e4964469cb05897d061aaa6419842c6b4c21f44a3a9641968aab0ab35c8d584783dd9964187a5f858f4bdc45aaacd011ba213495de6673200009cfe27f12a78d7f01c4ab30b86d7ad662fc1fa6bd3b4732f21872b27b8a0be9e465083e0b36228e3c6f8b1b9f64902637f1ba566275e78199b371fa2e6ecbe652edd95fac377105236fc349104f1a46ebbee7a5e8da1af29f802a60050f80ded0cc18842346fcda2a76f33a89577207960e75b503d0ce530a2ce4c4fa4fb8b8f105178202838abfdb8a6b748247cc340119f89de5d090b24916cb7293865532173b6d98e2a8b98b0e09e5ebd20da666f40f6edb64b02aed1c302cd1c9fd806a92737fdc8417554b1cc9afd3cf5da571fda5e145c90a9884c791755afe2aa90e7053266f348b1216e9d4a74aedd493817512b9317432dc96e7f113c5d3caac8466768a3897b3dd4676603883b88ad4490e7d0fc39102b8676369a1faa9fba902d2bde84aa6147b2ee935080c862068c90c1a04ff11d88425635a8889e83ed72a77a37efe2eb31cb5f698e25818c2bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h7fb31c381e98a88f819cc01f862eb921be68422b329496e9041b3b85a002e6a83673c762687406e0a72c89d47cacbb822c530c5aae7d84789872c36e8141faa2e1447693bd968b38eac311f01d4fc5b0085bfdff95f79290c22e3645861940b1ebbed9acd084d83db5b41f2c0b27df100ab09355d5ed885822aacc7a7ebccb8c63297c58cbe7915a3e10e1cf301ab979411f46165024d9a0a3ff74d85744490c2a6530554940ea8570325590c2606d3cee7f0bbf31b45802a6fa076caf361b2d446d62d9a974f12a71b11520b4e18e21316bf0928f4c71e241579287bb490c5be3ea16ca3c73039b58c9e9b5dbd03c2b469311bb49de941c79ce5787a087a97aa71e387e67b2ee3d038c357226d6c7171c53e1869b348cc28e7c9ea789f2ff2ac82343e5c9657395ca33d425641bac1eafd0b306a94f2efb417149be01ab6075217ed92d6b98c99036f5699c76f623c4f127907ec6a3951910254222606db4b4451f07ebdcaaa8981c9212f02a3fb45b484de82e4ef524c95a2d391b29f7c4d1b4886a0b979bbc753587c13a02b4ca337d972355966dde5c1c71a545b3cb5407dcdb9f45741fcb5f094ffb73e5adcfdacffd32122f85f90c993d044eb9447ad3fc7569014fd4274c710781949b79dea55848d328a9e2d7cb9e6071cd4f5356ffcf358a89fbb50dff6ff5192d94a52f6c59dbe1e4b801cf6a46c2d2445469fff9d66b6155e5a3e692cad9d9ae6eca2f931480747042721beaef4c01d6ce905b24a5d92615ed5e65551e38a2de0c96849cc670b9f6cb40027985cd2a58d5c95a3419ed2ffd6574d7306eb1bb2dd3fd0be5cd5aab90b3506448096af4776632a6b9737082157b19033594ee92285c8d23c341a186c3857cce289570e2359e8304a58d39518792dd0d04aa1a884a9a27177ff413cf526b030fef607d956cc37982e2dafc3255ae2383281c703cf70591e54eba6433142feeb783aba0541418c9b51ed1e7cef452a0aec9709afaa5ced8a5363e4408ad0af98572c4557904e75275e8c6404633c0bf8874241a90f0a7b220e9cc1dd90f1ac4132c071010735ed56827bbfaf61778e8e6ea5809c4802274eb3ea5cffe157ff54c71c31bdbcf3cb4323c2c1e73f676c4de57a24c7d8591fc3fdae55862a9764585223feefe6f181707571fae8ca48e99019c03fc2b5ac2b417d8ee04b2c6ce7bc4f22895b8f9b9a832c3be7505db54b7b285c99124a8268618e3804087870cf63f16295f77b57c8106886d03be7142bc52bd156c2cc4895c52677421b10eb7a222b93b4669b5d4bc07b944572cade46f839b73e8c3ff2329fb65416e6f42bf37f6e2ba2e980c6116af5808602e2ab9d7b11b184deb6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he2a897ad212d0018132a51548f3589c33afbcd522dc8924550de50243190e8dcc638835d739584a251d059fd1e31b06dbce641e7b682078df663680e10adb9d4f4bf62423d60305a48d143ddf653bc2be1e380594adf34df6c69e225d98ebb0a6f89b7a5f1ddeba99816fa0afd221124b6b96712d5c9eb0bf4abbe36a9c8537dbb5380ef0aa022901329fca7ea3b4c7df97159ae22677ae8a3a59ff6558383ddd6a895652365f7f981e28164a640e39a28a0cc3403ef41b6065d50584f4c1b492c210fa8af79103be8ad4af577e2cf83cd4f3b078c18ae0274200745509469bdfde1bc932476524c2608fb8de3f63492d6b101fddca6aa7c76ddb29e6e5bf716017fd326c26124dd1baddf45d0a81abebf57341848dfb24fe42b721a0853d8859e619c856fd2a994487366db37c8d856e39caa9a7cce4ffee873e769ef1e52eb9b4c61c58b7341f42dbc2ffc742248ce33e2e0848b7d467150cc73280b05cb8e7362f1a3ad56501d571ab276b538a06f19f382b08ca5ea1c3a664b00ff34ca6c4bc121e849da81cf414a156e1110f2cd69d3e781ba1a99f0ff65b41f8567fe64341f60249cc76a243f0a4ebab33af12f4f02eea9ae1ec431f779bdf57dbe7adfc7ef8b695daff35435d44f900e00e8495f1c4ef787c48d1670c07bfb16ec25f4969817e6014026cd8de7372f6f401df964cf272e980a658f286e9d196fab883cd075d23e31abbaa66c60a60ab7825e2da2c49968160501a295f6ca1ddcaeebc1b0a243b091eb9a76680b014967534e7446513f4a5a89ffaed3e6aa43f087588892c065cfe574da6d096d664b0f1b6cc1c63463339a3851882950fd0b64399f24ccfc0bc2f20fabb7d50d0e9a2259fd3d4c17086cd0d6becff0cd1a7500cec5088f631c1a15f1620a090de784b04ac1c048afbf63a16766e1027411322d077b53646c0c6f9f07080dccda59c45d210efb3ce99f3d71ad5fc9d5543069a21ee4002c71d5ececb1dc4c490ac3217503d0b2c7148a060e4942e9974eca0ad262829f593a757ec603e310783ac37b8cada610c8fc3ba28029da5a5d289de794937505d48564d7ff5439c8360dd851d66e088d84a3df2fa855296a83ccaa27ab91ebc36d88a8aa66d908ef26d538e7081efa88c06635a6242f83798b5623a93c104da304b8714c0b82aa130e680c20b72baa0f58e717176950ad78283591ad3ed2dfdaa2e1772ebc552c131dc0ff2a104823d68a911d9f1517b670b55c7cb85e70cdf0aadda88d6f3d2eb00587062df63b216ac384b67ad3d753295ae76775ac8549e2d7ed248a1be3855e3d18df455dc1659b9c327ee483e85a844c2ec7182edfcc44741424b8d5f95e87d37bec5;
        #1
        $finish();
    end
endmodule
