module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    compressor_CLA32_12 compressor_CLA32_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA32_12(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [0:0] comp_out16;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [17:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [13:0] stage1_4;
   wire [14:0] stage1_5;
   wire [16:0] stage1_6;
   wire [10:0] stage1_7;
   wire [21:0] stage1_8;
   wire [28:0] stage1_9;
   wire [24:0] stage1_10;
   wire [29:0] stage1_11;
   wire [2:0] stage1_12;
   wire [0:0] stage1_13;
   wire [7:0] stage2_0;
   wire [10:0] stage2_1;
   wire [1:0] stage2_2;
   wire [5:0] stage2_3;
   wire [6:0] stage2_4;
   wire [3:0] stage2_5;
   wire [5:0] stage2_6;
   wire [12:0] stage2_7;
   wire [5:0] stage2_8;
   wire [12:0] stage2_9;
   wire [11:0] stage2_10;
   wire [11:0] stage2_11;
   wire [8:0] stage2_12;
   wire [5:0] stage2_13;
   wire [7:0] stage3_0;
   wire [5:0] stage3_1;
   wire [2:0] stage3_2;
   wire [0:0] stage3_3;
   wire [2:0] stage3_4;
   wire [5:0] stage3_5;
   wire [0:0] stage3_6;
   wire [8:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [1:0] stage3_14;
   wire [0:0] stage3_15;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [0:0] stage4_15;
   wire [0:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc615_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[0]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc606_5 gpc9 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[0],stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_6[1]},
      {stage0_7[2]},
      {stage1_8[1],stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage1_8[2],stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12], stage0_6[13]},
      {stage1_8[3],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage1_9[0],stage1_8[4],stage1_7[4],stage1_6[6],stage1_5[11]}
   );
   gpc606_5 gpc15 (
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage1_9[1],stage1_8[5],stage1_7[5],stage1_6[7],stage1_5[12]}
   );
   gpc606_5 gpc16 (
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage1_9[2],stage1_8[6],stage1_7[6],stage1_6[8],stage1_5[13]}
   );
   gpc615_5 gpc17 (
      {stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_6[14]},
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage1_9[3],stage1_8[7],stage1_7[7],stage1_6[9],stage1_5[14]}
   );
   gpc606_5 gpc18 (
      {stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[8],stage1_7[8],stage1_6[10]}
   );
   gpc606_5 gpc19 (
      {stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[5],stage1_8[9],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc20 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31]},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[6],stage1_8[10],stage1_7[10]}
   );
   gpc615_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_9[6]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[7],stage1_8[11]}
   );
   gpc615_5 gpc22 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_9[7]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[8],stage1_8[12]}
   );
   gpc615_5 gpc23 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12]},
      {stage0_10[12]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[9]}
   );
   gpc1_1 gpc24 (
      {stage0_0[17]},
      {stage1_0[3]}
   );
   gpc1_1 gpc25 (
      {stage0_0[18]},
      {stage1_0[4]}
   );
   gpc1_1 gpc26 (
      {stage0_0[19]},
      {stage1_0[5]}
   );
   gpc1_1 gpc27 (
      {stage0_0[20]},
      {stage1_0[6]}
   );
   gpc1_1 gpc28 (
      {stage0_0[21]},
      {stage1_0[7]}
   );
   gpc1_1 gpc29 (
      {stage0_0[22]},
      {stage1_0[8]}
   );
   gpc1_1 gpc30 (
      {stage0_0[23]},
      {stage1_0[9]}
   );
   gpc1_1 gpc31 (
      {stage0_0[24]},
      {stage1_0[10]}
   );
   gpc1_1 gpc32 (
      {stage0_0[25]},
      {stage1_0[11]}
   );
   gpc1_1 gpc33 (
      {stage0_0[26]},
      {stage1_0[12]}
   );
   gpc1_1 gpc34 (
      {stage0_0[27]},
      {stage1_0[13]}
   );
   gpc1_1 gpc35 (
      {stage0_0[28]},
      {stage1_0[14]}
   );
   gpc1_1 gpc36 (
      {stage0_0[29]},
      {stage1_0[15]}
   );
   gpc1_1 gpc37 (
      {stage0_0[30]},
      {stage1_0[16]}
   );
   gpc1_1 gpc38 (
      {stage0_0[31]},
      {stage1_0[17]}
   );
   gpc1_1 gpc39 (
      {stage0_1[31]},
      {stage1_1[8]}
   );
   gpc1_1 gpc40 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc41 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc42 (
      {stage0_3[30]},
      {stage1_3[10]}
   );
   gpc1_1 gpc43 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc44 (
      {stage0_6[27]},
      {stage1_6[12]}
   );
   gpc1_1 gpc45 (
      {stage0_6[28]},
      {stage1_6[13]}
   );
   gpc1_1 gpc46 (
      {stage0_6[29]},
      {stage1_6[14]}
   );
   gpc1_1 gpc47 (
      {stage0_6[30]},
      {stage1_6[15]}
   );
   gpc1_1 gpc48 (
      {stage0_6[31]},
      {stage1_6[16]}
   );
   gpc1_1 gpc49 (
      {stage0_8[23]},
      {stage1_8[13]}
   );
   gpc1_1 gpc50 (
      {stage0_8[24]},
      {stage1_8[14]}
   );
   gpc1_1 gpc51 (
      {stage0_8[25]},
      {stage1_8[15]}
   );
   gpc1_1 gpc52 (
      {stage0_8[26]},
      {stage1_8[16]}
   );
   gpc1_1 gpc53 (
      {stage0_8[27]},
      {stage1_8[17]}
   );
   gpc1_1 gpc54 (
      {stage0_8[28]},
      {stage1_8[18]}
   );
   gpc1_1 gpc55 (
      {stage0_8[29]},
      {stage1_8[19]}
   );
   gpc1_1 gpc56 (
      {stage0_8[30]},
      {stage1_8[20]}
   );
   gpc1_1 gpc57 (
      {stage0_8[31]},
      {stage1_8[21]}
   );
   gpc1_1 gpc58 (
      {stage0_9[13]},
      {stage1_9[10]}
   );
   gpc1_1 gpc59 (
      {stage0_9[14]},
      {stage1_9[11]}
   );
   gpc1_1 gpc60 (
      {stage0_9[15]},
      {stage1_9[12]}
   );
   gpc1_1 gpc61 (
      {stage0_9[16]},
      {stage1_9[13]}
   );
   gpc1_1 gpc62 (
      {stage0_9[17]},
      {stage1_9[14]}
   );
   gpc1_1 gpc63 (
      {stage0_9[18]},
      {stage1_9[15]}
   );
   gpc1_1 gpc64 (
      {stage0_9[19]},
      {stage1_9[16]}
   );
   gpc1_1 gpc65 (
      {stage0_9[20]},
      {stage1_9[17]}
   );
   gpc1_1 gpc66 (
      {stage0_9[21]},
      {stage1_9[18]}
   );
   gpc1_1 gpc67 (
      {stage0_9[22]},
      {stage1_9[19]}
   );
   gpc1_1 gpc68 (
      {stage0_9[23]},
      {stage1_9[20]}
   );
   gpc1_1 gpc69 (
      {stage0_9[24]},
      {stage1_9[21]}
   );
   gpc1_1 gpc70 (
      {stage0_9[25]},
      {stage1_9[22]}
   );
   gpc1_1 gpc71 (
      {stage0_9[26]},
      {stage1_9[23]}
   );
   gpc1_1 gpc72 (
      {stage0_9[27]},
      {stage1_9[24]}
   );
   gpc1_1 gpc73 (
      {stage0_9[28]},
      {stage1_9[25]}
   );
   gpc1_1 gpc74 (
      {stage0_9[29]},
      {stage1_9[26]}
   );
   gpc1_1 gpc75 (
      {stage0_9[30]},
      {stage1_9[27]}
   );
   gpc1_1 gpc76 (
      {stage0_9[31]},
      {stage1_9[28]}
   );
   gpc1_1 gpc77 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc78 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc79 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc80 (
      {stage0_10[16]},
      {stage1_10[9]}
   );
   gpc1_1 gpc81 (
      {stage0_10[17]},
      {stage1_10[10]}
   );
   gpc1_1 gpc82 (
      {stage0_10[18]},
      {stage1_10[11]}
   );
   gpc1_1 gpc83 (
      {stage0_10[19]},
      {stage1_10[12]}
   );
   gpc1_1 gpc84 (
      {stage0_10[20]},
      {stage1_10[13]}
   );
   gpc1_1 gpc85 (
      {stage0_10[21]},
      {stage1_10[14]}
   );
   gpc1_1 gpc86 (
      {stage0_10[22]},
      {stage1_10[15]}
   );
   gpc1_1 gpc87 (
      {stage0_10[23]},
      {stage1_10[16]}
   );
   gpc1_1 gpc88 (
      {stage0_10[24]},
      {stage1_10[17]}
   );
   gpc1_1 gpc89 (
      {stage0_10[25]},
      {stage1_10[18]}
   );
   gpc1_1 gpc90 (
      {stage0_10[26]},
      {stage1_10[19]}
   );
   gpc1_1 gpc91 (
      {stage0_10[27]},
      {stage1_10[20]}
   );
   gpc1_1 gpc92 (
      {stage0_10[28]},
      {stage1_10[21]}
   );
   gpc1_1 gpc93 (
      {stage0_10[29]},
      {stage1_10[22]}
   );
   gpc1_1 gpc94 (
      {stage0_10[30]},
      {stage1_10[23]}
   );
   gpc1_1 gpc95 (
      {stage0_10[31]},
      {stage1_10[24]}
   );
   gpc1_1 gpc96 (
      {stage0_11[6]},
      {stage1_11[4]}
   );
   gpc1_1 gpc97 (
      {stage0_11[7]},
      {stage1_11[5]}
   );
   gpc1_1 gpc98 (
      {stage0_11[8]},
      {stage1_11[6]}
   );
   gpc1_1 gpc99 (
      {stage0_11[9]},
      {stage1_11[7]}
   );
   gpc1_1 gpc100 (
      {stage0_11[10]},
      {stage1_11[8]}
   );
   gpc1_1 gpc101 (
      {stage0_11[11]},
      {stage1_11[9]}
   );
   gpc1_1 gpc102 (
      {stage0_11[12]},
      {stage1_11[10]}
   );
   gpc1_1 gpc103 (
      {stage0_11[13]},
      {stage1_11[11]}
   );
   gpc1_1 gpc104 (
      {stage0_11[14]},
      {stage1_11[12]}
   );
   gpc1_1 gpc105 (
      {stage0_11[15]},
      {stage1_11[13]}
   );
   gpc1_1 gpc106 (
      {stage0_11[16]},
      {stage1_11[14]}
   );
   gpc1_1 gpc107 (
      {stage0_11[17]},
      {stage1_11[15]}
   );
   gpc1_1 gpc108 (
      {stage0_11[18]},
      {stage1_11[16]}
   );
   gpc1_1 gpc109 (
      {stage0_11[19]},
      {stage1_11[17]}
   );
   gpc1_1 gpc110 (
      {stage0_11[20]},
      {stage1_11[18]}
   );
   gpc1_1 gpc111 (
      {stage0_11[21]},
      {stage1_11[19]}
   );
   gpc1_1 gpc112 (
      {stage0_11[22]},
      {stage1_11[20]}
   );
   gpc1_1 gpc113 (
      {stage0_11[23]},
      {stage1_11[21]}
   );
   gpc1_1 gpc114 (
      {stage0_11[24]},
      {stage1_11[22]}
   );
   gpc1_1 gpc115 (
      {stage0_11[25]},
      {stage1_11[23]}
   );
   gpc1_1 gpc116 (
      {stage0_11[26]},
      {stage1_11[24]}
   );
   gpc1_1 gpc117 (
      {stage0_11[27]},
      {stage1_11[25]}
   );
   gpc1_1 gpc118 (
      {stage0_11[28]},
      {stage1_11[26]}
   );
   gpc1_1 gpc119 (
      {stage0_11[29]},
      {stage1_11[27]}
   );
   gpc1_1 gpc120 (
      {stage0_11[30]},
      {stage1_11[28]}
   );
   gpc1_1 gpc121 (
      {stage0_11[31]},
      {stage1_11[29]}
   );
   gpc606_5 gpc122 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc123 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc124 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc125 (
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc2135_5 gpc126 (
      {stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_5[12], stage1_5[13], stage1_5[14]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc127 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc615_5 gpc128 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc129 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[3]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[5],stage2_6[5]}
   );
   gpc615_5 gpc130 (
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[4]}
   );
   gpc615_5 gpc131 (
      {stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_9[1]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[5]}
   );
   gpc1163_5 gpc132 (
      {stage1_9[2], stage1_9[3], stage1_9[4]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_11[0]},
      {stage1_12[0]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[4],stage2_9[4]}
   );
   gpc615_5 gpc133 (
      {stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[18]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[5],stage2_9[5]}
   );
   gpc615_5 gpc134 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14]},
      {stage1_10[19]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc135 (
      {stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19]},
      {stage1_10[20]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[7],stage2_9[7]}
   );
   gpc615_5 gpc136 (
      {stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_10[21]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[8],stage2_9[8]}
   );
   gpc1_1 gpc137 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc138 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc139 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc140 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc141 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc142 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc143 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc144 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc145 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc146 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc147 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc148 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc149 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc150 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc151 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc152 (
      {stage1_3[10]},
      {stage2_3[4]}
   );
   gpc1_1 gpc153 (
      {stage1_3[11]},
      {stage2_3[5]}
   );
   gpc1_1 gpc154 (
      {stage1_4[13]},
      {stage2_4[6]}
   );
   gpc1_1 gpc155 (
      {stage1_7[4]},
      {stage2_7[6]}
   );
   gpc1_1 gpc156 (
      {stage1_7[5]},
      {stage2_7[7]}
   );
   gpc1_1 gpc157 (
      {stage1_7[6]},
      {stage2_7[8]}
   );
   gpc1_1 gpc158 (
      {stage1_7[7]},
      {stage2_7[9]}
   );
   gpc1_1 gpc159 (
      {stage1_7[8]},
      {stage2_7[10]}
   );
   gpc1_1 gpc160 (
      {stage1_7[9]},
      {stage2_7[11]}
   );
   gpc1_1 gpc161 (
      {stage1_7[10]},
      {stage2_7[12]}
   );
   gpc1_1 gpc162 (
      {stage1_9[25]},
      {stage2_9[9]}
   );
   gpc1_1 gpc163 (
      {stage1_9[26]},
      {stage2_9[10]}
   );
   gpc1_1 gpc164 (
      {stage1_9[27]},
      {stage2_9[11]}
   );
   gpc1_1 gpc165 (
      {stage1_9[28]},
      {stage2_9[12]}
   );
   gpc1_1 gpc166 (
      {stage1_10[22]},
      {stage2_10[9]}
   );
   gpc1_1 gpc167 (
      {stage1_10[23]},
      {stage2_10[10]}
   );
   gpc1_1 gpc168 (
      {stage1_10[24]},
      {stage2_10[11]}
   );
   gpc1_1 gpc169 (
      {stage1_11[25]},
      {stage2_11[7]}
   );
   gpc1_1 gpc170 (
      {stage1_11[26]},
      {stage2_11[8]}
   );
   gpc1_1 gpc171 (
      {stage1_11[27]},
      {stage2_11[9]}
   );
   gpc1_1 gpc172 (
      {stage1_11[28]},
      {stage2_11[10]}
   );
   gpc1_1 gpc173 (
      {stage1_11[29]},
      {stage2_11[11]}
   );
   gpc1_1 gpc174 (
      {stage1_12[1]},
      {stage2_12[7]}
   );
   gpc1_1 gpc175 (
      {stage1_12[2]},
      {stage2_12[8]}
   );
   gpc1_1 gpc176 (
      {stage1_13[0]},
      {stage2_13[5]}
   );
   gpc606_5 gpc177 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc178 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1]}
   );
   gpc606_5 gpc179 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[1]}
   );
   gpc615_5 gpc180 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc181 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[2],stage3_10[2],stage3_9[2]}
   );
   gpc606_5 gpc182 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[2],stage3_11[3],stage3_10[3]}
   );
   gpc615_5 gpc183 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[3],stage3_11[4]}
   );
   gpc1_1 gpc184 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc185 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc186 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc187 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc188 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc189 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc190 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc191 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc192 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc193 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc194 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc195 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc196 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc197 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
   gpc1_1 gpc198 (
      {stage2_2[1]},
      {stage3_2[2]}
   );
   gpc1_1 gpc199 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc200 (
      {stage2_5[0]},
      {stage3_5[2]}
   );
   gpc1_1 gpc201 (
      {stage2_5[1]},
      {stage3_5[3]}
   );
   gpc1_1 gpc202 (
      {stage2_5[2]},
      {stage3_5[4]}
   );
   gpc1_1 gpc203 (
      {stage2_5[3]},
      {stage3_5[5]}
   );
   gpc1_1 gpc204 (
      {stage2_7[6]},
      {stage3_7[2]}
   );
   gpc1_1 gpc205 (
      {stage2_7[7]},
      {stage3_7[3]}
   );
   gpc1_1 gpc206 (
      {stage2_7[8]},
      {stage3_7[4]}
   );
   gpc1_1 gpc207 (
      {stage2_7[9]},
      {stage3_7[5]}
   );
   gpc1_1 gpc208 (
      {stage2_7[10]},
      {stage3_7[6]}
   );
   gpc1_1 gpc209 (
      {stage2_7[11]},
      {stage3_7[7]}
   );
   gpc1_1 gpc210 (
      {stage2_7[12]},
      {stage3_7[8]}
   );
   gpc1_1 gpc211 (
      {stage2_8[5]},
      {stage3_8[3]}
   );
   gpc1_1 gpc212 (
      {stage2_11[11]},
      {stage3_11[5]}
   );
   gpc1_1 gpc213 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc214 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc207_4 gpc215 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5], stage3_0[6]},
      {stage3_2[0], stage3_2[1]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc2116_5 gpc216 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[2]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1]},
      {stage4_5[0],stage4_4[0],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc217 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1]}
   );
   gpc1343_5 gpc218 (
      {stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc219 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc220 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], 1'b0},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc221 (
      {stage3_0[7]},
      {stage4_0[1]}
   );
   gpc1_1 gpc222 (
      {stage3_4[2]},
      {stage4_4[1]}
   );
   gpc1_1 gpc223 (
      {stage3_6[0]},
      {stage4_6[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor_CLA32_12 compressor_CLA32_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h81b3a9b42d0ec2a32c11d4bdf239c37ea545081eecd06ee31be104e38bc7b133def3f1a801c993889fd48a9fedd1ad38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h84fb7507cd374fd3d89d9bf93ecfe69e60d50815ef5ea6b45f129588d9eb29426e8bed7fa0abb397422eb6aa0fac3ee0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h801140d3bd419adbd8100936192210f7e3906fdfe987997e13afa5b0ba9c933fcceb1fa4fd98276418b835434cce44a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3563b2615f6a03c931d5fe5084351a74fa2f5fd8f6665055facb784d3413f0de109c2efc8c39facbb531823362a94bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hdc479de0770079de38e2bf093b47432c8f99e0ec9e7be7cb2f33cf824591177ba80c0a766c13fb5967bd762a9422ee1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h27bdd755a2eebb059615dcd56ad6945e166288e59e96a5bcfc6042effee1771b5aed18fc4df8f48e07559351f13a6bb6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h797de45e7130bb51e9b924221c8b463d7eebd5be1d0f1749cc5af5ebf89c4ef5ab3e2f0d6c5ce8c6735c359ef332541f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h355280bf4adc32fe5800a2a3cc83cd6f7b5e25053a4f841860db9544a4115d6b6f040cc7a15db24389d55410b605628;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h67afbe6d36e354b4c20caf5aa9935aac82010259d7df1c78d5b46836011a79bac63543845178f4573d751fb0267b56a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'heb29556e65929aa98a8d75cdd55cc38cb820174806d796dc45c7ee887f29096d0ed9e0c78ad3c807e9fd257523a9c010;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbacc6e387cb2a00b6dfa0bdac23922353aad6d45d7df3bf1bbf573e4be84e8862935c740fa0d4f99545de41fe85772e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hec67210434ab91c14a161a6ef7a921fd66a09637417ee5f3727b52466c08d811a807779d9bfaab5d57456314f4d3c3c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h64193b6966b37ff7ed9ab3065b94317e03f99cc532d7f291a9efb0b3eec4bb961e4721bff209e77ab99a37ae7a8ce59c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h65a8c2caef0c4e9109531937ee2ba63664107f5e7ba65abe3f0d481c5823e47634e62aa4397ae5e350018cace7f1f437;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1a12407728eade3c9623d621634e35c8bf717b5bbf7f65355c058a87c346dc09ca782331e54b6d5c552a085f060013c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd9526b7253368b68d96c870fe77bba4acea63b667f07d1f049ceec65c706dcb75cca037f6b79827cd32de0fe90296d56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd85561738d87cd7270a220e59ad6159f4668c37b8014064f625151558611983c547a06934c845ff7051844ca07b266d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h26a27c0bb24588b74bacb5d63ced3e52c1f943f5c36a58576619c22ab7f4a4acca8552a0bd076dee9c1706a69a258a05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h12565ac2a3b82b4c5812b3b53209f73f4d3c5406e9ca04cebd63a4787a2b942a70d56fb612cb88ce8c52be8c33878ab4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb6f58e3e60a937dd1d28933decea9c43e2d84782f0d0fa0e832bd0fbbfa60d3b808f70d242b4da133b0c32da0d9aae70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h47dd4fa57adee21d748088a9441ba510e737ef505bf5086f28a41325ab273f6c138d47e2b5306033452eda68ab0a5796;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h54528cf5b69c3ca4de1900ad45bc8dff3e1e8184d55900793114dd4c1a04bd80b619db912d7c07967ca3e3f2c3a868c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4112a8ded8181d1aa9510daeb35abe846a58816ec6722e3d7b1164bbe31efa8b2495e5835da213cacb862f2db76065df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h482c556fac26108bdfe4a9ca16d5cb1f5368ee8dea7e69b7a3ee106cf83bfe49284b9be3b042fb76ec42ee905355bd15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h437db93b635005f7947c42111381582418a7ea5cb8686e8f0fdf262e0dd254bcafcb6a0f576583170f405c0bf2b1cade;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h848bf6feed51a80d847b48e36459c22ec044a62b2cdb658b150f02405424755a0de921313130ca595fc845ea991de93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf7d308421212164983d3060592a6266e9947f93b71c9108026880cc756c67aab3887aa393cc60f90f45878b30ff1cc94;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7072f744c23295c5c496d35d6f98923e3b1a465ff450678ab10b4a87f5712f83ef7634f1d629f5c84992ea07250d973f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hddd2eb7a04b5d7d8a98dc77b11daa79280f8f3b88ad0418fa2a3011a082fd6ee9b4ebcbfed3d9d5f9449e631cbd61ebe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h83d218b0275f47f08a9849a955f78be8d7b92aca0676efb98804efba1deec55a11a5e59ac4e512f8559e52828ae57f95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hed573248e71a2140876c9e81b2e0ac887a2c7487739745cb08ec561a7df2b610ef8b1ccf7d3583a30fb886436e324a8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h71fea28f60401b96e06f89900ceb158ac2fd4023aa3440bd8f84d70d95890ec71dc0e9da648d4940aa67f78b44075763;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h2f6659c44e25d0c3c0adac6726b4e82f73280d70251bcbf75986518e44464bf290d8e5076634b23ab4cb3cf42fa1b6de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3b3e0d091c63af3de10ed9465ae85b38dcaa30c56d19d99d3a83d3d9c74e4250b78e9dc0628ffa859e51722d7176037a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4e57ec18e578a99fd2b273184c1420b664d4a27c7c0b1d0de70f3de27f3d90f0dd4200f9ac17fab41c08a8e2eae47ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6d019f9b748c3045856590bfb0a05dfe3f7c50b8525bf420d6d5e720ef8aa1175aa093403b11bc6bdf454bd85045a0b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h959e0f712f106600108af45d7e900869f05bd87efc8de26a762bdce2feb12123d0a45e509cf09ee5255fff64c444d7e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4a8fa55f607b85237eaa30f5532287ac4a2f8ebfc3a1ccef6a091b4042f5248c18003574d1ac72ea777454d81fc82c5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'haf461fa7670fcc5277f6782b662804f35435cf84f5c295c0fe240e2ec8d592d5b59ef932c54fb0205d01471e7e38b070;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc46d142c0e6543f291467841e7375b39dfc6dea03c7b61270fef04a6390e6a3e74cc95dfdd20016e1f46c5aae6db5568;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h120311a51be11e60feedf6ffc139b22ed1a9bee7a38a69ba440767f33b753a74b76be8ec61c4df5f42f6d19aeb5f1acd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'heebd6817abc703082ad11ca2588e9d3ac6cc4d00b21de1281ddf69f0207c314a91ef9afc4363cfef35e2db3281210520;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha2ba73610653fb65ecf5ec4c06011bae099aa648adb87d78384990c6cfe7bd762c7decc579fe808811a5caf66a3f8b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h66d25dbb194926037c31a37ca52f346c527c1fc5bbed0e6fda542650eae69dc2f82b3926e659c9ec46ace061c65c4bcb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd9eff6a83c7c04270de30043fc7f7a771cb2cdf7ad82ff3d55d5ad4476b25c54336c9475d2628023c7572ab008f668aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1804d720f1357a28f91c2238eeb29f292fce464a78c92177ec0ac8f045b458c385381ac606ca75220f3211f099c24651;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3b3fd066241060506b8b98fc6f02a191506a0cae21b348a21eb42cfbb7b05a2141d45c908c70ec8e517e1244fd36e843;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h964e9d5277c6bf3259de48bf277176dea4ff379890e6d86cb9955bcebea790bc5b7db9473fefccc799bb240c88cac790;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hba3d3c3a814f558d951c3c0b3a37c7104f9b94401d05a874f7058a43465f67b4de34b321783eae4de82ced7bfbacc808;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hbd02c3ee8b6b96e8130cd5e4858ee06cc2f925d02ef6df951d67abc42a5b1334e972279df31c1f68f3643cf5cd6ec27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h220c7d4f62628e14fd00b9288af5db9e4bd0d65587791a76b75c3d32e2d6ccfa8e98cc0c8f2b4b96e1cd801facc3590e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1241f5f6ec93077530e79f7f85873d484f3c172fadc43264edbb5b92ebcc96f01122407852cb9796a1501bc060190dea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he8edcfaafff26fdc2a8315aad9839c6b9216c5eca305e5a89416512c01ea8f3fe96b1a3f71bba10ff6055fc6a733c2e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8119242eec355b5909526d572495d0a24c8538a8af52b4065aefee35f8e6d81454037cb77801ece6544bf894e35f777c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hadda99491a3311b61e3e9b04c29d2304c71c4fbc9e5617a99a5dcb9e1f02a3fb2d25a597029a37c4332562f3c488ca2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he03fd8be8921cb12a1f6f848e2f61d131d597c660efef657698566b9a5fec49e0e103f0abc9a9a5383f2fd888cedde2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8f09f2ceb0cc490001920e1c7423590d1ed51b5ead8bc0d07099f56b25509c090c761f233cb7cbb8a76e471d6653240f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hb0606258fd06aa5ca8e13627afe9d6edf8fdc76c844c3b4ed4bc6d5ed974ad68bbd8b18a9e787d376a90cab3ef6aa367;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h9917fd643a1510188f5e8c383fe6ccf4bedf491b4501f27ca631cfa025d0cd335585c42bd887bdc67721c5d9fe610965;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h7ee55f6f599c5cbff457568303fc39236272f15c851d723416266cef6b14a7a0b7d10e2eb0e20f9c51924279bffc4077;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3e4e56d1fe276eec258dced27a92b273014c2b377b7f36d6ffdb2d8a04e74820928167a5fe184e4474c3f3895dd1f5f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h83e1307c0a219b7817ebb019c7f03c60d9298950e53816bd453f91758b9e74695b210b69fcd63407d23e35a25f1cb691;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4564edb9512a24cab091dfe99fea746f56e9601eec35f79cad3bd176280dc6d1af2ffe98c654c122dd4a4dce4829b86e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he7bcf055561cb5902275ca3f0ab67748ca43f0b3251a4ba325711dbc49b95ea86b3ee5037d7a6902dc15567af5a03a38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hed9432050cb586e53833da8e03059f966e9754af194b09502c0fd861742b4b38d19f619e25c207c61a377431b2cff96f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h9528f2f5ac699e5d9a3c192acd0cc70e9c198c1e6a5fa1592ec6c62e3cf6087dc0e4dcd569d38773b7c29507fdf61c7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc68dcb4a0c2a7f7b7369696d72b50ef503ea42e4674a2c1f1a3e357725a039c725b83d208763a3f8c7e44745b7c85275;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h8934e1f17143b0cfb8e53ead27d6325f92405077816229bde84e6dc79824ff2644cf964adc7703633989369328dd2fb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4d8aa3fc8716b703e8559957e235325ba70689fe3968654cf7e41a993fabfce16da29cdf59dea83851080f830cab9c6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h392acec8b0d449e314cba1d9fef832207e742abfa70ba17c4fac381306e54e2efca431c9ad889857bf4f70ee7d70b30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hc78ff0e8c319f692a589438b513641e28309ec0cc5f137208858f9b30b83e16de484cf6f3308079129217f217741ca75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h453eafcfe89b2b6abe8cd656e26a07a395aecf32175ba280b4f3c5749eedc9253385cdf20f1cf9c23e5a8deed008c6a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hcda61046c5615d686ae41fff1e5a39d2432257dcb70202bb4155df8d1f9feefcc4c49ce6323356d86570f16ba582aed9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hfccbaff2f266784c56678bbf1a66c9d3c4bde1c733f19c4265baedd61ec788397d62099786393033ee5f9201248cdef1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'haa9e66513d22f0bb10f96279c3d969f65518d704a62ae13c9b71ab04f7928e88af6ecf2f5608be62b19d0d088aafd1ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h81db0fb5a6ff005a4b5e80bdca4adbc805c08de16a3a9c576d1266116d56bced8317a2914031740f52a9d755be5b7799;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hd01e205286ef3b56694420ebe72faefc47652bae15fe47d5b770b6ce482ec9df4e678d7b611e30ff628534087e53353d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hcc79a4441a6c2084f79f746d9cf4ce8338435527e66702cfa7280948b7207c8238fda6769dcc8142dff925e0d426b100;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h861d63bcb400329568f59917605e561e76a3139654f333019a7f9b32b2760af9ed6873b7ec3fb286df80618a6da16b80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1c355ab41d27548db5c510de2cb69e57369bccfd7e081d5a95f0b040de84797e884c39b707d7569ccf8819b78ca0156;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3c0da1c76c216294848672693d1a6cf9e3b8f8a77976aa57b254ed77c4addf647b0c8e8989c4a1e7bfe7688ba1828c02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h63890221a7b64526b67edf0f145f51749e2acf7be24c257c1a0d96a6a46c38113ef03f51bd412a8423cfe60bac444238;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'he69976df31f960c98330f8c3d0a71e4cbd29d48c7375df09304cb938ef9b8eb54d05ef69270c4b728924cb240f18c2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h822e1b857f1d78f59380a12be62bcad9dfabc9fa44309593759093ecc46e19484a9f175089c79868b0062e58c2b83419;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3d9412945a94752388b9432ac599a30cc0ddc1783043bf475e3a5dc40bbca8190c77abec1e13a2ddf2c35ba6b49cc05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha5118f7e29509ee2b7f502df00ef8b86528a168daf5b722635143b2c58b04a710dd7982eb44aa0edd0cbb261b3ac409c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h6582d56fbbb50eb8e1d43188e9513912f642a53c5ff2376ae142dea10b42bc81a83e846d6c8094b99d3ef8a85d8fdd58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3fb9eeb9102049a9e64b1643f09f388657e0b9f5933fb41104db25ac2464e07389ebb6e79143bb5a9588a7d4358d4f74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h4e2526e79cef07bbb9e234734401e1dc174842041138a3bfb459bf9daab39790ebfebc506e9a9df1d2dad55771b32a3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h87bb59acf0d1aeb9a58cbddc0ef2234243133927a3331af002ef0ee8f2740b45881e9e483657cb2f577f671e778c1ab1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h3799e0027066f3298fab089ce03caefbb62c978fddcef5b0316cff4ac6c1ada6339a4549c2cfabdd3821bc416e95f70c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h1b4ff1d091d8572e1a66ff491974ba985811008c9f1491466709e42ee9f35b95e9f267dd9cde5c7ebbed286184123791;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h5579fa38afbfe6fbec51a503d03342f26105108f44cc3c1b255912062feaf8f0dec98fbe2c8e7eb509dfb3ec4b825dc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h817c443afea71ede6d6b29cf82170703d291477096fbbd51e71352fafb3920bfe39850edd31b6c2992945b435e67c18e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h98f57459c7e931af108433422d8cc694ff6de89eaf666e7e640dc05f4dc096d405e0ab3ab0127e1f0809112b9f50d002;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hde4d00cacb473a7ad657b361b79251f604b0b98ab831970b6c9a7028a06fea8d4b53249017827e21cede69c3fd2509cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hdeee6f82535798a48754b4faf34b0a0e5acf35096909488dc22834d23dd8518d2080f884737a6ba95748d17e15f914bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'hf2134da512fb81cc29a00e3c0d8b9c3a32499ff3d7e9fdb011b71a7ba4370f95486c824c45e3889af8c6900beba0f806;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'h2170dcd8b2f36f38dd33aa0e19f5f153646f9bc15a4b714b15d2133d8d187737c32085c360591cd54265b7dc22600e8c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 384'ha03d011de104cad37b95eb66369f5624ac904cf8710b4e566d7dc2a857fa040a995cc023dcd5e79a1160ebee1c876dbe;
        #1
        $finish();
    end
endmodule
