module compressor_without_rowadder (
      input wire [0:0] src0,
      input wire [1:0] src1,
      input wire [2:0] src2,
      input wire [3:0] src3,
      input wire [4:0] src4,
      input wire [5:0] src5,
      input wire [6:0] src6,
      input wire [7:0] src7,
      input wire [8:0] src8,
      input wire [9:0] src9,
      input wire [10:0] src10,
      input wire [11:0] src11,
      input wire [12:0] src12,
      input wire [13:0] src13,
      input wire [14:0] src14,
      input wire [15:0] src15,
      input wire [16:0] src16,
      input wire [17:0] src17,
      input wire [18:0] src18,
      input wire [19:0] src19,
      input wire [20:0] src20,
      input wire [21:0] src21,
      input wire [22:0] src22,
      input wire [23:0] src23,
      input wire [24:0] src24,
      input wire [25:0] src25,
      input wire [26:0] src26,
      input wire [27:0] src27,
      input wire [28:0] src28,
      input wire [29:0] src29,
      input wire [28:0] src30,
      input wire [27:0] src31,
      input wire [26:0] src32,
      input wire [25:0] src33,
      input wire [24:0] src34,
      input wire [23:0] src35,
      input wire [22:0] src36,
      input wire [21:0] src37,
      input wire [20:0] src38,
      input wire [19:0] src39,
      input wire [18:0] src40,
      input wire [17:0] src41,
      input wire [16:0] src42,
      input wire [15:0] src43,
      input wire [14:0] src44,
      input wire [13:0] src45,
      input wire [12:0] src46,
      input wire [11:0] src47,
      input wire [10:0] src48,
      input wire [9:0] src49,
      input wire [8:0] src50,
      input wire [7:0] src51,
      input wire [6:0] src52,
      input wire [5:0] src53,
      input wire [4:0] src54,
      input wire [3:0] src55,
      input wire [2:0] src56,
      input wire [1:0] src57,
      input wire [0:0] src58,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [0:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [0:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [0:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [0:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [0:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [0:0] dst58,
      output wire [0:0] dst59);

   wire [0:0] stage0_0;
   wire [1:0] stage0_1;
   wire [2:0] stage0_2;
   wire [3:0] stage0_3;
   wire [4:0] stage0_4;
   wire [5:0] stage0_5;
   wire [6:0] stage0_6;
   wire [7:0] stage0_7;
   wire [8:0] stage0_8;
   wire [9:0] stage0_9;
   wire [10:0] stage0_10;
   wire [11:0] stage0_11;
   wire [12:0] stage0_12;
   wire [13:0] stage0_13;
   wire [14:0] stage0_14;
   wire [15:0] stage0_15;
   wire [16:0] stage0_16;
   wire [17:0] stage0_17;
   wire [18:0] stage0_18;
   wire [19:0] stage0_19;
   wire [20:0] stage0_20;
   wire [21:0] stage0_21;
   wire [22:0] stage0_22;
   wire [23:0] stage0_23;
   wire [24:0] stage0_24;
   wire [25:0] stage0_25;
   wire [26:0] stage0_26;
   wire [27:0] stage0_27;
   wire [28:0] stage0_28;
   wire [29:0] stage0_29;
   wire [28:0] stage0_30;
   wire [27:0] stage0_31;
   wire [26:0] stage0_32;
   wire [25:0] stage0_33;
   wire [24:0] stage0_34;
   wire [23:0] stage0_35;
   wire [22:0] stage0_36;
   wire [21:0] stage0_37;
   wire [20:0] stage0_38;
   wire [19:0] stage0_39;
   wire [18:0] stage0_40;
   wire [17:0] stage0_41;
   wire [16:0] stage0_42;
   wire [15:0] stage0_43;
   wire [14:0] stage0_44;
   wire [13:0] stage0_45;
   wire [12:0] stage0_46;
   wire [11:0] stage0_47;
   wire [10:0] stage0_48;
   wire [9:0] stage0_49;
   wire [8:0] stage0_50;
   wire [7:0] stage0_51;
   wire [6:0] stage0_52;
   wire [5:0] stage0_53;
   wire [4:0] stage0_54;
   wire [3:0] stage0_55;
   wire [2:0] stage0_56;
   wire [1:0] stage0_57;
   wire [0:0] stage0_58;
   wire [0:0] stage1_0;
   wire [1:0] stage1_1;
   wire [2:0] stage1_2;
   wire [3:0] stage1_3;
   wire [4:0] stage1_4;
   wire [0:0] stage1_5;
   wire [7:0] stage1_6;
   wire [2:0] stage1_7;
   wire [9:0] stage1_8;
   wire [6:0] stage1_9;
   wire [9:0] stage1_10;
   wire [4:0] stage1_11;
   wire [5:0] stage1_12;
   wire [5:0] stage1_13;
   wire [5:0] stage1_14;
   wire [5:0] stage1_15;
   wire [8:0] stage1_16;
   wire [8:0] stage1_17;
   wire [5:0] stage1_18;
   wire [20:0] stage1_19;
   wire [13:0] stage1_20;
   wire [5:0] stage1_21;
   wire [9:0] stage1_22;
   wire [7:0] stage1_23;
   wire [17:0] stage1_24;
   wire [19:0] stage1_25;
   wire [11:0] stage1_26;
   wire [17:0] stage1_27;
   wire [11:0] stage1_28;
   wire [12:0] stage1_29;
   wire [12:0] stage1_30;
   wire [13:0] stage1_31;
   wire [12:0] stage1_32;
   wire [21:0] stage1_33;
   wire [14:0] stage1_34;
   wire [17:0] stage1_35;
   wire [7:0] stage1_36;
   wire [19:0] stage1_37;
   wire [9:0] stage1_38;
   wire [18:0] stage1_39;
   wire [11:0] stage1_40;
   wire [7:0] stage1_41;
   wire [5:0] stage1_42;
   wire [13:0] stage1_43;
   wire [7:0] stage1_44;
   wire [5:0] stage1_45;
   wire [16:0] stage1_46;
   wire [7:0] stage1_47;
   wire [11:0] stage1_48;
   wire [6:0] stage1_49;
   wire [8:0] stage1_50;
   wire [2:0] stage1_51;
   wire [7:0] stage1_52;
   wire [6:0] stage1_53;
   wire [4:0] stage1_54;
   wire [3:0] stage1_55;
   wire [2:0] stage1_56;
   wire [1:0] stage1_57;
   wire [0:0] stage1_58;
   wire [0:0] stage2_0;
   wire [1:0] stage2_1;
   wire [0:0] stage2_2;
   wire [1:0] stage2_3;
   wire [1:0] stage2_4;
   wire [1:0] stage2_5;
   wire [5:0] stage2_6;
   wire [0:0] stage2_7;
   wire [7:0] stage2_8;
   wire [6:0] stage2_9;
   wire [5:0] stage2_10;
   wire [5:0] stage2_11;
   wire [0:0] stage2_12;
   wire [1:0] stage2_13;
   wire [2:0] stage2_14;
   wire [1:0] stage2_15;
   wire [4:0] stage2_16;
   wire [3:0] stage2_17;
   wire [6:0] stage2_18;
   wire [6:0] stage2_19;
   wire [15:0] stage2_20;
   wire [2:0] stage2_21;
   wire [5:0] stage2_22;
   wire [5:0] stage2_23;
   wire [4:0] stage2_24;
   wire [5:0] stage2_25;
   wire [5:0] stage2_26;
   wire [5:0] stage2_27;
   wire [8:0] stage2_28;
   wire [5:0] stage2_29;
   wire [3:0] stage2_30;
   wire [11:0] stage2_31;
   wire [5:0] stage2_32;
   wire [12:0] stage2_33;
   wire [4:0] stage2_34;
   wire [4:0] stage2_35;
   wire [9:0] stage2_36;
   wire [6:0] stage2_37;
   wire [4:0] stage2_38;
   wire [4:0] stage2_39;
   wire [6:0] stage2_40;
   wire [6:0] stage2_41;
   wire [2:0] stage2_42;
   wire [9:0] stage2_43;
   wire [5:0] stage2_44;
   wire [6:0] stage2_45;
   wire [7:0] stage2_46;
   wire [5:0] stage2_47;
   wire [8:0] stage2_48;
   wire [2:0] stage2_49;
   wire [5:0] stage2_50;
   wire [4:0] stage2_51;
   wire [2:0] stage2_52;
   wire [5:0] stage2_53;
   wire [4:0] stage2_54;
   wire [0:0] stage2_55;
   wire [2:0] stage2_56;
   wire [2:0] stage2_57;
   wire [0:0] stage2_58;
   wire [0:0] stage3_0;
   wire [1:0] stage3_1;
   wire [0:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [0:0] stage3_7;
   wire [1:0] stage3_8;
   wire [6:0] stage3_9;
   wire [1:0] stage3_10;
   wire [6:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [2:0] stage3_14;
   wire [1:0] stage3_15;
   wire [4:0] stage3_16;
   wire [0:0] stage3_17;
   wire [4:0] stage3_18;
   wire [1:0] stage3_19;
   wire [6:0] stage3_20;
   wire [5:0] stage3_21;
   wire [1:0] stage3_22;
   wire [6:0] stage3_23;
   wire [3:0] stage3_24;
   wire [0:0] stage3_25;
   wire [1:0] stage3_26;
   wire [2:0] stage3_27;
   wire [2:0] stage3_28;
   wire [2:0] stage3_29;
   wire [6:0] stage3_30;
   wire [2:0] stage3_31;
   wire [4:0] stage3_32;
   wire [3:0] stage3_33;
   wire [2:0] stage3_34;
   wire [5:0] stage3_35;
   wire [1:0] stage3_36;
   wire [4:0] stage3_37;
   wire [2:0] stage3_38;
   wire [1:0] stage3_39;
   wire [2:0] stage3_40;
   wire [4:0] stage3_41;
   wire [1:0] stage3_42;
   wire [5:0] stage3_43;
   wire [2:0] stage3_44;
   wire [2:0] stage3_45;
   wire [3:0] stage3_46;
   wire [1:0] stage3_47;
   wire [5:0] stage3_48;
   wire [4:0] stage3_49;
   wire [0:0] stage3_50;
   wire [1:0] stage3_51;
   wire [4:0] stage3_52;
   wire [0:0] stage3_53;
   wire [5:0] stage3_54;
   wire [1:0] stage3_55;
   wire [2:0] stage3_56;
   wire [2:0] stage3_57;
   wire [0:0] stage3_58;
   wire [0:0] stage4_0;
   wire [1:0] stage4_1;
   wire [0:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [0:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [0:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [0:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [0:0] stage4_26;
   wire [1:0] stage4_27;
   wire [1:0] stage4_28;
   wire [1:0] stage4_29;
   wire [1:0] stage4_30;
   wire [1:0] stage4_31;
   wire [1:0] stage4_32;
   wire [1:0] stage4_33;
   wire [1:0] stage4_34;
   wire [1:0] stage4_35;
   wire [1:0] stage4_36;
   wire [1:0] stage4_37;
   wire [1:0] stage4_38;
   wire [1:0] stage4_39;
   wire [1:0] stage4_40;
   wire [1:0] stage4_41;
   wire [1:0] stage4_42;
   wire [0:0] stage4_43;
   wire [1:0] stage4_44;
   wire [1:0] stage4_45;
   wire [1:0] stage4_46;
   wire [1:0] stage4_47;
   wire [1:0] stage4_48;
   wire [1:0] stage4_49;
   wire [1:0] stage4_50;
   wire [1:0] stage4_51;
   wire [1:0] stage4_52;
   wire [1:0] stage4_53;
   wire [0:0] stage4_54;
   wire [1:0] stage4_55;
   wire [1:0] stage4_56;
   wire [1:0] stage4_57;
   wire [0:0] stage4_58;
   wire [0:0] stage4_59;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;
   assign dst31 = stage4_31;
   assign dst32 = stage4_32;
   assign dst33 = stage4_33;
   assign dst34 = stage4_34;
   assign dst35 = stage4_35;
   assign dst36 = stage4_36;
   assign dst37 = stage4_37;
   assign dst38 = stage4_38;
   assign dst39 = stage4_39;
   assign dst40 = stage4_40;
   assign dst41 = stage4_41;
   assign dst42 = stage4_42;
   assign dst43 = stage4_43;
   assign dst44 = stage4_44;
   assign dst45 = stage4_45;
   assign dst46 = stage4_46;
   assign dst47 = stage4_47;
   assign dst48 = stage4_48;
   assign dst49 = stage4_49;
   assign dst50 = stage4_50;
   assign dst51 = stage4_51;
   assign dst52 = stage4_52;
   assign dst53 = stage4_53;
   assign dst54 = stage4_54;
   assign dst55 = stage4_55;
   assign dst56 = stage4_56;
   assign dst57 = stage4_57;
   assign dst58 = stage4_58;
   assign dst59 = stage4_59;

   gpc606_5 gpc0 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[0],stage1_7[0],stage1_6[0],stage1_5[0]}
   );
   gpc425_5 gpc1 (
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4]},
      {stage0_10[0], stage0_10[1]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3]},
      {stage1_13[0],stage1_12[0],stage1_11[0],stage1_10[0],stage1_9[1]}
   );
   gpc615_5 gpc2 (
      {stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8]},
      {stage0_12[0]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[1],stage1_12[1],stage1_11[1]}
   );
   gpc615_5 gpc3 (
      {stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage0_13[6]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[2],stage1_12[2]}
   );
   gpc615_5 gpc4 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10]},
      {stage0_13[7]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[3],stage1_12[3]}
   );
   gpc1415_5 gpc5 (
      {stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12]},
      {stage0_14[12]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3]},
      {stage0_16[0]},
      {stage1_17[0],stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[4]}
   );
   gpc606_5 gpc6 (
      {stage0_15[4], stage0_15[5], stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[0],stage1_17[1],stage1_16[3],stage1_15[4]}
   );
   gpc606_5 gpc7 (
      {stage0_15[10], stage0_15[11], stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[1],stage1_17[2],stage1_16[4],stage1_15[5]}
   );
   gpc615_5 gpc8 (
      {stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage0_17[12]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[2],stage1_18[2],stage1_17[3],stage1_16[5]}
   );
   gpc615_5 gpc9 (
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10]},
      {stage0_17[13]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[3],stage1_18[3],stage1_17[4],stage1_16[6]}
   );
   gpc615_5 gpc10 (
      {stage0_16[11], stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15]},
      {stage0_17[14]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[4],stage1_18[4],stage1_17[5],stage1_16[7]}
   );
   gpc615_5 gpc11 (
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4]},
      {stage0_20[0]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[0],stage1_20[3],stage1_19[5]}
   );
   gpc606_5 gpc12 (
      {stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5], stage0_20[6]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[1],stage1_22[1],stage1_21[1],stage1_20[4]}
   );
   gpc606_5 gpc13 (
      {stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[2],stage1_22[2],stage1_21[2],stage1_20[5]}
   );
   gpc606_5 gpc14 (
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[2],stage1_23[3],stage1_22[3],stage1_21[3]}
   );
   gpc615_5 gpc15 (
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16]},
      {stage0_22[12]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[3],stage1_23[4],stage1_22[4],stage1_21[4]}
   );
   gpc615_5 gpc16 (
      {stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21]},
      {stage0_22[13]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[4],stage1_23[5],stage1_22[5],stage1_21[5]}
   );
   gpc606_5 gpc17 (
      {stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17], stage0_22[18], stage0_22[19]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[3],stage1_24[5],stage1_23[6],stage1_22[6]}
   );
   gpc606_5 gpc18 (
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[4],stage1_24[6],stage1_23[7]}
   );
   gpc615_5 gpc19 (
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10]},
      {stage0_25[6]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[2],stage1_25[5],stage1_24[7]}
   );
   gpc615_5 gpc20 (
      {stage0_24[11], stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15]},
      {stage0_25[7]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[2],stage1_26[3],stage1_25[6],stage1_24[8]}
   );
   gpc606_5 gpc21 (
      {stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11], stage0_25[12], stage0_25[13]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[2],stage1_27[3],stage1_26[4],stage1_25[7]}
   );
   gpc425_5 gpc22 (
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16]},
      {stage0_27[6], stage0_27[7]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3]},
      {stage1_30[0],stage1_29[1],stage1_28[3],stage1_27[4],stage1_26[5]}
   );
   gpc615_5 gpc23 (
      {stage0_26[17], stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21]},
      {stage0_27[8]},
      {stage0_28[4], stage0_28[5], stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9]},
      {stage1_30[1],stage1_29[2],stage1_28[4],stage1_27[5],stage1_26[6]}
   );
   gpc615_5 gpc24 (
      {stage0_27[9], stage0_27[10], stage0_27[11], stage0_27[12], stage0_27[13]},
      {stage0_28[10]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[2],stage1_29[3],stage1_28[5],stage1_27[6]}
   );
   gpc1334_5 gpc25 (
      {stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage0_28[11], stage0_28[12], stage0_28[13]},
      {stage0_29[6], stage0_29[7], stage0_29[8]},
      {stage0_30[0]},
      {stage1_31[1],stage1_30[3],stage1_29[4],stage1_28[6],stage1_27[7]}
   );
   gpc606_5 gpc26 (
      {stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19]},
      {stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6]},
      {stage1_32[0],stage1_31[2],stage1_30[4],stage1_29[5],stage1_28[7]}
   );
   gpc1316_5 gpc27 (
      {stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25]},
      {stage0_29[9]},
      {stage0_30[7], stage0_30[8], stage0_30[9]},
      {stage0_31[0]},
      {stage1_32[1],stage1_31[3],stage1_30[5],stage1_29[6],stage1_28[8]}
   );
   gpc606_5 gpc28 (
      {stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15]},
      {stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6]},
      {stage1_33[0],stage1_32[2],stage1_31[4],stage1_30[6],stage1_29[7]}
   );
   gpc606_5 gpc29 (
      {stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21]},
      {stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12]},
      {stage1_33[1],stage1_32[3],stage1_31[5],stage1_30[7],stage1_29[8]}
   );
   gpc615_5 gpc30 (
      {stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25], stage0_29[26]},
      {stage0_30[10]},
      {stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18]},
      {stage1_33[2],stage1_32[4],stage1_31[6],stage1_30[8],stage1_29[9]}
   );
   gpc606_5 gpc31 (
      {stage0_30[11], stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[3],stage1_32[5],stage1_31[7],stage1_30[9]}
   );
   gpc606_5 gpc32 (
      {stage0_30[17], stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[4],stage1_32[6],stage1_31[8],stage1_30[10]}
   );
   gpc615_5 gpc33 (
      {stage0_30[23], stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27]},
      {stage0_31[19]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[5],stage1_32[7],stage1_31[9],stage1_30[11]}
   );
   gpc615_5 gpc34 (
      {stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24]},
      {stage0_32[18]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[3],stage1_33[6],stage1_32[8],stage1_31[10]}
   );
   gpc615_5 gpc35 (
      {stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage0_33[6]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[1],stage1_34[4],stage1_33[7],stage1_32[9]}
   );
   gpc606_5 gpc36 (
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[1],stage1_35[2],stage1_34[5],stage1_33[8]}
   );
   gpc606_5 gpc37 (
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[1],stage1_36[2],stage1_35[3],stage1_34[6]}
   );
   gpc606_5 gpc38 (
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[2],stage1_36[3],stage1_35[4],stage1_34[7]}
   );
   gpc606_5 gpc39 (
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[2],stage1_37[3],stage1_36[4],stage1_35[5]}
   );
   gpc615_5 gpc40 (
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16]},
      {stage0_37[6]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[1],stage1_38[3],stage1_37[4],stage1_36[5]}
   );
   gpc615_5 gpc41 (
      {stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21]},
      {stage0_37[7]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[2],stage1_38[4],stage1_37[5],stage1_36[6]}
   );
   gpc615_5 gpc42 (
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16]},
      {stage0_39[0]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[0],stage1_40[2],stage1_39[3],stage1_38[5]}
   );
   gpc615_5 gpc43 (
      {stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage0_40[6]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[1],stage1_41[1],stage1_40[3],stage1_39[4]}
   );
   gpc1171_5 gpc44 (
      {stage0_40[7]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11], stage0_41[12]},
      {stage0_42[0]},
      {stage0_43[0]},
      {stage1_44[0],stage1_43[1],stage1_42[2],stage1_41[2],stage1_40[4]}
   );
   gpc1415_5 gpc45 (
      {stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11], stage0_40[12]},
      {stage0_41[13]},
      {stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4]},
      {stage0_43[1]},
      {stage1_44[1],stage1_43[2],stage1_42[3],stage1_41[3],stage1_40[5]}
   );
   gpc606_5 gpc46 (
      {stage0_42[5], stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[0],stage1_44[2],stage1_43[3],stage1_42[4]}
   );
   gpc606_5 gpc47 (
      {stage0_42[11], stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[1],stage1_44[3],stage1_43[4],stage1_42[5]}
   );
   gpc606_5 gpc48 (
      {stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6], stage0_43[7]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[2],stage1_45[2],stage1_44[4],stage1_43[5]}
   );
   gpc606_5 gpc49 (
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[0],stage1_47[1],stage1_46[3],stage1_45[3]}
   );
   gpc615_5 gpc50 (
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4]},
      {stage0_50[0]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[0],stage1_51[0],stage1_50[0],stage1_49[1]}
   );
   gpc1_1 gpc51 (
      {stage0_0[0]},
      {stage1_0[0]}
   );
   gpc1_1 gpc52 (
      {stage0_1[0]},
      {stage1_1[0]}
   );
   gpc1_1 gpc53 (
      {stage0_1[1]},
      {stage1_1[1]}
   );
   gpc1_1 gpc54 (
      {stage0_2[0]},
      {stage1_2[0]}
   );
   gpc1_1 gpc55 (
      {stage0_2[1]},
      {stage1_2[1]}
   );
   gpc1_1 gpc56 (
      {stage0_2[2]},
      {stage1_2[2]}
   );
   gpc1_1 gpc57 (
      {stage0_3[0]},
      {stage1_3[0]}
   );
   gpc1_1 gpc58 (
      {stage0_3[1]},
      {stage1_3[1]}
   );
   gpc1_1 gpc59 (
      {stage0_3[2]},
      {stage1_3[2]}
   );
   gpc1_1 gpc60 (
      {stage0_3[3]},
      {stage1_3[3]}
   );
   gpc1_1 gpc61 (
      {stage0_4[0]},
      {stage1_4[0]}
   );
   gpc1_1 gpc62 (
      {stage0_4[1]},
      {stage1_4[1]}
   );
   gpc1_1 gpc63 (
      {stage0_4[2]},
      {stage1_4[2]}
   );
   gpc1_1 gpc64 (
      {stage0_4[3]},
      {stage1_4[3]}
   );
   gpc1_1 gpc65 (
      {stage0_4[4]},
      {stage1_4[4]}
   );
   gpc1_1 gpc66 (
      {stage0_6[0]},
      {stage1_6[1]}
   );
   gpc1_1 gpc67 (
      {stage0_6[1]},
      {stage1_6[2]}
   );
   gpc1_1 gpc68 (
      {stage0_6[2]},
      {stage1_6[3]}
   );
   gpc1_1 gpc69 (
      {stage0_6[3]},
      {stage1_6[4]}
   );
   gpc1_1 gpc70 (
      {stage0_6[4]},
      {stage1_6[5]}
   );
   gpc1_1 gpc71 (
      {stage0_6[5]},
      {stage1_6[6]}
   );
   gpc1_1 gpc72 (
      {stage0_6[6]},
      {stage1_6[7]}
   );
   gpc1_1 gpc73 (
      {stage0_7[6]},
      {stage1_7[1]}
   );
   gpc1_1 gpc74 (
      {stage0_7[7]},
      {stage1_7[2]}
   );
   gpc1_1 gpc75 (
      {stage0_8[0]},
      {stage1_8[1]}
   );
   gpc1_1 gpc76 (
      {stage0_8[1]},
      {stage1_8[2]}
   );
   gpc1_1 gpc77 (
      {stage0_8[2]},
      {stage1_8[3]}
   );
   gpc1_1 gpc78 (
      {stage0_8[3]},
      {stage1_8[4]}
   );
   gpc1_1 gpc79 (
      {stage0_8[4]},
      {stage1_8[5]}
   );
   gpc1_1 gpc80 (
      {stage0_8[5]},
      {stage1_8[6]}
   );
   gpc1_1 gpc81 (
      {stage0_8[6]},
      {stage1_8[7]}
   );
   gpc1_1 gpc82 (
      {stage0_8[7]},
      {stage1_8[8]}
   );
   gpc1_1 gpc83 (
      {stage0_8[8]},
      {stage1_8[9]}
   );
   gpc1_1 gpc84 (
      {stage0_9[5]},
      {stage1_9[2]}
   );
   gpc1_1 gpc85 (
      {stage0_9[6]},
      {stage1_9[3]}
   );
   gpc1_1 gpc86 (
      {stage0_9[7]},
      {stage1_9[4]}
   );
   gpc1_1 gpc87 (
      {stage0_9[8]},
      {stage1_9[5]}
   );
   gpc1_1 gpc88 (
      {stage0_9[9]},
      {stage1_9[6]}
   );
   gpc1_1 gpc89 (
      {stage0_10[2]},
      {stage1_10[1]}
   );
   gpc1_1 gpc90 (
      {stage0_10[3]},
      {stage1_10[2]}
   );
   gpc1_1 gpc91 (
      {stage0_10[4]},
      {stage1_10[3]}
   );
   gpc1_1 gpc92 (
      {stage0_10[5]},
      {stage1_10[4]}
   );
   gpc1_1 gpc93 (
      {stage0_10[6]},
      {stage1_10[5]}
   );
   gpc1_1 gpc94 (
      {stage0_10[7]},
      {stage1_10[6]}
   );
   gpc1_1 gpc95 (
      {stage0_10[8]},
      {stage1_10[7]}
   );
   gpc1_1 gpc96 (
      {stage0_10[9]},
      {stage1_10[8]}
   );
   gpc1_1 gpc97 (
      {stage0_10[10]},
      {stage1_10[9]}
   );
   gpc1_1 gpc98 (
      {stage0_11[9]},
      {stage1_11[2]}
   );
   gpc1_1 gpc99 (
      {stage0_11[10]},
      {stage1_11[3]}
   );
   gpc1_1 gpc100 (
      {stage0_11[11]},
      {stage1_11[4]}
   );
   gpc1_1 gpc101 (
      {stage0_12[11]},
      {stage1_12[4]}
   );
   gpc1_1 gpc102 (
      {stage0_12[12]},
      {stage1_12[5]}
   );
   gpc1_1 gpc103 (
      {stage0_13[13]},
      {stage1_13[5]}
   );
   gpc1_1 gpc104 (
      {stage0_14[13]},
      {stage1_14[4]}
   );
   gpc1_1 gpc105 (
      {stage0_14[14]},
      {stage1_14[5]}
   );
   gpc1_1 gpc106 (
      {stage0_16[16]},
      {stage1_16[8]}
   );
   gpc1_1 gpc107 (
      {stage0_17[15]},
      {stage1_17[6]}
   );
   gpc1_1 gpc108 (
      {stage0_17[16]},
      {stage1_17[7]}
   );
   gpc1_1 gpc109 (
      {stage0_17[17]},
      {stage1_17[8]}
   );
   gpc1_1 gpc110 (
      {stage0_18[18]},
      {stage1_18[5]}
   );
   gpc1_1 gpc111 (
      {stage0_19[5]},
      {stage1_19[6]}
   );
   gpc1_1 gpc112 (
      {stage0_19[6]},
      {stage1_19[7]}
   );
   gpc1_1 gpc113 (
      {stage0_19[7]},
      {stage1_19[8]}
   );
   gpc1_1 gpc114 (
      {stage0_19[8]},
      {stage1_19[9]}
   );
   gpc1_1 gpc115 (
      {stage0_19[9]},
      {stage1_19[10]}
   );
   gpc1_1 gpc116 (
      {stage0_19[10]},
      {stage1_19[11]}
   );
   gpc1_1 gpc117 (
      {stage0_19[11]},
      {stage1_19[12]}
   );
   gpc1_1 gpc118 (
      {stage0_19[12]},
      {stage1_19[13]}
   );
   gpc1_1 gpc119 (
      {stage0_19[13]},
      {stage1_19[14]}
   );
   gpc1_1 gpc120 (
      {stage0_19[14]},
      {stage1_19[15]}
   );
   gpc1_1 gpc121 (
      {stage0_19[15]},
      {stage1_19[16]}
   );
   gpc1_1 gpc122 (
      {stage0_19[16]},
      {stage1_19[17]}
   );
   gpc1_1 gpc123 (
      {stage0_19[17]},
      {stage1_19[18]}
   );
   gpc1_1 gpc124 (
      {stage0_19[18]},
      {stage1_19[19]}
   );
   gpc1_1 gpc125 (
      {stage0_19[19]},
      {stage1_19[20]}
   );
   gpc1_1 gpc126 (
      {stage0_20[13]},
      {stage1_20[6]}
   );
   gpc1_1 gpc127 (
      {stage0_20[14]},
      {stage1_20[7]}
   );
   gpc1_1 gpc128 (
      {stage0_20[15]},
      {stage1_20[8]}
   );
   gpc1_1 gpc129 (
      {stage0_20[16]},
      {stage1_20[9]}
   );
   gpc1_1 gpc130 (
      {stage0_20[17]},
      {stage1_20[10]}
   );
   gpc1_1 gpc131 (
      {stage0_20[18]},
      {stage1_20[11]}
   );
   gpc1_1 gpc132 (
      {stage0_20[19]},
      {stage1_20[12]}
   );
   gpc1_1 gpc133 (
      {stage0_20[20]},
      {stage1_20[13]}
   );
   gpc1_1 gpc134 (
      {stage0_22[20]},
      {stage1_22[7]}
   );
   gpc1_1 gpc135 (
      {stage0_22[21]},
      {stage1_22[8]}
   );
   gpc1_1 gpc136 (
      {stage0_22[22]},
      {stage1_22[9]}
   );
   gpc1_1 gpc137 (
      {stage0_24[16]},
      {stage1_24[9]}
   );
   gpc1_1 gpc138 (
      {stage0_24[17]},
      {stage1_24[10]}
   );
   gpc1_1 gpc139 (
      {stage0_24[18]},
      {stage1_24[11]}
   );
   gpc1_1 gpc140 (
      {stage0_24[19]},
      {stage1_24[12]}
   );
   gpc1_1 gpc141 (
      {stage0_24[20]},
      {stage1_24[13]}
   );
   gpc1_1 gpc142 (
      {stage0_24[21]},
      {stage1_24[14]}
   );
   gpc1_1 gpc143 (
      {stage0_24[22]},
      {stage1_24[15]}
   );
   gpc1_1 gpc144 (
      {stage0_24[23]},
      {stage1_24[16]}
   );
   gpc1_1 gpc145 (
      {stage0_24[24]},
      {stage1_24[17]}
   );
   gpc1_1 gpc146 (
      {stage0_25[14]},
      {stage1_25[8]}
   );
   gpc1_1 gpc147 (
      {stage0_25[15]},
      {stage1_25[9]}
   );
   gpc1_1 gpc148 (
      {stage0_25[16]},
      {stage1_25[10]}
   );
   gpc1_1 gpc149 (
      {stage0_25[17]},
      {stage1_25[11]}
   );
   gpc1_1 gpc150 (
      {stage0_25[18]},
      {stage1_25[12]}
   );
   gpc1_1 gpc151 (
      {stage0_25[19]},
      {stage1_25[13]}
   );
   gpc1_1 gpc152 (
      {stage0_25[20]},
      {stage1_25[14]}
   );
   gpc1_1 gpc153 (
      {stage0_25[21]},
      {stage1_25[15]}
   );
   gpc1_1 gpc154 (
      {stage0_25[22]},
      {stage1_25[16]}
   );
   gpc1_1 gpc155 (
      {stage0_25[23]},
      {stage1_25[17]}
   );
   gpc1_1 gpc156 (
      {stage0_25[24]},
      {stage1_25[18]}
   );
   gpc1_1 gpc157 (
      {stage0_25[25]},
      {stage1_25[19]}
   );
   gpc1_1 gpc158 (
      {stage0_26[22]},
      {stage1_26[7]}
   );
   gpc1_1 gpc159 (
      {stage0_26[23]},
      {stage1_26[8]}
   );
   gpc1_1 gpc160 (
      {stage0_26[24]},
      {stage1_26[9]}
   );
   gpc1_1 gpc161 (
      {stage0_26[25]},
      {stage1_26[10]}
   );
   gpc1_1 gpc162 (
      {stage0_26[26]},
      {stage1_26[11]}
   );
   gpc1_1 gpc163 (
      {stage0_27[18]},
      {stage1_27[8]}
   );
   gpc1_1 gpc164 (
      {stage0_27[19]},
      {stage1_27[9]}
   );
   gpc1_1 gpc165 (
      {stage0_27[20]},
      {stage1_27[10]}
   );
   gpc1_1 gpc166 (
      {stage0_27[21]},
      {stage1_27[11]}
   );
   gpc1_1 gpc167 (
      {stage0_27[22]},
      {stage1_27[12]}
   );
   gpc1_1 gpc168 (
      {stage0_27[23]},
      {stage1_27[13]}
   );
   gpc1_1 gpc169 (
      {stage0_27[24]},
      {stage1_27[14]}
   );
   gpc1_1 gpc170 (
      {stage0_27[25]},
      {stage1_27[15]}
   );
   gpc1_1 gpc171 (
      {stage0_27[26]},
      {stage1_27[16]}
   );
   gpc1_1 gpc172 (
      {stage0_27[27]},
      {stage1_27[17]}
   );
   gpc1_1 gpc173 (
      {stage0_28[26]},
      {stage1_28[9]}
   );
   gpc1_1 gpc174 (
      {stage0_28[27]},
      {stage1_28[10]}
   );
   gpc1_1 gpc175 (
      {stage0_28[28]},
      {stage1_28[11]}
   );
   gpc1_1 gpc176 (
      {stage0_29[27]},
      {stage1_29[10]}
   );
   gpc1_1 gpc177 (
      {stage0_29[28]},
      {stage1_29[11]}
   );
   gpc1_1 gpc178 (
      {stage0_29[29]},
      {stage1_29[12]}
   );
   gpc1_1 gpc179 (
      {stage0_30[28]},
      {stage1_30[12]}
   );
   gpc1_1 gpc180 (
      {stage0_31[25]},
      {stage1_31[11]}
   );
   gpc1_1 gpc181 (
      {stage0_31[26]},
      {stage1_31[12]}
   );
   gpc1_1 gpc182 (
      {stage0_31[27]},
      {stage1_31[13]}
   );
   gpc1_1 gpc183 (
      {stage0_32[24]},
      {stage1_32[10]}
   );
   gpc1_1 gpc184 (
      {stage0_32[25]},
      {stage1_32[11]}
   );
   gpc1_1 gpc185 (
      {stage0_32[26]},
      {stage1_32[12]}
   );
   gpc1_1 gpc186 (
      {stage0_33[13]},
      {stage1_33[9]}
   );
   gpc1_1 gpc187 (
      {stage0_33[14]},
      {stage1_33[10]}
   );
   gpc1_1 gpc188 (
      {stage0_33[15]},
      {stage1_33[11]}
   );
   gpc1_1 gpc189 (
      {stage0_33[16]},
      {stage1_33[12]}
   );
   gpc1_1 gpc190 (
      {stage0_33[17]},
      {stage1_33[13]}
   );
   gpc1_1 gpc191 (
      {stage0_33[18]},
      {stage1_33[14]}
   );
   gpc1_1 gpc192 (
      {stage0_33[19]},
      {stage1_33[15]}
   );
   gpc1_1 gpc193 (
      {stage0_33[20]},
      {stage1_33[16]}
   );
   gpc1_1 gpc194 (
      {stage0_33[21]},
      {stage1_33[17]}
   );
   gpc1_1 gpc195 (
      {stage0_33[22]},
      {stage1_33[18]}
   );
   gpc1_1 gpc196 (
      {stage0_33[23]},
      {stage1_33[19]}
   );
   gpc1_1 gpc197 (
      {stage0_33[24]},
      {stage1_33[20]}
   );
   gpc1_1 gpc198 (
      {stage0_33[25]},
      {stage1_33[21]}
   );
   gpc1_1 gpc199 (
      {stage0_34[18]},
      {stage1_34[8]}
   );
   gpc1_1 gpc200 (
      {stage0_34[19]},
      {stage1_34[9]}
   );
   gpc1_1 gpc201 (
      {stage0_34[20]},
      {stage1_34[10]}
   );
   gpc1_1 gpc202 (
      {stage0_34[21]},
      {stage1_34[11]}
   );
   gpc1_1 gpc203 (
      {stage0_34[22]},
      {stage1_34[12]}
   );
   gpc1_1 gpc204 (
      {stage0_34[23]},
      {stage1_34[13]}
   );
   gpc1_1 gpc205 (
      {stage0_34[24]},
      {stage1_34[14]}
   );
   gpc1_1 gpc206 (
      {stage0_35[12]},
      {stage1_35[6]}
   );
   gpc1_1 gpc207 (
      {stage0_35[13]},
      {stage1_35[7]}
   );
   gpc1_1 gpc208 (
      {stage0_35[14]},
      {stage1_35[8]}
   );
   gpc1_1 gpc209 (
      {stage0_35[15]},
      {stage1_35[9]}
   );
   gpc1_1 gpc210 (
      {stage0_35[16]},
      {stage1_35[10]}
   );
   gpc1_1 gpc211 (
      {stage0_35[17]},
      {stage1_35[11]}
   );
   gpc1_1 gpc212 (
      {stage0_35[18]},
      {stage1_35[12]}
   );
   gpc1_1 gpc213 (
      {stage0_35[19]},
      {stage1_35[13]}
   );
   gpc1_1 gpc214 (
      {stage0_35[20]},
      {stage1_35[14]}
   );
   gpc1_1 gpc215 (
      {stage0_35[21]},
      {stage1_35[15]}
   );
   gpc1_1 gpc216 (
      {stage0_35[22]},
      {stage1_35[16]}
   );
   gpc1_1 gpc217 (
      {stage0_35[23]},
      {stage1_35[17]}
   );
   gpc1_1 gpc218 (
      {stage0_36[22]},
      {stage1_36[7]}
   );
   gpc1_1 gpc219 (
      {stage0_37[8]},
      {stage1_37[6]}
   );
   gpc1_1 gpc220 (
      {stage0_37[9]},
      {stage1_37[7]}
   );
   gpc1_1 gpc221 (
      {stage0_37[10]},
      {stage1_37[8]}
   );
   gpc1_1 gpc222 (
      {stage0_37[11]},
      {stage1_37[9]}
   );
   gpc1_1 gpc223 (
      {stage0_37[12]},
      {stage1_37[10]}
   );
   gpc1_1 gpc224 (
      {stage0_37[13]},
      {stage1_37[11]}
   );
   gpc1_1 gpc225 (
      {stage0_37[14]},
      {stage1_37[12]}
   );
   gpc1_1 gpc226 (
      {stage0_37[15]},
      {stage1_37[13]}
   );
   gpc1_1 gpc227 (
      {stage0_37[16]},
      {stage1_37[14]}
   );
   gpc1_1 gpc228 (
      {stage0_37[17]},
      {stage1_37[15]}
   );
   gpc1_1 gpc229 (
      {stage0_37[18]},
      {stage1_37[16]}
   );
   gpc1_1 gpc230 (
      {stage0_37[19]},
      {stage1_37[17]}
   );
   gpc1_1 gpc231 (
      {stage0_37[20]},
      {stage1_37[18]}
   );
   gpc1_1 gpc232 (
      {stage0_37[21]},
      {stage1_37[19]}
   );
   gpc1_1 gpc233 (
      {stage0_38[17]},
      {stage1_38[6]}
   );
   gpc1_1 gpc234 (
      {stage0_38[18]},
      {stage1_38[7]}
   );
   gpc1_1 gpc235 (
      {stage0_38[19]},
      {stage1_38[8]}
   );
   gpc1_1 gpc236 (
      {stage0_38[20]},
      {stage1_38[9]}
   );
   gpc1_1 gpc237 (
      {stage0_39[6]},
      {stage1_39[5]}
   );
   gpc1_1 gpc238 (
      {stage0_39[7]},
      {stage1_39[6]}
   );
   gpc1_1 gpc239 (
      {stage0_39[8]},
      {stage1_39[7]}
   );
   gpc1_1 gpc240 (
      {stage0_39[9]},
      {stage1_39[8]}
   );
   gpc1_1 gpc241 (
      {stage0_39[10]},
      {stage1_39[9]}
   );
   gpc1_1 gpc242 (
      {stage0_39[11]},
      {stage1_39[10]}
   );
   gpc1_1 gpc243 (
      {stage0_39[12]},
      {stage1_39[11]}
   );
   gpc1_1 gpc244 (
      {stage0_39[13]},
      {stage1_39[12]}
   );
   gpc1_1 gpc245 (
      {stage0_39[14]},
      {stage1_39[13]}
   );
   gpc1_1 gpc246 (
      {stage0_39[15]},
      {stage1_39[14]}
   );
   gpc1_1 gpc247 (
      {stage0_39[16]},
      {stage1_39[15]}
   );
   gpc1_1 gpc248 (
      {stage0_39[17]},
      {stage1_39[16]}
   );
   gpc1_1 gpc249 (
      {stage0_39[18]},
      {stage1_39[17]}
   );
   gpc1_1 gpc250 (
      {stage0_39[19]},
      {stage1_39[18]}
   );
   gpc1_1 gpc251 (
      {stage0_40[13]},
      {stage1_40[6]}
   );
   gpc1_1 gpc252 (
      {stage0_40[14]},
      {stage1_40[7]}
   );
   gpc1_1 gpc253 (
      {stage0_40[15]},
      {stage1_40[8]}
   );
   gpc1_1 gpc254 (
      {stage0_40[16]},
      {stage1_40[9]}
   );
   gpc1_1 gpc255 (
      {stage0_40[17]},
      {stage1_40[10]}
   );
   gpc1_1 gpc256 (
      {stage0_40[18]},
      {stage1_40[11]}
   );
   gpc1_1 gpc257 (
      {stage0_41[14]},
      {stage1_41[4]}
   );
   gpc1_1 gpc258 (
      {stage0_41[15]},
      {stage1_41[5]}
   );
   gpc1_1 gpc259 (
      {stage0_41[16]},
      {stage1_41[6]}
   );
   gpc1_1 gpc260 (
      {stage0_41[17]},
      {stage1_41[7]}
   );
   gpc1_1 gpc261 (
      {stage0_43[8]},
      {stage1_43[6]}
   );
   gpc1_1 gpc262 (
      {stage0_43[9]},
      {stage1_43[7]}
   );
   gpc1_1 gpc263 (
      {stage0_43[10]},
      {stage1_43[8]}
   );
   gpc1_1 gpc264 (
      {stage0_43[11]},
      {stage1_43[9]}
   );
   gpc1_1 gpc265 (
      {stage0_43[12]},
      {stage1_43[10]}
   );
   gpc1_1 gpc266 (
      {stage0_43[13]},
      {stage1_43[11]}
   );
   gpc1_1 gpc267 (
      {stage0_43[14]},
      {stage1_43[12]}
   );
   gpc1_1 gpc268 (
      {stage0_43[15]},
      {stage1_43[13]}
   );
   gpc1_1 gpc269 (
      {stage0_44[12]},
      {stage1_44[5]}
   );
   gpc1_1 gpc270 (
      {stage0_44[13]},
      {stage1_44[6]}
   );
   gpc1_1 gpc271 (
      {stage0_44[14]},
      {stage1_44[7]}
   );
   gpc1_1 gpc272 (
      {stage0_45[12]},
      {stage1_45[4]}
   );
   gpc1_1 gpc273 (
      {stage0_45[13]},
      {stage1_45[5]}
   );
   gpc1_1 gpc274 (
      {stage0_46[0]},
      {stage1_46[4]}
   );
   gpc1_1 gpc275 (
      {stage0_46[1]},
      {stage1_46[5]}
   );
   gpc1_1 gpc276 (
      {stage0_46[2]},
      {stage1_46[6]}
   );
   gpc1_1 gpc277 (
      {stage0_46[3]},
      {stage1_46[7]}
   );
   gpc1_1 gpc278 (
      {stage0_46[4]},
      {stage1_46[8]}
   );
   gpc1_1 gpc279 (
      {stage0_46[5]},
      {stage1_46[9]}
   );
   gpc1_1 gpc280 (
      {stage0_46[6]},
      {stage1_46[10]}
   );
   gpc1_1 gpc281 (
      {stage0_46[7]},
      {stage1_46[11]}
   );
   gpc1_1 gpc282 (
      {stage0_46[8]},
      {stage1_46[12]}
   );
   gpc1_1 gpc283 (
      {stage0_46[9]},
      {stage1_46[13]}
   );
   gpc1_1 gpc284 (
      {stage0_46[10]},
      {stage1_46[14]}
   );
   gpc1_1 gpc285 (
      {stage0_46[11]},
      {stage1_46[15]}
   );
   gpc1_1 gpc286 (
      {stage0_46[12]},
      {stage1_46[16]}
   );
   gpc1_1 gpc287 (
      {stage0_47[6]},
      {stage1_47[2]}
   );
   gpc1_1 gpc288 (
      {stage0_47[7]},
      {stage1_47[3]}
   );
   gpc1_1 gpc289 (
      {stage0_47[8]},
      {stage1_47[4]}
   );
   gpc1_1 gpc290 (
      {stage0_47[9]},
      {stage1_47[5]}
   );
   gpc1_1 gpc291 (
      {stage0_47[10]},
      {stage1_47[6]}
   );
   gpc1_1 gpc292 (
      {stage0_47[11]},
      {stage1_47[7]}
   );
   gpc1_1 gpc293 (
      {stage0_48[0]},
      {stage1_48[1]}
   );
   gpc1_1 gpc294 (
      {stage0_48[1]},
      {stage1_48[2]}
   );
   gpc1_1 gpc295 (
      {stage0_48[2]},
      {stage1_48[3]}
   );
   gpc1_1 gpc296 (
      {stage0_48[3]},
      {stage1_48[4]}
   );
   gpc1_1 gpc297 (
      {stage0_48[4]},
      {stage1_48[5]}
   );
   gpc1_1 gpc298 (
      {stage0_48[5]},
      {stage1_48[6]}
   );
   gpc1_1 gpc299 (
      {stage0_48[6]},
      {stage1_48[7]}
   );
   gpc1_1 gpc300 (
      {stage0_48[7]},
      {stage1_48[8]}
   );
   gpc1_1 gpc301 (
      {stage0_48[8]},
      {stage1_48[9]}
   );
   gpc1_1 gpc302 (
      {stage0_48[9]},
      {stage1_48[10]}
   );
   gpc1_1 gpc303 (
      {stage0_48[10]},
      {stage1_48[11]}
   );
   gpc1_1 gpc304 (
      {stage0_49[5]},
      {stage1_49[2]}
   );
   gpc1_1 gpc305 (
      {stage0_49[6]},
      {stage1_49[3]}
   );
   gpc1_1 gpc306 (
      {stage0_49[7]},
      {stage1_49[4]}
   );
   gpc1_1 gpc307 (
      {stage0_49[8]},
      {stage1_49[5]}
   );
   gpc1_1 gpc308 (
      {stage0_49[9]},
      {stage1_49[6]}
   );
   gpc1_1 gpc309 (
      {stage0_50[1]},
      {stage1_50[1]}
   );
   gpc1_1 gpc310 (
      {stage0_50[2]},
      {stage1_50[2]}
   );
   gpc1_1 gpc311 (
      {stage0_50[3]},
      {stage1_50[3]}
   );
   gpc1_1 gpc312 (
      {stage0_50[4]},
      {stage1_50[4]}
   );
   gpc1_1 gpc313 (
      {stage0_50[5]},
      {stage1_50[5]}
   );
   gpc1_1 gpc314 (
      {stage0_50[6]},
      {stage1_50[6]}
   );
   gpc1_1 gpc315 (
      {stage0_50[7]},
      {stage1_50[7]}
   );
   gpc1_1 gpc316 (
      {stage0_50[8]},
      {stage1_50[8]}
   );
   gpc1_1 gpc317 (
      {stage0_51[6]},
      {stage1_51[1]}
   );
   gpc1_1 gpc318 (
      {stage0_51[7]},
      {stage1_51[2]}
   );
   gpc1_1 gpc319 (
      {stage0_52[0]},
      {stage1_52[1]}
   );
   gpc1_1 gpc320 (
      {stage0_52[1]},
      {stage1_52[2]}
   );
   gpc1_1 gpc321 (
      {stage0_52[2]},
      {stage1_52[3]}
   );
   gpc1_1 gpc322 (
      {stage0_52[3]},
      {stage1_52[4]}
   );
   gpc1_1 gpc323 (
      {stage0_52[4]},
      {stage1_52[5]}
   );
   gpc1_1 gpc324 (
      {stage0_52[5]},
      {stage1_52[6]}
   );
   gpc1_1 gpc325 (
      {stage0_52[6]},
      {stage1_52[7]}
   );
   gpc1_1 gpc326 (
      {stage0_53[0]},
      {stage1_53[1]}
   );
   gpc1_1 gpc327 (
      {stage0_53[1]},
      {stage1_53[2]}
   );
   gpc1_1 gpc328 (
      {stage0_53[2]},
      {stage1_53[3]}
   );
   gpc1_1 gpc329 (
      {stage0_53[3]},
      {stage1_53[4]}
   );
   gpc1_1 gpc330 (
      {stage0_53[4]},
      {stage1_53[5]}
   );
   gpc1_1 gpc331 (
      {stage0_53[5]},
      {stage1_53[6]}
   );
   gpc1_1 gpc332 (
      {stage0_54[0]},
      {stage1_54[0]}
   );
   gpc1_1 gpc333 (
      {stage0_54[1]},
      {stage1_54[1]}
   );
   gpc1_1 gpc334 (
      {stage0_54[2]},
      {stage1_54[2]}
   );
   gpc1_1 gpc335 (
      {stage0_54[3]},
      {stage1_54[3]}
   );
   gpc1_1 gpc336 (
      {stage0_54[4]},
      {stage1_54[4]}
   );
   gpc1_1 gpc337 (
      {stage0_55[0]},
      {stage1_55[0]}
   );
   gpc1_1 gpc338 (
      {stage0_55[1]},
      {stage1_55[1]}
   );
   gpc1_1 gpc339 (
      {stage0_55[2]},
      {stage1_55[2]}
   );
   gpc1_1 gpc340 (
      {stage0_55[3]},
      {stage1_55[3]}
   );
   gpc1_1 gpc341 (
      {stage0_56[0]},
      {stage1_56[0]}
   );
   gpc1_1 gpc342 (
      {stage0_56[1]},
      {stage1_56[1]}
   );
   gpc1_1 gpc343 (
      {stage0_56[2]},
      {stage1_56[2]}
   );
   gpc1_1 gpc344 (
      {stage0_57[0]},
      {stage1_57[0]}
   );
   gpc1_1 gpc345 (
      {stage0_57[1]},
      {stage1_57[1]}
   );
   gpc1_1 gpc346 (
      {stage0_58[0]},
      {stage1_58[0]}
   );
   gpc433_5 gpc347 (
      {stage1_2[0], stage1_2[1], stage1_2[2]},
      {stage1_3[0], stage1_3[1], stage1_3[2]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3]},
      {stage2_6[0],stage2_5[0],stage2_4[0],stage2_3[0],stage2_2[0]}
   );
   gpc1334_5 gpc348 (
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3]},
      {stage1_7[0], stage1_7[1], stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2]},
      {stage1_9[0]},
      {stage2_10[0],stage2_9[0],stage2_8[0],stage2_7[0],stage2_6[1]}
   );
   gpc606_5 gpc349 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[1]}
   );
   gpc606_5 gpc350 (
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[0],stage2_14[1],stage2_13[1]}
   );
   gpc606_5 gpc351 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[1],stage2_14[2]}
   );
   gpc606_5 gpc352 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[0],stage2_19[0],stage2_18[1],stage2_17[2]}
   );
   gpc623_5 gpc353 (
      {stage1_17[6], stage1_17[7], stage1_17[8]},
      {stage1_18[0], stage1_18[1]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[1],stage2_19[1],stage2_18[2],stage2_17[3]}
   );
   gpc615_5 gpc354 (
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[2],stage2_20[2],stage2_19[2]}
   );
   gpc606_5 gpc355 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[0],stage2_24[0],stage2_23[1],stage2_22[1]}
   );
   gpc615_5 gpc356 (
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4]},
      {stage1_24[6]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[1],stage2_25[1],stage2_24[1],stage2_23[2]}
   );
   gpc615_5 gpc357 (
      {stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage1_25[6]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[1],stage2_26[2],stage2_25[2],stage2_24[2]}
   );
   gpc615_5 gpc358 (
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16]},
      {stage1_25[7]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[2],stage2_26[3],stage2_25[3],stage2_24[3]}
   );
   gpc606_5 gpc359 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[3],stage2_26[4],stage2_25[4]}
   );
   gpc606_5 gpc360 (
      {stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18], stage1_25[19]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[3],stage2_27[4],stage2_26[5],stage2_25[5]}
   );
   gpc606_5 gpc361 (
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[0],stage2_29[2],stage2_28[4],stage2_27[5]}
   );
   gpc615_5 gpc362 (
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4]},
      {stage1_29[6]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[1],stage2_30[1],stage2_29[3],stage2_28[5]}
   );
   gpc615_5 gpc363 (
      {stage1_28[5], stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9]},
      {stage1_29[7]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[2],stage2_30[2],stage2_29[4],stage2_28[6]}
   );
   gpc615_5 gpc364 (
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11], stage1_29[12]},
      {stage1_30[12]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[2],stage2_31[3],stage2_30[3],stage2_29[5]}
   );
   gpc606_5 gpc365 (
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[0],stage2_34[0],stage2_33[1],stage2_32[3]}
   );
   gpc606_5 gpc366 (
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[1],stage2_34[1],stage2_33[2],stage2_32[4]}
   );
   gpc615_5 gpc367 (
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4]},
      {stage1_34[12]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[2],stage2_35[2],stage2_34[2],stage2_33[3]}
   );
   gpc615_5 gpc368 (
      {stage1_33[5], stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9]},
      {stage1_34[13]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[3],stage2_35[3],stage2_34[3],stage2_33[4]}
   );
   gpc615_5 gpc369 (
      {stage1_33[10], stage1_33[11], stage1_33[12], stage1_33[13], stage1_33[14]},
      {stage1_34[14]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[4],stage2_35[4],stage2_34[4],stage2_33[5]}
   );
   gpc1244_5 gpc370 (
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3]},
      {stage1_38[0], stage1_38[1]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[0],stage2_38[0],stage2_37[3],stage2_36[5]}
   );
   gpc606_5 gpc371 (
      {stage1_37[4], stage1_37[5], stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[1],stage2_39[1],stage2_38[1],stage2_37[4]}
   );
   gpc615_5 gpc372 (
      {stage1_37[10], stage1_37[11], stage1_37[12], stage1_37[13], stage1_37[14]},
      {stage1_38[2]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[2],stage2_39[2],stage2_38[2],stage2_37[5]}
   );
   gpc615_5 gpc373 (
      {stage1_37[15], stage1_37[16], stage1_37[17], stage1_37[18], stage1_37[19]},
      {stage1_38[3]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[3],stage2_39[3],stage2_38[3],stage2_37[6]}
   );
   gpc606_5 gpc374 (
      {stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[3],stage2_40[4],stage2_39[4],stage2_38[4]}
   );
   gpc615_5 gpc375 (
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10]},
      {stage1_41[0]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[1],stage2_41[4],stage2_40[5]}
   );
   gpc606_5 gpc376 (
      {stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5], stage1_41[6]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[1],stage2_43[1],stage2_42[2],stage2_41[5]}
   );
   gpc615_5 gpc377 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[0]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[0],stage2_46[0],stage2_45[1],stage2_44[2]}
   );
   gpc425_5 gpc378 (
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10]},
      {stage1_47[0], stage1_47[1]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3]},
      {stage2_50[0],stage2_49[0],stage2_48[1],stage2_47[1],stage2_46[1]}
   );
   gpc623_5 gpc379 (
      {stage1_47[2], stage1_47[3], stage1_47[4]},
      {stage1_48[4], stage1_48[5]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[1],stage2_49[1],stage2_48[2],stage2_47[2]}
   );
   gpc606_5 gpc380 (
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage1_52[0], stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5]},
      {stage2_54[0],stage2_53[0],stage2_52[0],stage2_51[1],stage2_50[2]}
   );
   gpc1423_5 gpc381 (
      {stage1_53[0], stage1_53[1], stage1_53[2]},
      {stage1_54[0], stage1_54[1]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3]},
      {stage1_56[0]},
      {stage2_57[0],stage2_56[0],stage2_55[0],stage2_54[1],stage2_53[1]}
   );
   gpc1_1 gpc382 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc383 (
      {stage1_1[0]},
      {stage2_1[0]}
   );
   gpc1_1 gpc384 (
      {stage1_1[1]},
      {stage2_1[1]}
   );
   gpc1_1 gpc385 (
      {stage1_3[3]},
      {stage2_3[1]}
   );
   gpc1_1 gpc386 (
      {stage1_4[4]},
      {stage2_4[1]}
   );
   gpc1_1 gpc387 (
      {stage1_5[0]},
      {stage2_5[1]}
   );
   gpc1_1 gpc388 (
      {stage1_6[4]},
      {stage2_6[2]}
   );
   gpc1_1 gpc389 (
      {stage1_6[5]},
      {stage2_6[3]}
   );
   gpc1_1 gpc390 (
      {stage1_6[6]},
      {stage2_6[4]}
   );
   gpc1_1 gpc391 (
      {stage1_6[7]},
      {stage2_6[5]}
   );
   gpc1_1 gpc392 (
      {stage1_8[3]},
      {stage2_8[1]}
   );
   gpc1_1 gpc393 (
      {stage1_8[4]},
      {stage2_8[2]}
   );
   gpc1_1 gpc394 (
      {stage1_8[5]},
      {stage2_8[3]}
   );
   gpc1_1 gpc395 (
      {stage1_8[6]},
      {stage2_8[4]}
   );
   gpc1_1 gpc396 (
      {stage1_8[7]},
      {stage2_8[5]}
   );
   gpc1_1 gpc397 (
      {stage1_8[8]},
      {stage2_8[6]}
   );
   gpc1_1 gpc398 (
      {stage1_8[9]},
      {stage2_8[7]}
   );
   gpc1_1 gpc399 (
      {stage1_9[1]},
      {stage2_9[1]}
   );
   gpc1_1 gpc400 (
      {stage1_9[2]},
      {stage2_9[2]}
   );
   gpc1_1 gpc401 (
      {stage1_9[3]},
      {stage2_9[3]}
   );
   gpc1_1 gpc402 (
      {stage1_9[4]},
      {stage2_9[4]}
   );
   gpc1_1 gpc403 (
      {stage1_9[5]},
      {stage2_9[5]}
   );
   gpc1_1 gpc404 (
      {stage1_9[6]},
      {stage2_9[6]}
   );
   gpc1_1 gpc405 (
      {stage1_10[6]},
      {stage2_10[2]}
   );
   gpc1_1 gpc406 (
      {stage1_10[7]},
      {stage2_10[3]}
   );
   gpc1_1 gpc407 (
      {stage1_10[8]},
      {stage2_10[4]}
   );
   gpc1_1 gpc408 (
      {stage1_10[9]},
      {stage2_10[5]}
   );
   gpc1_1 gpc409 (
      {stage1_11[0]},
      {stage2_11[1]}
   );
   gpc1_1 gpc410 (
      {stage1_11[1]},
      {stage2_11[2]}
   );
   gpc1_1 gpc411 (
      {stage1_11[2]},
      {stage2_11[3]}
   );
   gpc1_1 gpc412 (
      {stage1_11[3]},
      {stage2_11[4]}
   );
   gpc1_1 gpc413 (
      {stage1_11[4]},
      {stage2_11[5]}
   );
   gpc1_1 gpc414 (
      {stage1_16[6]},
      {stage2_16[2]}
   );
   gpc1_1 gpc415 (
      {stage1_16[7]},
      {stage2_16[3]}
   );
   gpc1_1 gpc416 (
      {stage1_16[8]},
      {stage2_16[4]}
   );
   gpc1_1 gpc417 (
      {stage1_18[2]},
      {stage2_18[3]}
   );
   gpc1_1 gpc418 (
      {stage1_18[3]},
      {stage2_18[4]}
   );
   gpc1_1 gpc419 (
      {stage1_18[4]},
      {stage2_18[5]}
   );
   gpc1_1 gpc420 (
      {stage1_18[5]},
      {stage2_18[6]}
   );
   gpc1_1 gpc421 (
      {stage1_19[17]},
      {stage2_19[3]}
   );
   gpc1_1 gpc422 (
      {stage1_19[18]},
      {stage2_19[4]}
   );
   gpc1_1 gpc423 (
      {stage1_19[19]},
      {stage2_19[5]}
   );
   gpc1_1 gpc424 (
      {stage1_19[20]},
      {stage2_19[6]}
   );
   gpc1_1 gpc425 (
      {stage1_20[1]},
      {stage2_20[3]}
   );
   gpc1_1 gpc426 (
      {stage1_20[2]},
      {stage2_20[4]}
   );
   gpc1_1 gpc427 (
      {stage1_20[3]},
      {stage2_20[5]}
   );
   gpc1_1 gpc428 (
      {stage1_20[4]},
      {stage2_20[6]}
   );
   gpc1_1 gpc429 (
      {stage1_20[5]},
      {stage2_20[7]}
   );
   gpc1_1 gpc430 (
      {stage1_20[6]},
      {stage2_20[8]}
   );
   gpc1_1 gpc431 (
      {stage1_20[7]},
      {stage2_20[9]}
   );
   gpc1_1 gpc432 (
      {stage1_20[8]},
      {stage2_20[10]}
   );
   gpc1_1 gpc433 (
      {stage1_20[9]},
      {stage2_20[11]}
   );
   gpc1_1 gpc434 (
      {stage1_20[10]},
      {stage2_20[12]}
   );
   gpc1_1 gpc435 (
      {stage1_20[11]},
      {stage2_20[13]}
   );
   gpc1_1 gpc436 (
      {stage1_20[12]},
      {stage2_20[14]}
   );
   gpc1_1 gpc437 (
      {stage1_20[13]},
      {stage2_20[15]}
   );
   gpc1_1 gpc438 (
      {stage1_22[6]},
      {stage2_22[2]}
   );
   gpc1_1 gpc439 (
      {stage1_22[7]},
      {stage2_22[3]}
   );
   gpc1_1 gpc440 (
      {stage1_22[8]},
      {stage2_22[4]}
   );
   gpc1_1 gpc441 (
      {stage1_22[9]},
      {stage2_22[5]}
   );
   gpc1_1 gpc442 (
      {stage1_23[5]},
      {stage2_23[3]}
   );
   gpc1_1 gpc443 (
      {stage1_23[6]},
      {stage2_23[4]}
   );
   gpc1_1 gpc444 (
      {stage1_23[7]},
      {stage2_23[5]}
   );
   gpc1_1 gpc445 (
      {stage1_24[17]},
      {stage2_24[4]}
   );
   gpc1_1 gpc446 (
      {stage1_28[10]},
      {stage2_28[7]}
   );
   gpc1_1 gpc447 (
      {stage1_28[11]},
      {stage2_28[8]}
   );
   gpc1_1 gpc448 (
      {stage1_31[6]},
      {stage2_31[4]}
   );
   gpc1_1 gpc449 (
      {stage1_31[7]},
      {stage2_31[5]}
   );
   gpc1_1 gpc450 (
      {stage1_31[8]},
      {stage2_31[6]}
   );
   gpc1_1 gpc451 (
      {stage1_31[9]},
      {stage2_31[7]}
   );
   gpc1_1 gpc452 (
      {stage1_31[10]},
      {stage2_31[8]}
   );
   gpc1_1 gpc453 (
      {stage1_31[11]},
      {stage2_31[9]}
   );
   gpc1_1 gpc454 (
      {stage1_31[12]},
      {stage2_31[10]}
   );
   gpc1_1 gpc455 (
      {stage1_31[13]},
      {stage2_31[11]}
   );
   gpc1_1 gpc456 (
      {stage1_32[12]},
      {stage2_32[5]}
   );
   gpc1_1 gpc457 (
      {stage1_33[15]},
      {stage2_33[6]}
   );
   gpc1_1 gpc458 (
      {stage1_33[16]},
      {stage2_33[7]}
   );
   gpc1_1 gpc459 (
      {stage1_33[17]},
      {stage2_33[8]}
   );
   gpc1_1 gpc460 (
      {stage1_33[18]},
      {stage2_33[9]}
   );
   gpc1_1 gpc461 (
      {stage1_33[19]},
      {stage2_33[10]}
   );
   gpc1_1 gpc462 (
      {stage1_33[20]},
      {stage2_33[11]}
   );
   gpc1_1 gpc463 (
      {stage1_33[21]},
      {stage2_33[12]}
   );
   gpc1_1 gpc464 (
      {stage1_36[4]},
      {stage2_36[6]}
   );
   gpc1_1 gpc465 (
      {stage1_36[5]},
      {stage2_36[7]}
   );
   gpc1_1 gpc466 (
      {stage1_36[6]},
      {stage2_36[8]}
   );
   gpc1_1 gpc467 (
      {stage1_36[7]},
      {stage2_36[9]}
   );
   gpc1_1 gpc468 (
      {stage1_40[11]},
      {stage2_40[6]}
   );
   gpc1_1 gpc469 (
      {stage1_41[7]},
      {stage2_41[6]}
   );
   gpc1_1 gpc470 (
      {stage1_43[6]},
      {stage2_43[2]}
   );
   gpc1_1 gpc471 (
      {stage1_43[7]},
      {stage2_43[3]}
   );
   gpc1_1 gpc472 (
      {stage1_43[8]},
      {stage2_43[4]}
   );
   gpc1_1 gpc473 (
      {stage1_43[9]},
      {stage2_43[5]}
   );
   gpc1_1 gpc474 (
      {stage1_43[10]},
      {stage2_43[6]}
   );
   gpc1_1 gpc475 (
      {stage1_43[11]},
      {stage2_43[7]}
   );
   gpc1_1 gpc476 (
      {stage1_43[12]},
      {stage2_43[8]}
   );
   gpc1_1 gpc477 (
      {stage1_43[13]},
      {stage2_43[9]}
   );
   gpc1_1 gpc478 (
      {stage1_44[5]},
      {stage2_44[3]}
   );
   gpc1_1 gpc479 (
      {stage1_44[6]},
      {stage2_44[4]}
   );
   gpc1_1 gpc480 (
      {stage1_44[7]},
      {stage2_44[5]}
   );
   gpc1_1 gpc481 (
      {stage1_45[1]},
      {stage2_45[2]}
   );
   gpc1_1 gpc482 (
      {stage1_45[2]},
      {stage2_45[3]}
   );
   gpc1_1 gpc483 (
      {stage1_45[3]},
      {stage2_45[4]}
   );
   gpc1_1 gpc484 (
      {stage1_45[4]},
      {stage2_45[5]}
   );
   gpc1_1 gpc485 (
      {stage1_45[5]},
      {stage2_45[6]}
   );
   gpc1_1 gpc486 (
      {stage1_46[11]},
      {stage2_46[2]}
   );
   gpc1_1 gpc487 (
      {stage1_46[12]},
      {stage2_46[3]}
   );
   gpc1_1 gpc488 (
      {stage1_46[13]},
      {stage2_46[4]}
   );
   gpc1_1 gpc489 (
      {stage1_46[14]},
      {stage2_46[5]}
   );
   gpc1_1 gpc490 (
      {stage1_46[15]},
      {stage2_46[6]}
   );
   gpc1_1 gpc491 (
      {stage1_46[16]},
      {stage2_46[7]}
   );
   gpc1_1 gpc492 (
      {stage1_47[5]},
      {stage2_47[3]}
   );
   gpc1_1 gpc493 (
      {stage1_47[6]},
      {stage2_47[4]}
   );
   gpc1_1 gpc494 (
      {stage1_47[7]},
      {stage2_47[5]}
   );
   gpc1_1 gpc495 (
      {stage1_48[6]},
      {stage2_48[3]}
   );
   gpc1_1 gpc496 (
      {stage1_48[7]},
      {stage2_48[4]}
   );
   gpc1_1 gpc497 (
      {stage1_48[8]},
      {stage2_48[5]}
   );
   gpc1_1 gpc498 (
      {stage1_48[9]},
      {stage2_48[6]}
   );
   gpc1_1 gpc499 (
      {stage1_48[10]},
      {stage2_48[7]}
   );
   gpc1_1 gpc500 (
      {stage1_48[11]},
      {stage2_48[8]}
   );
   gpc1_1 gpc501 (
      {stage1_49[6]},
      {stage2_49[2]}
   );
   gpc1_1 gpc502 (
      {stage1_50[6]},
      {stage2_50[3]}
   );
   gpc1_1 gpc503 (
      {stage1_50[7]},
      {stage2_50[4]}
   );
   gpc1_1 gpc504 (
      {stage1_50[8]},
      {stage2_50[5]}
   );
   gpc1_1 gpc505 (
      {stage1_51[0]},
      {stage2_51[2]}
   );
   gpc1_1 gpc506 (
      {stage1_51[1]},
      {stage2_51[3]}
   );
   gpc1_1 gpc507 (
      {stage1_51[2]},
      {stage2_51[4]}
   );
   gpc1_1 gpc508 (
      {stage1_52[6]},
      {stage2_52[1]}
   );
   gpc1_1 gpc509 (
      {stage1_52[7]},
      {stage2_52[2]}
   );
   gpc1_1 gpc510 (
      {stage1_53[3]},
      {stage2_53[2]}
   );
   gpc1_1 gpc511 (
      {stage1_53[4]},
      {stage2_53[3]}
   );
   gpc1_1 gpc512 (
      {stage1_53[5]},
      {stage2_53[4]}
   );
   gpc1_1 gpc513 (
      {stage1_53[6]},
      {stage2_53[5]}
   );
   gpc1_1 gpc514 (
      {stage1_54[2]},
      {stage2_54[2]}
   );
   gpc1_1 gpc515 (
      {stage1_54[3]},
      {stage2_54[3]}
   );
   gpc1_1 gpc516 (
      {stage1_54[4]},
      {stage2_54[4]}
   );
   gpc1_1 gpc517 (
      {stage1_56[1]},
      {stage2_56[1]}
   );
   gpc1_1 gpc518 (
      {stage1_56[2]},
      {stage2_56[2]}
   );
   gpc1_1 gpc519 (
      {stage1_57[0]},
      {stage2_57[1]}
   );
   gpc1_1 gpc520 (
      {stage1_57[1]},
      {stage2_57[2]}
   );
   gpc1_1 gpc521 (
      {stage1_58[0]},
      {stage2_58[0]}
   );
   gpc1325_5 gpc522 (
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4]},
      {stage2_7[0], 1'b0},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[0]}
   );
   gpc615_5 gpc523 (
      {stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_9[1]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[1],stage3_8[1]}
   );
   gpc615_5 gpc524 (
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], 1'b0},
      {stage2_18[0]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[0],stage3_17[0]}
   );
   gpc623_5 gpc525 (
      {stage2_18[1], stage2_18[2], stage2_18[3]},
      {stage2_19[6], 1'b0},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[1],stage3_20[1],stage3_19[1],stage3_18[1]}
   );
   gpc606_5 gpc526 (
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[0],stage3_22[1],stage3_21[2],stage3_20[2]}
   );
   gpc2063_5 gpc527 (
      {stage2_24[0], stage2_24[1], stage2_24[2]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage2_27[0], stage2_27[1]},
      {stage3_28[0],stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[1]}
   );
   gpc606_5 gpc528 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[1]}
   );
   gpc135_4 gpc529 (
      {stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5], 1'b0},
      {stage2_28[6], stage2_28[7], stage2_28[8]},
      {stage2_29[0]},
      {stage3_30[1],stage3_29[1],stage3_28[2],stage3_27[2]}
   );
   gpc2206_5 gpc530 (
      {stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5], 1'b0},
      {stage2_31[0], stage2_31[1]},
      {stage2_32[0], stage2_32[1]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[2],stage3_29[2]}
   );
   gpc615_5 gpc531 (
      {stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5], stage2_31[6]},
      {stage2_32[2]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[1],stage3_32[1],stage3_31[1]}
   );
   gpc615_5 gpc532 (
      {stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage2_32[3]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[1],stage3_33[2],stage3_32[2],stage3_31[2]}
   );
   gpc425_5 gpc533 (
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4]},
      {stage2_35[0], stage2_35[1]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3]},
      {stage3_38[0],stage3_37[0],stage3_36[0],stage3_35[2],stage3_34[2]}
   );
   gpc606_5 gpc534 (
      {stage2_36[4], stage2_36[5], stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], 1'b0},
      {stage3_40[0],stage3_39[0],stage3_38[1],stage3_37[1],stage3_36[1]}
   );
   gpc615_5 gpc535 (
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4]},
      {1'b0},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], 1'b0},
      {stage3_41[0],stage3_40[1],stage3_39[1],stage3_38[2],stage3_37[2]}
   );
   gpc207_4 gpc536 (
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5], stage2_40[6]},
      {stage2_42[0], stage2_42[1]},
      {stage3_43[0],stage3_42[0],stage3_41[1],stage3_40[2]}
   );
   gpc615_5 gpc537 (
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4]},
      {stage2_42[2]},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[0],stage3_43[1],stage3_42[1],stage3_41[2]}
   );
   gpc615_5 gpc538 (
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4]},
      {stage2_45[0]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[0],stage3_46[0],stage3_45[1],stage3_44[1]}
   );
   gpc606_5 gpc539 (
      {stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5], stage2_45[6]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[1],stage3_47[1],stage3_46[1],stage3_45[2]}
   );
   gpc606_5 gpc540 (
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[0],stage3_50[0],stage3_49[1],stage3_48[2]}
   );
   gpc606_5 gpc541 (
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], 1'b0},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[0],stage3_52[1],stage3_51[1]}
   );
   gpc1_1 gpc542 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc543 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc544 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc545 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc546 (
      {stage2_3[0]},
      {stage3_3[0]}
   );
   gpc1_1 gpc547 (
      {stage2_3[1]},
      {stage3_3[1]}
   );
   gpc1_1 gpc548 (
      {stage2_4[0]},
      {stage3_4[0]}
   );
   gpc1_1 gpc549 (
      {stage2_4[1]},
      {stage3_4[1]}
   );
   gpc1_1 gpc550 (
      {stage2_5[0]},
      {stage3_5[0]}
   );
   gpc1_1 gpc551 (
      {stage2_5[1]},
      {stage3_5[1]}
   );
   gpc1_1 gpc552 (
      {stage2_6[5]},
      {stage3_6[1]}
   );
   gpc1_1 gpc553 (
      {stage2_9[2]},
      {stage3_9[2]}
   );
   gpc1_1 gpc554 (
      {stage2_9[3]},
      {stage3_9[3]}
   );
   gpc1_1 gpc555 (
      {stage2_9[4]},
      {stage3_9[4]}
   );
   gpc1_1 gpc556 (
      {stage2_9[5]},
      {stage3_9[5]}
   );
   gpc1_1 gpc557 (
      {stage2_9[6]},
      {stage3_9[6]}
   );
   gpc1_1 gpc558 (
      {stage2_11[0]},
      {stage3_11[1]}
   );
   gpc1_1 gpc559 (
      {stage2_11[1]},
      {stage3_11[2]}
   );
   gpc1_1 gpc560 (
      {stage2_11[2]},
      {stage3_11[3]}
   );
   gpc1_1 gpc561 (
      {stage2_11[3]},
      {stage3_11[4]}
   );
   gpc1_1 gpc562 (
      {stage2_11[4]},
      {stage3_11[5]}
   );
   gpc1_1 gpc563 (
      {stage2_11[5]},
      {stage3_11[6]}
   );
   gpc1_1 gpc564 (
      {stage2_12[0]},
      {stage3_12[1]}
   );
   gpc1_1 gpc565 (
      {stage2_13[0]},
      {stage3_13[0]}
   );
   gpc1_1 gpc566 (
      {stage2_13[1]},
      {stage3_13[1]}
   );
   gpc1_1 gpc567 (
      {stage2_14[0]},
      {stage3_14[0]}
   );
   gpc1_1 gpc568 (
      {stage2_14[1]},
      {stage3_14[1]}
   );
   gpc1_1 gpc569 (
      {stage2_14[2]},
      {stage3_14[2]}
   );
   gpc1_1 gpc570 (
      {stage2_15[0]},
      {stage3_15[0]}
   );
   gpc1_1 gpc571 (
      {stage2_15[1]},
      {stage3_15[1]}
   );
   gpc1_1 gpc572 (
      {stage2_16[0]},
      {stage3_16[0]}
   );
   gpc1_1 gpc573 (
      {stage2_16[1]},
      {stage3_16[1]}
   );
   gpc1_1 gpc574 (
      {stage2_16[2]},
      {stage3_16[2]}
   );
   gpc1_1 gpc575 (
      {stage2_16[3]},
      {stage3_16[3]}
   );
   gpc1_1 gpc576 (
      {stage2_16[4]},
      {stage3_16[4]}
   );
   gpc1_1 gpc577 (
      {stage2_18[4]},
      {stage3_18[2]}
   );
   gpc1_1 gpc578 (
      {stage2_18[5]},
      {stage3_18[3]}
   );
   gpc1_1 gpc579 (
      {stage2_18[6]},
      {stage3_18[4]}
   );
   gpc1_1 gpc580 (
      {stage2_20[12]},
      {stage3_20[3]}
   );
   gpc1_1 gpc581 (
      {stage2_20[13]},
      {stage3_20[4]}
   );
   gpc1_1 gpc582 (
      {stage2_20[14]},
      {stage3_20[5]}
   );
   gpc1_1 gpc583 (
      {stage2_20[15]},
      {stage3_20[6]}
   );
   gpc1_1 gpc584 (
      {stage2_21[0]},
      {stage3_21[3]}
   );
   gpc1_1 gpc585 (
      {stage2_21[1]},
      {stage3_21[4]}
   );
   gpc1_1 gpc586 (
      {stage2_21[2]},
      {stage3_21[5]}
   );
   gpc1_1 gpc587 (
      {stage2_23[0]},
      {stage3_23[1]}
   );
   gpc1_1 gpc588 (
      {stage2_23[1]},
      {stage3_23[2]}
   );
   gpc1_1 gpc589 (
      {stage2_23[2]},
      {stage3_23[3]}
   );
   gpc1_1 gpc590 (
      {stage2_23[3]},
      {stage3_23[4]}
   );
   gpc1_1 gpc591 (
      {stage2_23[4]},
      {stage3_23[5]}
   );
   gpc1_1 gpc592 (
      {stage2_23[5]},
      {stage3_23[6]}
   );
   gpc1_1 gpc593 (
      {stage2_24[3]},
      {stage3_24[2]}
   );
   gpc1_1 gpc594 (
      {stage2_24[4]},
      {stage3_24[3]}
   );
   gpc1_1 gpc595 (
      {stage2_30[0]},
      {stage3_30[3]}
   );
   gpc1_1 gpc596 (
      {stage2_30[1]},
      {stage3_30[4]}
   );
   gpc1_1 gpc597 (
      {stage2_30[2]},
      {stage3_30[5]}
   );
   gpc1_1 gpc598 (
      {stage2_30[3]},
      {stage3_30[6]}
   );
   gpc1_1 gpc599 (
      {stage2_32[4]},
      {stage3_32[3]}
   );
   gpc1_1 gpc600 (
      {stage2_32[5]},
      {stage3_32[4]}
   );
   gpc1_1 gpc601 (
      {stage2_33[12]},
      {stage3_33[3]}
   );
   gpc1_1 gpc602 (
      {stage2_35[2]},
      {stage3_35[3]}
   );
   gpc1_1 gpc603 (
      {stage2_35[3]},
      {stage3_35[4]}
   );
   gpc1_1 gpc604 (
      {stage2_35[4]},
      {stage3_35[5]}
   );
   gpc1_1 gpc605 (
      {stage2_37[5]},
      {stage3_37[3]}
   );
   gpc1_1 gpc606 (
      {stage2_37[6]},
      {stage3_37[4]}
   );
   gpc1_1 gpc607 (
      {stage2_41[5]},
      {stage3_41[3]}
   );
   gpc1_1 gpc608 (
      {stage2_41[6]},
      {stage3_41[4]}
   );
   gpc1_1 gpc609 (
      {stage2_43[6]},
      {stage3_43[2]}
   );
   gpc1_1 gpc610 (
      {stage2_43[7]},
      {stage3_43[3]}
   );
   gpc1_1 gpc611 (
      {stage2_43[8]},
      {stage3_43[4]}
   );
   gpc1_1 gpc612 (
      {stage2_43[9]},
      {stage3_43[5]}
   );
   gpc1_1 gpc613 (
      {stage2_44[5]},
      {stage3_44[2]}
   );
   gpc1_1 gpc614 (
      {stage2_46[6]},
      {stage3_46[2]}
   );
   gpc1_1 gpc615 (
      {stage2_46[7]},
      {stage3_46[3]}
   );
   gpc1_1 gpc616 (
      {stage2_48[6]},
      {stage3_48[3]}
   );
   gpc1_1 gpc617 (
      {stage2_48[7]},
      {stage3_48[4]}
   );
   gpc1_1 gpc618 (
      {stage2_48[8]},
      {stage3_48[5]}
   );
   gpc1_1 gpc619 (
      {stage2_49[0]},
      {stage3_49[2]}
   );
   gpc1_1 gpc620 (
      {stage2_49[1]},
      {stage3_49[3]}
   );
   gpc1_1 gpc621 (
      {stage2_49[2]},
      {stage3_49[4]}
   );
   gpc1_1 gpc622 (
      {stage2_52[0]},
      {stage3_52[2]}
   );
   gpc1_1 gpc623 (
      {stage2_52[1]},
      {stage3_52[3]}
   );
   gpc1_1 gpc624 (
      {stage2_52[2]},
      {stage3_52[4]}
   );
   gpc1_1 gpc625 (
      {stage2_54[0]},
      {stage3_54[1]}
   );
   gpc1_1 gpc626 (
      {stage2_54[1]},
      {stage3_54[2]}
   );
   gpc1_1 gpc627 (
      {stage2_54[2]},
      {stage3_54[3]}
   );
   gpc1_1 gpc628 (
      {stage2_54[3]},
      {stage3_54[4]}
   );
   gpc1_1 gpc629 (
      {stage2_54[4]},
      {stage3_54[5]}
   );
   gpc1_1 gpc630 (
      {stage2_55[0]},
      {stage3_55[1]}
   );
   gpc1_1 gpc631 (
      {stage2_56[0]},
      {stage3_56[0]}
   );
   gpc1_1 gpc632 (
      {stage2_56[1]},
      {stage3_56[1]}
   );
   gpc1_1 gpc633 (
      {stage2_56[2]},
      {stage3_56[2]}
   );
   gpc1_1 gpc634 (
      {stage2_57[0]},
      {stage3_57[0]}
   );
   gpc1_1 gpc635 (
      {stage2_57[1]},
      {stage3_57[1]}
   );
   gpc1_1 gpc636 (
      {stage2_57[2]},
      {stage3_57[2]}
   );
   gpc1_1 gpc637 (
      {stage2_58[0]},
      {stage3_58[0]}
   );
   gpc1261_5 gpc638 (
      {stage3_8[0]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_10[0], stage3_10[1]},
      {stage3_11[0]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[0],stage4_8[0]}
   );
   gpc126_4 gpc639 (
      {stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5], stage3_11[6]},
      {stage3_12[0], stage3_12[1]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[1]}
   );
   gpc615_5 gpc640 (
      {stage3_14[0], stage3_14[1], stage3_14[2], 1'b0, 1'b0},
      {stage3_15[0]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], 1'b0},
      {stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[0],stage4_14[1]}
   );
   gpc615_5 gpc641 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4]},
      {stage3_19[0]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[1]}
   );
   gpc2126_5 gpc642 (
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage3_22[0], stage3_22[1]},
      {stage3_23[0]},
      {stage3_24[0], stage3_24[1]},
      {stage4_25[0],stage4_24[0],stage4_23[0],stage4_22[1],stage4_21[1]}
   );
   gpc2126_5 gpc643 (
      {stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[2], stage3_24[3]},
      {stage3_25[0]},
      {stage3_26[0], stage3_26[1]},
      {stage4_27[0],stage4_26[0],stage4_25[1],stage4_24[1],stage4_23[1]}
   );
   gpc3023_5 gpc644 (
      {stage3_27[0], stage3_27[1], stage3_27[2]},
      {stage3_28[0], stage3_28[1]},
      {stage3_30[0], stage3_30[1], stage3_30[2]},
      {stage4_31[0],stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1]}
   );
   gpc1343_5 gpc645 (
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6]},
      {stage3_31[0], stage3_31[1], stage3_31[2]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[1]}
   );
   gpc44_4 gpc646 (
      {stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3]},
      {stage4_35[0],stage4_34[0],stage4_33[1],stage4_32[1]}
   );
   gpc1163_5 gpc647 (
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage3_36[0]},
      {stage3_37[0]},
      {stage4_38[0],stage4_37[0],stage4_36[0],stage4_35[1],stage4_34[1]}
   );
   gpc2135_5 gpc648 (
      {stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], 1'b0},
      {stage3_38[0], stage3_38[1], stage3_38[2]},
      {stage3_39[0]},
      {stage3_40[0], stage3_40[1]},
      {stage4_41[0],stage4_40[0],stage4_39[0],stage4_38[1],stage4_37[1]}
   );
   gpc615_5 gpc649 (
      {stage3_41[0], stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4]},
      {stage3_42[0]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[0],stage4_41[1]}
   );
   gpc1334_5 gpc650 (
      {stage3_44[0], stage3_44[1], stage3_44[2], 1'b0},
      {stage3_45[0], stage3_45[1], stage3_45[2]},
      {stage3_46[0], stage3_46[1], stage3_46[2]},
      {stage3_47[0]},
      {stage4_48[0],stage4_47[0],stage4_46[0],stage4_45[1],stage4_44[1]}
   );
   gpc615_5 gpc651 (
      {stage3_46[3], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_47[1]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[1],stage4_47[1],stage4_46[1]}
   );
   gpc126_4 gpc652 (
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], 1'b0},
      {stage3_50[0], 1'b0},
      {stage3_51[0]},
      {stage4_52[0],stage4_51[0],stage4_50[1],stage4_49[1]}
   );
   gpc606_5 gpc653 (
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], 1'b0},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[0],stage4_54[0],stage4_53[0],stage4_52[1]}
   );
   gpc1244_5 gpc654 (
      {stage3_55[0], stage3_55[1], 1'b0, 1'b0},
      {stage3_56[0], stage3_56[1], stage3_56[2], 1'b0},
      {stage3_57[0], stage3_57[1]},
      {stage3_58[0]},
      {stage4_59[0],stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[1]}
   );
   gpc1_1 gpc655 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc656 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc657 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc658 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc659 (
      {stage3_3[0]},
      {stage4_3[0]}
   );
   gpc1_1 gpc660 (
      {stage3_3[1]},
      {stage4_3[1]}
   );
   gpc1_1 gpc661 (
      {stage3_4[0]},
      {stage4_4[0]}
   );
   gpc1_1 gpc662 (
      {stage3_4[1]},
      {stage4_4[1]}
   );
   gpc1_1 gpc663 (
      {stage3_5[0]},
      {stage4_5[0]}
   );
   gpc1_1 gpc664 (
      {stage3_5[1]},
      {stage4_5[1]}
   );
   gpc1_1 gpc665 (
      {stage3_6[0]},
      {stage4_6[0]}
   );
   gpc1_1 gpc666 (
      {stage3_6[1]},
      {stage4_6[1]}
   );
   gpc1_1 gpc667 (
      {stage3_7[0]},
      {stage4_7[0]}
   );
   gpc1_1 gpc668 (
      {stage3_8[1]},
      {stage4_8[1]}
   );
   gpc1_1 gpc669 (
      {stage3_9[6]},
      {stage4_9[1]}
   );
   gpc1_1 gpc670 (
      {stage3_13[1]},
      {stage4_13[1]}
   );
   gpc1_1 gpc671 (
      {stage3_15[1]},
      {stage4_15[1]}
   );
   gpc1_1 gpc672 (
      {stage3_17[0]},
      {stage4_17[1]}
   );
   gpc1_1 gpc673 (
      {stage3_19[1]},
      {stage4_19[1]}
   );
   gpc1_1 gpc674 (
      {stage3_20[6]},
      {stage4_20[1]}
   );
   gpc1_1 gpc675 (
      {stage3_28[2]},
      {stage4_28[1]}
   );
   gpc1_1 gpc676 (
      {stage3_36[1]},
      {stage4_36[1]}
   );
   gpc1_1 gpc677 (
      {stage3_39[1]},
      {stage4_39[1]}
   );
   gpc1_1 gpc678 (
      {stage3_40[2]},
      {stage4_40[1]}
   );
   gpc1_1 gpc679 (
      {stage3_42[1]},
      {stage4_42[1]}
   );
   gpc1_1 gpc680 (
      {stage3_51[1]},
      {stage4_51[1]}
   );
   gpc1_1 gpc681 (
      {stage3_53[0]},
      {stage4_53[1]}
   );
   gpc1_1 gpc682 (
      {stage3_57[2]},
      {stage4_57[1]}
   );
endmodule
module cascade_fa_60(input [1:0] src0, input [1:0] src1, input [1:0] src2, input [1:0] src3, input [1:0] src4, input [1:0] src5, input [1:0] src6, input [1:0] src7, input [1:0] src8, input [1:0] src9, input [1:0] src10, input [1:0] src11, input [1:0] src12, input [1:0] src13, input [1:0] src14, input [1:0] src15, input [1:0] src16, input [1:0] src17, input [1:0] src18, input [1:0] src19, input [1:0] src20, input [1:0] src21, input [1:0] src22, input [1:0] src23, input [1:0] src24, input [1:0] src25, input [1:0] src26, input [1:0] src27, input [1:0] src28, input [1:0] src29, input [1:0] src30, input [1:0] src31, input [1:0] src32, input [1:0] src33, input [1:0] src34, input [1:0] src35, input [1:0] src36, input [1:0] src37, input [1:0] src38, input [1:0] src39, input [1:0] src40, input [1:0] src41, input [1:0] src42, input [1:0] src43, input [1:0] src44, input [1:0] src45, input [1:0] src46, input [1:0] src47, input [1:0] src48, input [1:0] src49, input [1:0] src50, input [1:0] src51, input [1:0] src52, input [1:0] src53, input [1:0] src54, input [1:0] src55, input [1:0] src56, input [1:0] src57, input [1:0] src58, input [1:0] src59, output [60:0] dst);
    wire [59:0] gene;
    wire [59:0] prop;
    wire [59:0] out;
    wire [59:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene0(
        .O(gene[0]),
        .I0(src0[0]),
        .I1(src0[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop0(
        .O(prop[0]),
        .I0(src0[0]),
        .I1(src0[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene1(
        .O(gene[1]),
        .I0(src1[0]),
        .I1(src1[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop1(
        .O(prop[1]),
        .I0(src1[0]),
        .I1(src1[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene2(
        .O(gene[2]),
        .I0(src2[0]),
        .I1(src2[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop2(
        .O(prop[2]),
        .I0(src2[0]),
        .I1(src2[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene3(
        .O(gene[3]),
        .I0(src3[0]),
        .I1(src3[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop3(
        .O(prop[3]),
        .I0(src3[0]),
        .I1(src3[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene4(
        .O(gene[4]),
        .I0(src4[0]),
        .I1(src4[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop4(
        .O(prop[4]),
        .I0(src4[0]),
        .I1(src4[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene5(
        .O(gene[5]),
        .I0(src5[0]),
        .I1(src5[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop5(
        .O(prop[5]),
        .I0(src5[0]),
        .I1(src5[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene6(
        .O(gene[6]),
        .I0(src6[0]),
        .I1(src6[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop6(
        .O(prop[6]),
        .I0(src6[0]),
        .I1(src6[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene7(
        .O(gene[7]),
        .I0(src7[0]),
        .I1(src7[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop7(
        .O(prop[7]),
        .I0(src7[0]),
        .I1(src7[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene8(
        .O(gene[8]),
        .I0(src8[0]),
        .I1(src8[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop8(
        .O(prop[8]),
        .I0(src8[0]),
        .I1(src8[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene9(
        .O(gene[9]),
        .I0(src9[0]),
        .I1(src9[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop9(
        .O(prop[9]),
        .I0(src9[0]),
        .I1(src9[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene10(
        .O(gene[10]),
        .I0(src10[0]),
        .I1(src10[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop10(
        .O(prop[10]),
        .I0(src10[0]),
        .I1(src10[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene11(
        .O(gene[11]),
        .I0(src11[0]),
        .I1(src11[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop11(
        .O(prop[11]),
        .I0(src11[0]),
        .I1(src11[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene12(
        .O(gene[12]),
        .I0(src12[0]),
        .I1(src12[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop12(
        .O(prop[12]),
        .I0(src12[0]),
        .I1(src12[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene13(
        .O(gene[13]),
        .I0(src13[0]),
        .I1(src13[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop13(
        .O(prop[13]),
        .I0(src13[0]),
        .I1(src13[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene14(
        .O(gene[14]),
        .I0(src14[0]),
        .I1(src14[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop14(
        .O(prop[14]),
        .I0(src14[0]),
        .I1(src14[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene15(
        .O(gene[15]),
        .I0(src15[0]),
        .I1(src15[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop15(
        .O(prop[15]),
        .I0(src15[0]),
        .I1(src15[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene16(
        .O(gene[16]),
        .I0(src16[0]),
        .I1(src16[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop16(
        .O(prop[16]),
        .I0(src16[0]),
        .I1(src16[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene17(
        .O(gene[17]),
        .I0(src17[0]),
        .I1(src17[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop17(
        .O(prop[17]),
        .I0(src17[0]),
        .I1(src17[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene18(
        .O(gene[18]),
        .I0(src18[0]),
        .I1(src18[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop18(
        .O(prop[18]),
        .I0(src18[0]),
        .I1(src18[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene19(
        .O(gene[19]),
        .I0(src19[0]),
        .I1(src19[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop19(
        .O(prop[19]),
        .I0(src19[0]),
        .I1(src19[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene20(
        .O(gene[20]),
        .I0(src20[0]),
        .I1(src20[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop20(
        .O(prop[20]),
        .I0(src20[0]),
        .I1(src20[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene21(
        .O(gene[21]),
        .I0(src21[0]),
        .I1(src21[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop21(
        .O(prop[21]),
        .I0(src21[0]),
        .I1(src21[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene22(
        .O(gene[22]),
        .I0(src22[0]),
        .I1(src22[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop22(
        .O(prop[22]),
        .I0(src22[0]),
        .I1(src22[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene23(
        .O(gene[23]),
        .I0(src23[0]),
        .I1(src23[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop23(
        .O(prop[23]),
        .I0(src23[0]),
        .I1(src23[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene24(
        .O(gene[24]),
        .I0(src24[0]),
        .I1(src24[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop24(
        .O(prop[24]),
        .I0(src24[0]),
        .I1(src24[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene25(
        .O(gene[25]),
        .I0(src25[0]),
        .I1(src25[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop25(
        .O(prop[25]),
        .I0(src25[0]),
        .I1(src25[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene26(
        .O(gene[26]),
        .I0(src26[0]),
        .I1(src26[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop26(
        .O(prop[26]),
        .I0(src26[0]),
        .I1(src26[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene27(
        .O(gene[27]),
        .I0(src27[0]),
        .I1(src27[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop27(
        .O(prop[27]),
        .I0(src27[0]),
        .I1(src27[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene28(
        .O(gene[28]),
        .I0(src28[0]),
        .I1(src28[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop28(
        .O(prop[28]),
        .I0(src28[0]),
        .I1(src28[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene29(
        .O(gene[29]),
        .I0(src29[0]),
        .I1(src29[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop29(
        .O(prop[29]),
        .I0(src29[0]),
        .I1(src29[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene30(
        .O(gene[30]),
        .I0(src30[0]),
        .I1(src30[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop30(
        .O(prop[30]),
        .I0(src30[0]),
        .I1(src30[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene31(
        .O(gene[31]),
        .I0(src31[0]),
        .I1(src31[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop31(
        .O(prop[31]),
        .I0(src31[0]),
        .I1(src31[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene32(
        .O(gene[32]),
        .I0(src32[0]),
        .I1(src32[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop32(
        .O(prop[32]),
        .I0(src32[0]),
        .I1(src32[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene33(
        .O(gene[33]),
        .I0(src33[0]),
        .I1(src33[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop33(
        .O(prop[33]),
        .I0(src33[0]),
        .I1(src33[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene34(
        .O(gene[34]),
        .I0(src34[0]),
        .I1(src34[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop34(
        .O(prop[34]),
        .I0(src34[0]),
        .I1(src34[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene35(
        .O(gene[35]),
        .I0(src35[0]),
        .I1(src35[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop35(
        .O(prop[35]),
        .I0(src35[0]),
        .I1(src35[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene36(
        .O(gene[36]),
        .I0(src36[0]),
        .I1(src36[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop36(
        .O(prop[36]),
        .I0(src36[0]),
        .I1(src36[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene37(
        .O(gene[37]),
        .I0(src37[0]),
        .I1(src37[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop37(
        .O(prop[37]),
        .I0(src37[0]),
        .I1(src37[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene38(
        .O(gene[38]),
        .I0(src38[0]),
        .I1(src38[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop38(
        .O(prop[38]),
        .I0(src38[0]),
        .I1(src38[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene39(
        .O(gene[39]),
        .I0(src39[0]),
        .I1(src39[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop39(
        .O(prop[39]),
        .I0(src39[0]),
        .I1(src39[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene40(
        .O(gene[40]),
        .I0(src40[0]),
        .I1(src40[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop40(
        .O(prop[40]),
        .I0(src40[0]),
        .I1(src40[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene41(
        .O(gene[41]),
        .I0(src41[0]),
        .I1(src41[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop41(
        .O(prop[41]),
        .I0(src41[0]),
        .I1(src41[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene42(
        .O(gene[42]),
        .I0(src42[0]),
        .I1(src42[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop42(
        .O(prop[42]),
        .I0(src42[0]),
        .I1(src42[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene43(
        .O(gene[43]),
        .I0(src43[0]),
        .I1(src43[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop43(
        .O(prop[43]),
        .I0(src43[0]),
        .I1(src43[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene44(
        .O(gene[44]),
        .I0(src44[0]),
        .I1(src44[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop44(
        .O(prop[44]),
        .I0(src44[0]),
        .I1(src44[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene45(
        .O(gene[45]),
        .I0(src45[0]),
        .I1(src45[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop45(
        .O(prop[45]),
        .I0(src45[0]),
        .I1(src45[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene46(
        .O(gene[46]),
        .I0(src46[0]),
        .I1(src46[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop46(
        .O(prop[46]),
        .I0(src46[0]),
        .I1(src46[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene47(
        .O(gene[47]),
        .I0(src47[0]),
        .I1(src47[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop47(
        .O(prop[47]),
        .I0(src47[0]),
        .I1(src47[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene48(
        .O(gene[48]),
        .I0(src48[0]),
        .I1(src48[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop48(
        .O(prop[48]),
        .I0(src48[0]),
        .I1(src48[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene49(
        .O(gene[49]),
        .I0(src49[0]),
        .I1(src49[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop49(
        .O(prop[49]),
        .I0(src49[0]),
        .I1(src49[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene50(
        .O(gene[50]),
        .I0(src50[0]),
        .I1(src50[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop50(
        .O(prop[50]),
        .I0(src50[0]),
        .I1(src50[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene51(
        .O(gene[51]),
        .I0(src51[0]),
        .I1(src51[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop51(
        .O(prop[51]),
        .I0(src51[0]),
        .I1(src51[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene52(
        .O(gene[52]),
        .I0(src52[0]),
        .I1(src52[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop52(
        .O(prop[52]),
        .I0(src52[0]),
        .I1(src52[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene53(
        .O(gene[53]),
        .I0(src53[0]),
        .I1(src53[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop53(
        .O(prop[53]),
        .I0(src53[0]),
        .I1(src53[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene54(
        .O(gene[54]),
        .I0(src54[0]),
        .I1(src54[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop54(
        .O(prop[54]),
        .I0(src54[0]),
        .I1(src54[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene55(
        .O(gene[55]),
        .I0(src55[0]),
        .I1(src55[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop55(
        .O(prop[55]),
        .I0(src55[0]),
        .I1(src55[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene56(
        .O(gene[56]),
        .I0(src56[0]),
        .I1(src56[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop56(
        .O(prop[56]),
        .I0(src56[0]),
        .I1(src56[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene57(
        .O(gene[57]),
        .I0(src57[0]),
        .I1(src57[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop57(
        .O(prop[57]),
        .I0(src57[0]),
        .I1(src57[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene58(
        .O(gene[58]),
        .I0(src58[0]),
        .I1(src58[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop58(
        .O(prop[58]),
        .I0(src58[0]),
        .I1(src58[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene59(
        .O(gene[59]),
        .I0(src59[0]),
        .I1(src59[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop59(
        .O(prop[59]),
        .I0(src59[0]),
        .I1(src59[1])
    );
    CARRY4 carry4_inst0(
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CYINIT(1'h0),
        .CI(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_inst1(
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CYINIT(1'h0),
        .CI(carryout[3]),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_inst2(
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CYINIT(1'h0),
        .CI(carryout[7]),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_inst3(
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CYINIT(1'h0),
        .CI(carryout[11]),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_inst4(
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CYINIT(1'h0),
        .CI(carryout[15]),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_inst5(
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CYINIT(1'h0),
        .CI(carryout[19]),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_inst6(
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CYINIT(1'h0),
        .CI(carryout[23]),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_inst7(
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CYINIT(1'h0),
        .CI(carryout[27]),
        .DI(gene[31:28]),
        .S(prop[31:28])
    );
    CARRY4 carry4_inst8(
        .CO(carryout[35:32]),
        .O(out[35:32]),
        .CYINIT(1'h0),
        .CI(carryout[31]),
        .DI(gene[35:32]),
        .S(prop[35:32])
    );
    CARRY4 carry4_inst9(
        .CO(carryout[39:36]),
        .O(out[39:36]),
        .CYINIT(1'h0),
        .CI(carryout[35]),
        .DI(gene[39:36]),
        .S(prop[39:36])
    );
    CARRY4 carry4_inst10(
        .CO(carryout[43:40]),
        .O(out[43:40]),
        .CYINIT(1'h0),
        .CI(carryout[39]),
        .DI(gene[43:40]),
        .S(prop[43:40])
    );
    CARRY4 carry4_inst11(
        .CO(carryout[47:44]),
        .O(out[47:44]),
        .CYINIT(1'h0),
        .CI(carryout[43]),
        .DI(gene[47:44]),
        .S(prop[47:44])
    );
    CARRY4 carry4_inst12(
        .CO(carryout[51:48]),
        .O(out[51:48]),
        .CYINIT(1'h0),
        .CI(carryout[47]),
        .DI(gene[51:48]),
        .S(prop[51:48])
    );
    CARRY4 carry4_inst13(
        .CO(carryout[55:52]),
        .O(out[55:52]),
        .CYINIT(1'h0),
        .CI(carryout[51]),
        .DI(gene[55:52]),
        .S(prop[55:52])
    );
    CARRY4 carry4_inst14(
        .CO(carryout[59:56]),
        .O(out[59:56]),
        .CYINIT(1'h0),
        .CI(carryout[55]),
        .DI(gene[59:56]),
        .S(prop[59:56])
    );
    assign dst = {carryout[59], out[59], out[58], out[57], out[56], out[55], out[54], out[53], out[52], out[51], out[50], out[49], out[48], out[47], out[46], out[45], out[44], out[43], out[42], out[41], out[40], out[39], out[38], out[37], out[36], out[35], out[34], out[33], out[32], out[31], out[30], out[29], out[28], out[27], out[26], out[25], out[24], out[23], out[22], out[21], out[20], out[19], out[18], out[17], out[16], out[15], out[14], out[13], out[12], out[11], out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], out[1], out[0]};
endmodule

module rowadder2_1_60_(input [59:0] src0, input [59:0] src1, output [60:0] dst0);
    cascade_fa_60 cascade_fa_60(.src0({src0[0], src1[0]}), .src1({src0[1], src1[1]}), .src2({src0[2], src1[2]}), .src3({src0[3], src1[3]}), .src4({src0[4], src1[4]}), .src5({src0[5], src1[5]}), .src6({src0[6], src1[6]}), .src7({src0[7], src1[7]}), .src8({src0[8], src1[8]}), .src9({src0[9], src1[9]}), .src10({src0[10], src1[10]}), .src11({src0[11], src1[11]}), .src12({src0[12], src1[12]}), .src13({src0[13], src1[13]}), .src14({src0[14], src1[14]}), .src15({src0[15], src1[15]}), .src16({src0[16], src1[16]}), .src17({src0[17], src1[17]}), .src18({src0[18], src1[18]}), .src19({src0[19], src1[19]}), .src20({src0[20], src1[20]}), .src21({src0[21], src1[21]}), .src22({src0[22], src1[22]}), .src23({src0[23], src1[23]}), .src24({src0[24], src1[24]}), .src25({src0[25], src1[25]}), .src26({src0[26], src1[26]}), .src27({src0[27], src1[27]}), .src28({src0[28], src1[28]}), .src29({src0[29], src1[29]}), .src30({src0[30], src1[30]}), .src31({src0[31], src1[31]}), .src32({src0[32], src1[32]}), .src33({src0[33], src1[33]}), .src34({src0[34], src1[34]}), .src35({src0[35], src1[35]}), .src36({src0[36], src1[36]}), .src37({src0[37], src1[37]}), .src38({src0[38], src1[38]}), .src39({src0[39], src1[39]}), .src40({src0[40], src1[40]}), .src41({src0[41], src1[41]}), .src42({src0[42], src1[42]}), .src43({src0[43], src1[43]}), .src44({src0[44], src1[44]}), .src45({src0[45], src1[45]}), .src46({src0[46], src1[46]}), .src47({src0[47], src1[47]}), .src48({src0[48], src1[48]}), .src49({src0[49], src1[49]}), .src50({src0[50], src1[50]}), .src51({src0[51], src1[51]}), .src52({src0[52], src1[52]}), .src53({src0[53], src1[53]}), .src54({src0[54], src1[54]}), .src55({src0[55], src1[55]}), .src56({src0[56], src1[56]}), .src57({src0[57], src1[57]}), .src58({src0[58], src1[58]}), .src59({src0[59], src1[59]}), .dst(dst0));
endmodule


module rowadder(input [1:0] src0, input [1:0] src1, input [1:0] src2, input [1:0] src3, input [1:0] src4, input [1:0] src5, input [1:0] src6, input [1:0] src7, input [1:0] src8, input [1:0] src9, input [1:0] src10, input [1:0] src11, input [1:0] src12, input [1:0] src13, input [1:0] src14, input [1:0] src15, input [1:0] src16, input [1:0] src17, input [1:0] src18, input [1:0] src19, input [1:0] src20, input [1:0] src21, input [1:0] src22, input [1:0] src23, input [1:0] src24, input [1:0] src25, input [1:0] src26, input [1:0] src27, input [1:0] src28, input [1:0] src29, input [1:0] src30, input [1:0] src31, input [1:0] src32, input [1:0] src33, input [1:0] src34, input [1:0] src35, input [1:0] src36, input [1:0] src37, input [1:0] src38, input [1:0] src39, input [1:0] src40, input [1:0] src41, input [1:0] src42, input [1:0] src43, input [1:0] src44, input [1:0] src45, input [1:0] src46, input [1:0] src47, input [1:0] src48, input [1:0] src49, input [1:0] src50, input [1:0] src51, input [1:0] src52, input [1:0] src53, input [1:0] src54, input [1:0] src55, input [1:0] src56, input [1:0] src57, input [1:0] src58, input [1:0] src59, output dst0, output dst1, output dst2, output dst3, output dst4, output dst5, output dst6, output dst7, output dst8, output dst9, output dst10, output dst11, output dst12, output dst13, output dst14, output dst15, output dst16, output dst17, output dst18, output dst19, output dst20, output dst21, output dst22, output dst23, output dst24, output dst25, output dst26, output dst27, output dst28, output dst29, output dst30, output dst31, output dst32, output dst33, output dst34, output dst35, output dst36, output dst37, output dst38, output dst39, output dst40, output dst41, output dst42, output dst43, output dst44, output dst45, output dst46, output dst47, output dst48, output dst49, output dst50, output dst51, output dst52, output dst53, output dst54, output dst55, output dst56, output dst57, output dst58, output dst59, output dst60);
    rowadder_rowwise ra(.src0({src59[0], src58[0], src57[0], src56[0], src55[0], src54[0], src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}), .src1({src59[1], src58[1], src57[1], src56[1], src55[1], src54[1], src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}), .dst0({dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0}));
endmodule
module rowadder_rowwise(input [59:0] src0, input [59:0] src1, output [60:0] dst0);
    wire [60:0] internal0;
    assign dst0 = internal0;
    rowadder2_1_60_ rowadder_0(.src0(src0), .src1(src1), .dst0(internal0));
endmodule

module compressor(input [0:0] src0, input [1:0] src1, input [2:0] src2, input [3:0] src3, input [4:0] src4, input [5:0] src5, input [6:0] src6, input [7:0] src7, input [8:0] src8, input [9:0] src9, input [10:0] src10, input [11:0] src11, input [12:0] src12, input [13:0] src13, input [14:0] src14, input [15:0] src15, input [16:0] src16, input [17:0] src17, input [18:0] src18, input [19:0] src19, input [20:0] src20, input [21:0] src21, input [22:0] src22, input [23:0] src23, input [24:0] src24, input [25:0] src25, input [26:0] src26, input [27:0] src27, input [28:0] src28, input [29:0] src29, input [28:0] src30, input [27:0] src31, input [26:0] src32, input [25:0] src33, input [24:0] src34, input [23:0] src35, input [22:0] src36, input [21:0] src37, input [20:0] src38, input [19:0] src39, input [18:0] src40, input [17:0] src41, input [16:0] src42, input [15:0] src43, input [14:0] src44, input [13:0] src45, input [12:0] src46, input [11:0] src47, input [10:0] src48, input [9:0] src49, input [8:0] src50, input [7:0] src51, input [6:0] src52, input [5:0] src53, input [4:0] src54, input [3:0] src55, input [2:0] src56, input [1:0] src57, input [0:0] src58, output dst0, output dst1, output dst2, output dst3, output dst4, output dst5, output dst6, output dst7, output dst8, output dst9, output dst10, output dst11, output dst12, output dst13, output dst14, output dst15, output dst16, output dst17, output dst18, output dst19, output dst20, output dst21, output dst22, output dst23, output dst24, output dst25, output dst26, output dst27, output dst28, output dst29, output dst30, output dst31, output dst32, output dst33, output dst34, output dst35, output dst36, output dst37, output dst38, output dst39, output dst40, output dst41, output dst42, output dst43, output dst44, output dst45, output dst46, output dst47, output dst48, output dst49, output dst50, output dst51, output dst52, output dst53, output dst54, output dst55, output dst56, output dst57, output dst58, output dst59, output dst60);
    wire [0:0] compdst0;
    wire [1:0] compdst1;
    wire [0:0] compdst2;
    wire [1:0] compdst3;
    wire [1:0] compdst4;
    wire [1:0] compdst5;
    wire [1:0] compdst6;
    wire [0:0] compdst7;
    wire [1:0] compdst8;
    wire [1:0] compdst9;
    wire [0:0] compdst10;
    wire [1:0] compdst11;
    wire [1:0] compdst12;
    wire [1:0] compdst13;
    wire [1:0] compdst14;
    wire [1:0] compdst15;
    wire [0:0] compdst16;
    wire [1:0] compdst17;
    wire [1:0] compdst18;
    wire [1:0] compdst19;
    wire [1:0] compdst20;
    wire [1:0] compdst21;
    wire [1:0] compdst22;
    wire [1:0] compdst23;
    wire [1:0] compdst24;
    wire [1:0] compdst25;
    wire [0:0] compdst26;
    wire [1:0] compdst27;
    wire [1:0] compdst28;
    wire [1:0] compdst29;
    wire [1:0] compdst30;
    wire [1:0] compdst31;
    wire [1:0] compdst32;
    wire [1:0] compdst33;
    wire [1:0] compdst34;
    wire [1:0] compdst35;
    wire [1:0] compdst36;
    wire [1:0] compdst37;
    wire [1:0] compdst38;
    wire [1:0] compdst39;
    wire [1:0] compdst40;
    wire [1:0] compdst41;
    wire [1:0] compdst42;
    wire [0:0] compdst43;
    wire [1:0] compdst44;
    wire [1:0] compdst45;
    wire [1:0] compdst46;
    wire [1:0] compdst47;
    wire [1:0] compdst48;
    wire [1:0] compdst49;
    wire [1:0] compdst50;
    wire [1:0] compdst51;
    wire [1:0] compdst52;
    wire [1:0] compdst53;
    wire [0:0] compdst54;
    wire [1:0] compdst55;
    wire [1:0] compdst56;
    wire [1:0] compdst57;
    wire [0:0] compdst58;
    wire [0:0] compdst59;
    compressor_without_rowadder comp(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .src54(src54), .src55(src55), .src56(src56), .src57(src57), .src58(src58), .dst0(compdst0), .dst1(compdst1), .dst2(compdst2), .dst3(compdst3), .dst4(compdst4), .dst5(compdst5), .dst6(compdst6), .dst7(compdst7), .dst8(compdst8), .dst9(compdst9), .dst10(compdst10), .dst11(compdst11), .dst12(compdst12), .dst13(compdst13), .dst14(compdst14), .dst15(compdst15), .dst16(compdst16), .dst17(compdst17), .dst18(compdst18), .dst19(compdst19), .dst20(compdst20), .dst21(compdst21), .dst22(compdst22), .dst23(compdst23), .dst24(compdst24), .dst25(compdst25), .dst26(compdst26), .dst27(compdst27), .dst28(compdst28), .dst29(compdst29), .dst30(compdst30), .dst31(compdst31), .dst32(compdst32), .dst33(compdst33), .dst34(compdst34), .dst35(compdst35), .dst36(compdst36), .dst37(compdst37), .dst38(compdst38), .dst39(compdst39), .dst40(compdst40), .dst41(compdst41), .dst42(compdst42), .dst43(compdst43), .dst44(compdst44), .dst45(compdst45), .dst46(compdst46), .dst47(compdst47), .dst48(compdst48), .dst49(compdst49), .dst50(compdst50), .dst51(compdst51), .dst52(compdst52), .dst53(compdst53), .dst54(compdst54), .dst55(compdst55), .dst56(compdst56), .dst57(compdst57), .dst58(compdst58), .dst59(compdst59));
    rowadder ra(.src0({1'h0, compdst0}), .src1(compdst1), .src2({1'h0, compdst2}), .src3(compdst3), .src4(compdst4), .src5(compdst5), .src6(compdst6), .src7({1'h0, compdst7}), .src8(compdst8), .src9(compdst9), .src10({1'h0, compdst10}), .src11(compdst11), .src12(compdst12), .src13(compdst13), .src14(compdst14), .src15(compdst15), .src16({1'h0, compdst16}), .src17(compdst17), .src18(compdst18), .src19(compdst19), .src20(compdst20), .src21(compdst21), .src22(compdst22), .src23(compdst23), .src24(compdst24), .src25(compdst25), .src26({1'h0, compdst26}), .src27(compdst27), .src28(compdst28), .src29(compdst29), .src30(compdst30), .src31(compdst31), .src32(compdst32), .src33(compdst33), .src34(compdst34), .src35(compdst35), .src36(compdst36), .src37(compdst37), .src38(compdst38), .src39(compdst39), .src40(compdst40), .src41(compdst41), .src42(compdst42), .src43({1'h0, compdst43}), .src44(compdst44), .src45(compdst45), .src46(compdst46), .src47(compdst47), .src48(compdst48), .src49(compdst49), .src50(compdst50), .src51(compdst51), .src52(compdst52), .src53(compdst53), .src54({1'h0, compdst54}), .src55(compdst55), .src56(compdst56), .src57(compdst57), .src58({1'h0, compdst58}), .src59({1'h0, compdst59}), .dst0(dst0), .dst1(dst1), .dst2(dst2), .dst3(dst3), .dst4(dst4), .dst5(dst5), .dst6(dst6), .dst7(dst7), .dst8(dst8), .dst9(dst9), .dst10(dst10), .dst11(dst11), .dst12(dst12), .dst13(dst13), .dst14(dst14), .dst15(dst15), .dst16(dst16), .dst17(dst17), .dst18(dst18), .dst19(dst19), .dst20(dst20), .dst21(dst21), .dst22(dst22), .dst23(dst23), .dst24(dst24), .dst25(dst25), .dst26(dst26), .dst27(dst27), .dst28(dst28), .dst29(dst29), .dst30(dst30), .dst31(dst31), .dst32(dst32), .dst33(dst33), .dst34(dst34), .dst35(dst35), .dst36(dst36), .dst37(dst37), .dst38(dst38), .dst39(dst39), .dst40(dst40), .dst41(dst41), .dst42(dst42), .dst43(dst43), .dst44(dst44), .dst45(dst45), .dst46(dst46), .dst47(dst47), .dst48(dst48), .dst49(dst49), .dst50(dst50), .dst51(dst51), .dst52(dst52), .dst53(dst53), .dst54(dst54), .dst55(dst55), .dst56(dst56), .dst57(dst57), .dst58(dst58), .dst59(dst59), .dst60(dst60));
endmodule

