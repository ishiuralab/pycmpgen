module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [19:0] src21;
    reg [18:0] src22;
    reg [17:0] src23;
    reg [16:0] src24;
    reg [15:0] src25;
    reg [14:0] src26;
    reg [13:0] src27;
    reg [12:0] src28;
    reg [11:0] src29;
    reg [10:0] src30;
    reg [9:0] src31;
    reg [8:0] src32;
    reg [7:0] src33;
    reg [6:0] src34;
    reg [5:0] src35;
    reg [4:0] src36;
    reg [3:0] src37;
    reg [2:0] src38;
    reg [1:0] src39;
    reg [0:0] src40;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [41:0] srcsum;
    wire [41:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3])<<37) + ((src38[0] + src38[1] + src38[2])<<38) + ((src39[0] + src39[1])<<39) + ((src40[0])<<40);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1495263acc0b26512d62b5ec67c7cc3c1172f4c5d08b10ec307714054a9ca072893216aa7d81368e6c26a57912acd20711c98513481596c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d0cb0c87cc0a653b6184f81f97aecdd5a8b3dfd545f5510816b3e07fa218d2a37b62bc41bdaa3e0dc6ecf05948dd0bfb467d725fd152b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11dcc6399494e3c3d70124cb6804014928566f15ddda2d2a494a3fb33d259b8dcec2abe4b630908d6a56a2f9d5b3df5ba5653f251f47f9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4a45197e0bf50965ae62cf2a230f1ba0a900510763489a03cdad04c51444d432c5439bdba78c42ce4c3bfd5f9043baa5c99b75fc50d6f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d077647e31baadf8cc3a7f9384294a15e2a7b2c17b8d963962c4a3412a23032c65fb737eeb33740c95aa8edabeb82b08b3fe1dc5dd31ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5f3b43de27b320c39e90cca9779872d9b974da2204011523d4ac556c176425eed69676c318fda61b249318ff3f3845c7a7820634b5e8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81716f0d52d0b13389ce96c392bea338a1281b19b6faeb0f778c4a2261bbf5e0807ec4330f0f6a134819b5c82e58ab30821c65fed57392;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad4057f857940d2dc3f03a576b25def6eadb4863276d810eb544e6b059757afc789d96e4f7e09a1342451af6df94da4219748303face98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b042babd122ab1e782458f16ffe4c9e877043b29a4390feb12605928ef35fda2a57d850aa9b9c7852f5d30eb65f42dfbf178756e345dec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10883a58721d3a2103dea66ba590c4f50d60bb70bbb9748e3ddafc4ba1ce629df0d6968a658e06d415f5dc512bf398bbc9b44294252c53e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae628efaf8c608acd604a324b8840d3b67ff0560742a7f366abd163fcce1b3aa485ec4f75c90902c77d48e8cb834e0a330667e2cf76d38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2978a15ec0c6adab4d60d9f7503a06b8f0e9fa5c1963d64bc3938e3e4b26b3ad563481958d7b782632c11ea3832ecd38b2f90fbcf099a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha61ffb6374e9caea3ed08058d15a86e64b4994a135f2706bc754463e1a9aef991429bff0f5e200cbed0b4b869e1cf49884124116e81910;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175547ff1029cf7e9d5dd96ac1f6a30e94595dabc4eb5d891882cab2060909327f7604358cba6768069b9371f83200819f5ba2150ec38cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58b3d21a4388aaae94535e040158f75662e30b09c08a11198602fc1025955143b277c3b6537909424772329b8f19b04b3568f03e207490;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152a82d08446be1fe93c8b253b2b957a9f0be08aa3e2a18b3b01d0a82f0367bdf0ff6ab7ceeb3f9d27ac5e171997f7800aaf5b61c99044c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he25f630d9e4fb96536ca71874f830da809f57659bad92be9c856959a6eedb686812774b29a5b87651e47ad3be83083ac0272d7d5662239;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16232cf817923ee6b1a23fd2599402123db7246063941809726734dcebf0211d058de1fae87a879fe4ecf844136bfcf9b48baa575ef6891;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179d741babf2206892250381b19e9c30c610851ee4130633fc908ccd0416835b77e4278b5f15542ca8f5690be35e912452ef78c82c97694;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1461edea203b7488f7d9cdf54bda9384605f5cb23bbc024225648539073c6421af8212a9ac884fc5a3bfc6e50893fef6a456dfca4c8f236;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e1ba990fe03074689a580d388bda4508785b43fdb787a965e65bb974cf8e6f57ea39da37852c79dad1b7199deeb4a4ef583c959ea6449;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h863e8fc65380b95d498d0036a70b2d2da5ae56e064aef912c80654ec4bde7ae5cff3e26c972802de19839442d7cd58dd88c3e72732800a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h119e55c926205707039c795027c9708441c86239433af377972b7f741a8ce6481dfa572bccc1d9ce5239b21db203bf961a2a7d321eb1160;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a8fae4ceca559d71dc264e97723297364ba838d65dcf0dbdebc44562ebf8fa56b02b1674c00efa6f410812893ae4c5534760ad9d3faa6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a13dee92d8b132d7326b0022d650ab29fe6da295f00f6906a14520b3c72f092a9ebf6f6976a2013845dcc7c873f6d0bd3e585ef1347f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb70a30acafe377968a3881f1f146b918697a8658ece176ad317a661baeff44208fb0caed2f06a5a4d0010ab52e6dc35250bd05f3d17c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49e79fa4417d2b243c0402c272cdbe27c73770b2b16b20cbd752317d8ed700fd6ef1f2ab1c95d3eefe630f847a6511e533f1ad678911f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140b0800f60edf2e49c23f898149828f4975161163701bf81f3a9fe76a4babd0616016e71f9fa7645645041814f427827561f3be9fb5114;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11206dd767666094f1a159c3f944bc963a837c27d27dd195992a3b1aac757dc8f4055527dcff4e9310e6809a2d5068bc4f70fc7fd516ac0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82de6481d724aad2b5ad291e178ff6e1efcb135c38a6ff50487535a65174d4f672c264d67eb3f98d1460ac55cf5de56fb9d0fcfb704a45;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75cd1e4dc6c28f54d386916c903ad5a528744cbb2196f618a4e4dc5cf496cf7a602c49ed048bfdb0ec665041b8555ac3b24a6101a6d585;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4aba8be95b50528d437c241ea0a77440fee8074d8035da2b296377849e1b6902dceebc0b91a449650a60311eb191d131790f4462d57c35;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57848fdd0dcf7eeccd09ea25df70f3b5ae6f49866423ee6c8a8872fa3d654dc2cf72482c37fd65bb06d7bbfced6d0a33a76cc818a168b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h48dd1a16f12357565f227b08663b3cecb5775a74fe302f6ee1127e801bdb1c260994c2e733783fd95f40aebdf6fae535d5b9d680ca4987;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130f93617dc2c1c4e38bdd9833b927b1816790944fea82e601a81ba6de0f15f9b02d780ffc875a6a6b019da05262ebdc457fdf05ad39afc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb797dadecfbf0ac32dd7036d1d1602a72389b13d7eae70d393e45d5905e4eda468380994d059e638a19932c2f486a83bab48902dd4f9f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31971fb564d2279e638a025cd0068ce4b75ad0eba70e3f46e0696c14a6d00ac745fe2d0c8373c678d5a51e4c6f04ea1026487c2a7f60f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164de9089b40d50cf4833c50bbe0f9354c7d0ffde312aee0ceca6b36f539e65b8b6eb50ec67ea0240ba73cb9572860123a5df43ec45758;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10787d55529d876766765a9acc6d4b9112cb4e0fc52edb171a646c4864b71a45d4c400e6488bec63cbb5ea5e1cc1ca6ef9e7d4a877b9d75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e783a2fb8aca21f6c4a309e6393537418a1f7773464b16c037a8cb53b7a60e243117095f7e5688932a690d1c938b7c78484f1632ab397d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb96b2979d1a5ee197406f77966af72c56cc2c2cc1d912e307c3a99027a0a868fb591a887eb5314755b5e4aa67de9ebd20b17e2c569b28c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf72f459d8f16bfb76965ed934ebd6e071c3adcc170cd5bf83a8774bc0a5a32a6f481c0c90b1b705f2e92dae2f414be19b3b99235ad43f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e26ef120f3087909e4026c9b9a9e376322d9c13d23736044fa2629a0fe794ddc7b42326f7f9235b17b7ed6d7ac54d1e64627d775e777a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f174c432f1ed1ce812b86e7098d760533a76c0b57ddc83644d291b59a4b11bcef1ff5090091d6cdf2834666f5cc16bba905065abf07a99;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b49b90dc41aea7a38a484e30b44b6f8ae5e0dcf9eee06e081674d650c80c0a294380f58b0ff02263df71a3b247b7a52547b573b088a0ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e4199c71b8caffb425298ccbb90e8211cf6283ac7e3ccc3764a6c2cddd6cf97de4b36b6e7088762289b21094ac4367b8b08414818a389;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a112a6aebcbf55d3ab84f078557d1eeaca96bb00a90bd15ef92bc763feba79eb1c27ccf3c49a3173a4ad08b0d91e3cb494199ff4bcb7c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c1d5da8258b7c9f1a744e06cbb551d63574a70bda8aa3747309dbe4e4f9494cb5c53ae9537c772606eb8661d334ed1a795947135004f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h50c72260c573d036ea19209a975e8df77ff07bb6c4282d13a626eb188c37cbb93a7599cee38a3584daa8021e88e0786b9d3d6f39f7ad41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11071056aaf7aaa3270949859715b8bd64384b463a52f95932a31de677abedcd836029d21f03b183133e974fa6314dd7e624d6e8b5e35f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h350f21bd9acc62814439cc01b2363e83a70e6f713d6c3fd8bf698918e8baa58da8f35faea83eea8789de036957b95d3cee860d04601465;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3a276ff2302d2a6c7d5d0e108250562a4e0246d5e4532c7234485a09743f3d09c9d14a5598f8d1eb3c508c9db1d25d68863b0e7299af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132a89b2412bdbf393c706948ff5b83993bd5bef2c4841d4a1ac0ad7d4cd3c7525f43a810d16d58222b73f9bcc009ddb320ede408d2699f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de499b896e385fabee54f9e3b58682020977203cb66cc7ddc2232e335a84b5180aec896154980ac26860668e37a1847e00bb698f762c2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f8314b566eacf1874b61af9d137bc628e69159dff0bfb7acd181882f48337ef7f9fc9045bddabfd2b1940b47e683d7129812b2ac50627;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1208c54256e178ac71fd05a6a45cd023a2aedba82933910e8298a54b947fbd2e31756ced33ac720ea672629de08d34079bbfb194faeb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h773de7e410af9f38640050579c9a2217af5d4b6f12381c0a1740fc43e10e484b145fdc391b8d44a6a4e01ba09499ab4f0168abb7a8dd15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h661b7ed2d2b3d4995e37c93334013c8a330f478bcf8572e4d0ec800ec6d8a8677b215f7de6b27bf706fcd2849f7d2add74b6cf23ab790a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd67d5d1fbb0d7365a36474bec2b39d5d2fd0817a4e7d0060f716755e9f111025e6c61f902e80c768b37deb8c2ece6e9bf978438b3d60d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca8ed99119bd96c8a37536e3add55105c81a538b9b62f3e2fa1e6c36fd081ba0ec475da566f21b2d52da8e53fb1ed16cee7c8a6141b76f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f6280b8497422ac07daf72d270e259e10e20e458a22b7852e82ea02f2c640bf71469ac594184e4e1ff57eb11c932b661927872e376d42;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3c5a59ce4dfa30da0366aba3bc36b142d3e0cfe72214b548e9354a5c0da907da4939d1c5012329d14e5ed3a93f23af12ad1eb1e2b2959;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e8e103aaefd5aa794c8f3359017b6cdf0021369f3629254f82ee1607d593404b6295b8becabadf3ee97b9bff27f13c8cb11d2024176c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1599364746a0ddb9def6866e3080f83ce18c47245bb1533cee8d6e6eac7cb7cb2d26ae73c1fcb995f1ec4ef34934172dc9d8e10ecd94016;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1501247364a3a53274c2395954e950ae6462566bb0057ee87f6f353cad56967318ddf46a8493c0cda9731e2641d02c682992f764b20a446;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf98602fc089f7f554579241f1cbcb93d4eacf5c204a95289358057a679f3840862f912d42cff961fef826c26040995ea1bbf8c897e178;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hccf016c005bcc7da9b0b5b99ccd27be6d31fb56234f56418a606d971a290c76863b4d196ffb1fc5c5c3774d06dff0b9e7bbc0d0817b42c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habcfd61704038f97d8f995b1b28610ccbdfffc7c627817b064798e303a2f03d9b096b27aac381a11f35e592b86e49767e78430382c6ebf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cbf3a9b38a54709bdf085382179d6f0b6e05145d9953c125666bc82518e5a22a32a72ecd10abeb0d597580f192df4303f2fcffb93c1f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h797cfd6baeefbc87b04322e3a079cbf37df0c70bdba7b073e37edfe7b5ac7f01d7a8022b5c1129a31eafb398d49d192e17238fe396d498;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23950f207d69c0dd478e0040181775ae7ccd92bac3fa9bbf2706114cb6cc57163a196f5d972455561245ff905c46ae61eb97e1a704fea8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19363875905500990e25b640c7d434a66901f749f5470f9239d7a0c06be215c78f09f09e6b72ecda2b10c6e8bbf874915f18ba382052db6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a7c5cf18b00695a31dd4b16b2063257cca67cf95d13d2b158405f9f59ad8715f2613ba7ada5b130e7ea18c34196e7c835fcf0c4980f69;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de37fc53c125c8eaa23401f4b406c57df6798ad94940cf01a1043c4761dc217e15781958723cb474636a04fa60fc63ebfaea07b3c7a04d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124ac52d5a9c06ecfae6a1f2def6b257d9ad5407c2ae4c7fff6e8bfd78b08231882ce1f772a679f7fe988c79ab57553305f79639d115f0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb6d42d034069a6c83b0bb4f35e115024dfbb53f63148757934f6a6729ec70a972b086a46aead5ee22fe27583f02cd30a583eb981846b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe34b7bcca1b84982055a380a7920043f38e4d14cd46667d5f8b8b6077c4416155f4aa9334d911aaca32702c31bc838d1e85cea124bfde;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdeb2220c21e9328c3e70c98bf644c512e06c9de88857324a86cf742f278b6de91b5736e9dd7f8e73538666d441c0e1bd91c739a0af1c2e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60756d2f7b365d505d722f2cdb8e4c0fed1d585b6143bd0d4fbf4079a8f34321f860dafc42780e5c7570718cc6f6a361a90769c59501ce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc54c4e014861e3f590c7edc5ae6d66a0a5d90028d18c67a46d467d6f435a6420369ec8b75d2c9303167789aa7ecbcae2c8105794d45622;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12fae8d7f8e289e5fbf065e3773d169d06cebfe877f17fee4219edaa000e0210d49c0d0e8be372215d59b3e9f508258ea5b5b1693cbe910;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e8f4dabcd4dff87225a14a7ff40fbef059e3d41cf4deb93ed4468990099104c94ed00640c7c0bb0513342223080174ce7560e66a5a4c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a38fbc4af3483bf2bc9f9ed6402a6d331bc4be7fa44a9fb0d1893e2608887bccaea3c6dc41daf9beb6d7b3fd80168e4a663321eb72d64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7991a36b56f6b50090caafed6225817493d90906f9e7e4b2f9de3fde3336afa003d0c06992aa76e613cc28219461dca3313f85d35a967;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd22ecac91c664179db1acc4d6ff3c7001a5e6d017e54e80dfd3bb52985e4e32912fa3c35ba6e3ca731d8e7f3ffa421972eedc6253db73c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h920a93301cacaf733287e7257acc73e0bf2aa954bc5b25e2e16f05076a7edfea3fb9dc0bad98717445710e5128580a63a0a790bd87ae0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h833818cd7b4598f0e5525cc1bdd63d3521f946e4625955e5defd13767f1b32c54780955a5dc9dd0f61b5e254eed939eeef6b27eb12cf83;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d302dee423e1e3c0075541dc0943249b0093ca11ff9b57a050da3541f076cc6c45427d22c82e8f48e1ca23b4a0125e792c29785f5fd47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191aad7bfbf99784bb005da49db92d42983de2f569923aa642e98a213538b15b917154dd7c3b0e23b84b515a7e69161a7e1c567a7b4f974;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffa6a09080bb3a90909f564f0860c968f22216d76a09ce05156f170a0f741f7215f3293b985632c284052abdfe56de13f40562c32d2785;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe1e24ae8f1165cee779cd01ba488061320392775f6115fb54917fc3d9be55acca36567ddf98f8c95b65e9be3a80d66a972b174019cd66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abf3d8116a0faafc803051b3f8331ed936d026116807ca71ecd0a7229a669cbbf57b4ac2c1ef3a8a3622574c788b72236a083b28d7e07a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ab7d5f52a11bd03acc5612bef766b69ad1cada50f579aae76d923c6070f3b503ac6a7224db348659cf466494fbe685650e1ccaee16fd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb66dbc733c9dd145bc7e9b43ad6dd0d3ca2d593883c80f0fcee51f6db74cae5cf44ab3b7a94f464ff8a859f71e1b17e265da1a0689622b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178c33a6f3c94ada53640c3caf6d8c9b3e77bfec88554fdabe0b85acac5c39ced571d25dd6680d88f00b92518ea48fb7224fc74fc88b0c7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1542544ed770d59a984851300ebd8384140f0e9a87de5d49c824bf4c98b453aa0eeb7050e154f9670d66b65a2fecd264c094ecdfcbd64b1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd322861219ec80a265854664576d7ad74aeacac982dd2e5a1028a4206effb6fa6ce57c70820bb2f9b96adfc645ff3bfaba2f35951fd95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15af855d85e5e404b46d41b649b62df1fb41721fd5afd38ecf9cbd9424e4792fc73c0bc7b5293b6132c965d5894c5281cea7bbf60158b5f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9728cf255157c6bef2c5ded00824f5eea92e42322455fc26830cb0e1ff2d1b57f124d2f85e407de75e710b70781878bfab5ad8a21f1ee7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4edd60bbce643c8213c67a6524fe82a9e22bea5bf5f42bfa7f2906f61a53b25116e85a6c06cd5f67fd190285d78d1c9cea25392a0e878c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1651915f7567ab464f0e11df960a208309e4b8c7d897481c76fc04b5f7f3cfb618e0968c30da35534f54aa9fcda1ee01241fc8db39e1603;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2bf8ac3e5145ebae8c958d51dfd2548d36675c5e7a1911696e8d7966692f34dbcc05eb03fd832458fad7bf74e276b4df9ccc50d137d7f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h795bd749377d73cadfb93c1ec5c119dcfcb1c38628a3fb8714a783f5f9e09874e90d8cb4fa68234d08c75b11bc5a026f9b1087ac433f47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bb275602eefb0c08dcffa889a36f0491fb7c53754f8f3a3c0993f4eb4b22631606f1a7941f93e0c83cf00d0accf36802bc0d2d02b8126;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea72f23421d27d8b272ec4270b5892d92acecd61e0c9c66039db4aa0ea33949fd4b053b7ffd27b1c8cc873023e73df86be7db0b5080d9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134d54a9c7bea1b915f2c17d6c021f763f715a4dacc40f4f607965bab765c293a79969005a2fe92bafdab7ace0876b2e6551ff929727285;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb853f334d428ea3b4020632234e817e5861bca6970e18f159bf69ba5c009703552082c3f06710b4b28f6cd87cfff781993126d9bcd8c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha75143b7ee78cd402b2a016261662885f3e1a925725bd853725a13604d1b27d06ff2dc43f0507982d2999e303ccdee8fb5d4efdaa2bdfe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heec4c98143be125ebb180afd44d7338d32e271a87e5cdf4a184441ded0002842b196c28f11aed9a752a6c802d0409388d4f7daa4c9bdf3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144ea775e822387ad92e9c84e700d64ab79576953ddb35f710905cdfdb499bbd26f95cb9f3e0611912c7bd3aa0ff576f48a3b73f8ba071e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4f90e454d6ddfa67dea377d4bd2da769407ca841301ba23f190cdf3ace2ddeb4fcae5eb379a73c17d323b8a125e108293b97eb34b76a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6bd029b161d9165b7f521f8ead5f0eaf9efa5a060db1cf096016ccc29fce57fc7af1f468fe068f76744125089eaece14698eebc58fc07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb67c30cca306475197240bfef2ede5c6f43a6ffcad49925eb8ea3ea29b9e548fb837570f9dac915b8883e657a2e3141ce9b6eac6b388;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f974ae990faa52601dd0cb2422f170561ba1f6f97dce7a16ecd611b1f6781d49b4fbbe4db18d3a21446d7f36fad7f361f39ca16348fec3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a9ad29ac0a01fc2414455da68d57a31f19deab860e45bdab2be3e9f6c625ded99db790b1e3d1dcef1dd2bcc521dde9975298426755e56;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd62d769c469c309013be58a63ddb35d05a6b5693a43eb649daf6539c23b88fcc000b1fc93037ca79079c8151791744b8a28dca439f654b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16379f3f74561cdfd2bc6885f6e738565d6185d726156b08ded6f104d45710e9e62841106cc4c244652ab88650a8e9a52661a10a62456f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfe512d1df5e539721de03c1dcb91227093cca54dd8e733ba2faba98c5f39b5f2352e0882dbd1ebc59698a90f9ff486f1a6a23fd3c7142;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfddcbbe3ca9d678d13c63650c005d55af3e5568c88eb40eb932772de6da319b409985bf692bda48d406acf30e209387685fe3d5f17db2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1899c2d94563903c65208f68ddd9a49ba0913319d58461640301c6683dbab7c8f320fdd16ea453083712febf5c466f10ae97207ad6341;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha87e063e9d7a66d6299e5503132f851911d7208706fb3536309c90e47b39e9bf89d86c30e500d4df4603bd17673af0c32a447a3b3925e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed213c20860bc09a1e87a16609a9acffcb6d1173ed29fc1d30d4145e9c19cb3a11a0c7c9f6e7d205fde5fd574f3e568605f0832ebf89fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1752746214ee56d50acd28333441609ae798f816ca9f6f255de93f675c621ef96147ad705b0ef99110bc07dc9c455d864513cb31e8eef74;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a6cc6c8ebbce65b7e62356fe3698cc6c1013a62c80eab36d97002939aac75b5e219ceda36c3751d9cbc4c9aa62d39ba5e5aa258e1d60d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162bc26045ece433eb83bd1753e3bd369d66d86e46fbe61ce3e73aff02c72e83a4749c754056c761321f6cb6affcf039a2cf6867fd304cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h210030bd924902cd7262cca9d347bb9da47bfcf2df77a850032ff6a91a0dca61578d532bc0505de6c73321848616b59fa03ff88abfa735;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b3efa8cd5f03a7e23cbfa3aee3fabff90a7ed7a57c1885370b62bbd4fb2b092453c52ab46c86ff1048da97f7ce0356be97dd827b72450;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129b8d585738f65e5bbae63465150f99300575ca38bf052e004c9c0dfc9d87c30ee77b45c1e1776ff35aa5e1d27365170b2e93d8fb7601;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba77df07e4e26415b483fbadce5be7d95e411cde5a81b42ed4b235187f95e8fcc1e70a4338e4e26d23dff05f252710b94bf62c953353f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a67fa98fc58ce494d30e6bfd2c319eb5faf7bb47892deb1aaa483c78082a6dc82ee3c6b7a77ddc1ac7af4f17940585cd8b1d0af23a4c7a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1805eb9f69ca2c317f2338655d880c54b84721521a5f95509f9fffdf5db80657278a5e1820556c543a66e13f1c61fa3fd204fd6180c1d7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb33db9903eb16eba196a69ec28079e3c314e22d926da5ffaa39583bd091374b6e406cd8c0c86a62be239dc9752bdd04a80a500f7b624fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3228f160af48322b3179fdf3bd68dac522471b46e5edee682ca61eb49abcc500c192aba20b207389d56d4017ed1a5ce70d698190affc9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f05cdd5bf42a5502bbb9f0b4e420ecbd101175b8e6370c8a6a98e15f1f42003b85c87367b90c5e3ed404fa5c014a0446c6074bfa1026;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0e3268e944ddc1e876829475fb7f02407b66ffe2d31e95156c55e6ec9614e006eef63e3a50e45adeb31711eb9042c5e6977c6c7ce99ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4f93f7e8a833908d677acc03876888ffba93cc9c5180859354496b394b9d96864164162daecb2c7c7a9dbe1e9f4d55c23ded9cb6190b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127f1df4ec028820416952916eba709140fff8b0ad75baecfa76e1405d19ca38d0f742a6b3a9d546fe2010b70a66d6a313cbeda5ddac12f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d8ce6aa87013d096503eff667f6721bbebd893523aa2d40a7e7e9f5e8d213ca31a14378279760bfd0714f7b8f6092cf53710a8f02667b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d58c20f7102f7636db81c07ef5f5562efe0d40708b746513ab091b5d3a789960041ba4c6c82e9b65cb513004058bd550c35259e93a454f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb89beae6dfa1fffebf4291c13752c35690dae1e48274437592dcd3fa1f275f341450af5f413c409569ca482e259d1a946619e2cd007c66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1798b3424f860e933a2a5b4df8701a42382fb534e2bdeb745e4312f5941f4627acda1230d3c1b7fa18c68c1d68185d5862876d8746261e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2913f884edf6999bcddb62402eb359278f7a2d8528869e1d64a4451fd60be52b5c14fab00ae4ea874b16e1caa18230c9745aaa2155440e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf221bae413b5d7140e4f8878158c0ff5780367c02993e8d146425e3e4b4e0107a970b0fd92ddfb83b39c7fb62a79663aeccb08aeb86579;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1c7432a331ea24d177ce5336fc93e69aa8ae0eeedab6749f411aab9599d0249085ea3baf32a924e42c2821a0fd6a36d51163a2a4f4bd5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h408e8655cff722fddc4e8909b2f1154360810b18ff154111f1a49ea580997747b184890c30243adc20a13e7476d2563ba7a54493451843;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d589edf44e400f9f578dc234acbbaaf271f4c0f92100a188a8267802fd4893b65405752ae351724a0c7f28ba95f424511d68116c0e6acc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1078f07eda4c4add63015af7f992ad52d07dbe17ca19af1f9e6f499196a6885e488f23f77204d805c471b010c5ae9c7c6624adec1cff5b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10377366e8f106cdaaacc01193c6ca095055c981a8c3361cd70d8a446f25ed4b70dc6324e400c6b9178e87d242a252e5a7c487620104f81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e48c1e9cc140087045435705560718880c94aed1408815962d44b66e0d9260ca455b1c4483753de81a8af5852844942889814ee3bdc6a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c6c7cfacd912e3edacd418af0542d2b17dd8a86d3239a16b58fceab31e8e189ebf5614b5d4f06bd7ba466ead12419fd708dd8fa870948;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec8824c513a696220d5415cf9294a92f509b3596857808ee4e8f58fbec21c331f51fa64ff3cc665e788588a6f890280ef43af0e9a8cee0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d3cfa5141a0f5a2aa730b9088eb390440818d6c39b7cbfcf97afd8e6787d9f010a6699a303065d71109018aee71bf49d419481e2228e5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53d386356d4315d9fa798bf43bb278246dd13609604fee0461338e6b8d8c71b5d1c80a51380aa9000253e3ffb0c6e8a9b549f7deebf0e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120900e621a8e848657e8799d987bd397990e3b1902464820c1f7a220f37686bed9f45060cfd317d15da0227ac52aad81252a449e1fff86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b78fa23f5fb7f6b0acff2d6b0a70dac22f87bc0ceea200b27915b4f54333f6733156a7676ed1cbdd0a4392a8c214a1ad87e795c162db5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5803ba199c8d0a042e986024613b25c05caee4e7a5e48c7577b207f2187283040b1041ad43fca0eacfbcdb890cf9b0693c6f3d3ef1247;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd62c6062cb8fa8fa4cbd8bb2a4d105ab1f9b47191c0e68e4f2a7c5df35c0cbfc78416cfaf833eb2878f93fac81950978f608f8110188a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbbe65b4e9ca3b7eb9e74a6ee3a4b0a5b01020b09d637f221ca3303d263590e46542089d6b11c686ddc85ca074690ef13eb26d58e84ca73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ebe993077a47ab809a07ac358eb13ab80a577cc86081d25ebd03926075b454aa73712a2b50db75bc45dae0b8219517a790a5a31adb78a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db74bb2a2d9adfec24cacbe01232728abe467be6a49d1130f5e704dac71dec0c8f5eb21fe699784c66f5bb3f903ab1ee3cc15d5167541;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4519c0f26f2902e37b5d1b383cb254e519e0cfad3373c419d7314f7680fb652de4ea65badec005af4e0fc6e43c51d1de17c40d473d515;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb94d7eeca1298d9ae5ab6f01142312574d343a2b72e3c564260f028439f1e2f728482eb6852a151139a7172858d8fb98053ec245709081;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1f00e0e69575b3a6e5794b7159702b060cb109be1cacb76646efa1eada67e1cdfff1406cc70e65947e1ed8409c5ac7695a38017f5647d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f564dd400156c10418277f05658de09870b8ed3fe11e2530da3e6c3f20b369b6d3b522882a0fec41ca08a4b7f5cdc8d47c7b9d430a854;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3317ed16110bd8d8175ea0825b946e2f4f720479c0c4f7a45ee994eb73b235396064c5bcaeb0d143582242a11a2455fa87d9ecb4430ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176773f595e2e29c37eaeb72c6092b0c6ef22e80fee5bf0eced5b7f0a42dad0854177b9045c42b59f11c221ca8cf40aa99dc3e72e1805ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e69476fe6e1d7b6a980eca204f3dd56115205d0ad150322f155746a32d5d4faffc2172de830440b1409daa47d4510b9cbc9fa796e9a25a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1268dd3c1ddcef51d991c9598c06e3fb3c3671d02a469f43eb654a78b478a070295ea5621b904b9b1335447a8dfe50accd44607250ddca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a6b9f7916c47846599219808244b0e7f18786483716eb528c347f124f47c7f844e1a1e5fabeab716c6cdad85bd7b42d0d630511bdb44;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af077e8c32ae5a5e5b263a3d38ee3560db4b72963c13bd3e4c9393541bb91dd96fed0fc26575d61eaf900d1085586c9fbf8d28b13fb4e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab58864aa93317f2b4052e1dd06fa5fb2bfef5ed12581c48559394142de2a331c9770e974f628b44ea1eb7db993debcbe8cdfdeda4ca5f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31e1eb6a9e9c05c86eedaebf1e117e32b9b1722fcc6e38e1695130c7365da216946173db3e2c040a02adbe6e7347318b65cc33f1e26de0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14520c14b8b0d90dd3bc80f7957aea858b9709ff12f3d2d08976ba0a84a04334d6cbf351bedee95cd7d2e7761da14e891e8691f470c0ca3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180a6d052c7af5a57a41b757c71b57f50ce81767cfcb00132409f99d444e10d8ad3e055c8c1d38f73a3e93d838501d768d17310e44bf00f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habd2e33ce614c1b282f30f371ae43866fd6284dc0b10634c91c2f22d70650410b2c4de65e54020d23239a94b76d1114ae12436f3124d26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3de7645014f6f5456cdd2b91e1074552c15d7e07fef38e32231432433be24a585cdef184c2496e7e88a14b0d53022a85518c355805a8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda7db355796c3c014140a556e6299357e12028546608bf0f74fefb538692ed5ad783f8083f112fafcca62670ff8c0d4fe7e987b7fe647f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ebb0bd2673b2a8404c442dd5d0c85985e6ac1f661e44904a890c32694cac824da4f923524d5ba6fa73723df8566898877c2db58e4b492d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h162d7db83f282b34ce16aba09ab98dca772d2baf972ea94084cbd09e21d008ac21130216020e182b4c9b0a1f02e5511bdecb3bfc7562b50;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69fd3baf6815dfa0381dc492b33fe0a33dbf6771591b3f427737a8c535c5a4891d82740acbc1a42c27d9e045413d6ee773b6cd935446cf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39a4d64915ebf6e50481be0899f37d493b1502c92bb7611fb1d1a632f483d0d63a74c9107133182d65e903364fe2786f9b12d01858fef1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a0bd0d3c647775cbdb35b32d63595e3a234e7873d26b1428d6752635546248fa602c9c3bc116a98afb7ea1151fd5e5fb0df82cb95c7c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5f12d3e27213ac65af54d2ddb15fc515c2f71a5a8ea40ac02846d7a66b14cf59484c4b4b1ee8f8c38a2f20ab12761742b5fbae64758f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de40fd3040ef2f095df2641963417575bf1dc362aa6f7d55156ae7c019ddf6ed74fa8e733721c26c10a2d8862d674d6df9f36ec95fba9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2f6ce2dfb3f36340d5d4f9d5a4caea25ca005a9ae4974faedfd5bdb5df07ea6771dc31ea99bfc7dd30de5069cd36e3fddcf83cdb63e4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc66a0373b580b59df915647fe57d23ad4a27dc2662b0891732e668ac1047dbf1f11d19d3f8dc886846bd67b0733aef89672b68c2db7307;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adc148f88db2517b2c60e31c3c670213d9a34ecbf825c7553c928e7444e71ef56c8fa3fb5d858569a30f4b4b338e15a026bf24e0f50499;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc399c27dad84ca34af14e1dd2cdf874372c9fcd5ab50c5b902996640384f60202f69c2d3f2fc603faeedb8813d76728fc14309c17b03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1277b139c3851b2478fce0715c02c34f052ce1c70fe1b4cff954db844b982925d49bb22eaae98943019f717d964337cfc6989dc0b574cd7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1981e6b321f5d463b0759f9bf85a6e0d676c09f578ef7478d5b939430fc4cc0e7484ae0850e8995332cc695a3bdcacad110bd19a1b3c6d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1834d0b28dd8885a8c431491fa1a22badaa62094c4575540740a9e450938df8d62c6d2ab61968face579efe9b9f7246716d964f8697044d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h288dbdfe213d424138881ff9fdeadf7b287a5e98fd36cb1d5f5f6a08430fe3a125550005f0150ab0481186593d544cb24541d4f5cf0072;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ca3fe5354975968d30a792a13d2f329273afa921f8ccc457ac223308a5f3bff44f439e7768e7cd7e596bd1e03b3959ab4fd23be0c3b84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a827cd4cd3413f0e5af195c31c548bce2bc5db743c04fe9037b00f1ba9c3aa3ad9f0c233401e1046f329c66bdac28eb4c721e8e138c6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5cceff941e4f91dbe9eafcf3b6febbf721ee5ce29be2c252d5e3ba7df95cfb428bb69ce62cc369e14664efaa64da1bd94b908d53462a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175f58b89dcaac059ee93a82b95c6d807e61b252485ad436fffdc6c0e64463e5b32d81e12e92ef59ced63d4d5d1b546e5446678c6f5888b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7345e7df20f611accd1e43454eda5ab1c24ad3a8b2752cba17a2407348bad0b85f99d869a8552e7dff0c5efd5d989ab5190913d34800ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a56f50ee4f3e72e4aa2505eef2d9405de8f62b321981049fe97c76a33c5058b177132bcde13b1081bb4e88de71e6c9eca816aea0826ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a5439e4af4ce51656349bd63a2058483ccf69591260a2912c03c3b6fae9d94e8b559d70031457c8b61aa8ea29f53e5faf2697fdfa30f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b8d2761563797d0a4f9552af86883a63698d1421901649ba0d74bc2ae1502fd129509daed5b5c73f4456f8c7c9fd146e05b28c4c7f195;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1293534cda8780f1f3fbf72c5fd51e963781396423795f73519f8e5c1c4673d59b92f04d6028bb9f6331c062a58498cc49225540da38d4a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c66ca3541bda25858b96153be03fc37a4b4953dc50698fc1a7601db1b19dbe4df37bd1ef043ba8302ba3222cd5ee681ff2415c4e13f61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h429b1f3780aedee2b9780fbd11f075b7ebacbe533a92356466646777b9e4ad3e34eb0d1f4b722b5819f35ca196b23aca998bd312eedef2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17beb780d9da41dd0b2c23dfd895b10c3315568fa79d1407d4398658b8056d4daddf34d08923d66884c9edc1fdeb728adebcd1850164701;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h867df6e2267e4c3b8d9df792e0f906b66adcb9d4bcf4673a8fc4f0a3a18d94dbc872aa1fb565a0ca9f8bdbd264f45d5d4c8926eca245bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb0f9c36711a858e9c1cda64edf193c55469ca60473a8bcd1d7d60a024228d5961bc5dd4e69f02d72fc0c5b34efde0c41e2cc71bc7c541;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94a8194250b94cf7770c785adfa001e6ec95b975d7bd58be6baad8f0aea32d1d0a5d670bbbc8c249a335b899ff3540b598ab1002b57a01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84bb8f9c94f305c9d1aabf7536dbf6c52e1b87f32f61195c3318f0862ceb500217b32ea9cf28272d514e1dbfbfb888b6f80d069fd559d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac9fa80defbe8a9071850ba841e90b35c186178e7c8c050f33a8c5a776c1eb26ef45515c81e10d272343e57413ffaf75b65573413ace92;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3125f4715ad4397c3dcbd304cdaa627f88bef7d762099c2a7f50301a59133b25dc5325e6b45f7272946c821d2850782d95bd252860209c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19284e9fd63be37a5705e176a1c49c7115be9aa507fec4a934fbed4d1f56b661c305e4483d50f72ed0da4a8af82a18581423919a2963f81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8210bb7a1b3278230eefcac557116d47af398bf7025552f387c02b451595a47a567b6553a1fc3a8ecb1c9129284570b34bc9256453cb8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ccee8a4a6f7307644dcb371d13342a42ce2962aede7beada28d2bab0cbd14ff6c76557a26fe1ad3ac246e02276de15e91f4ca227b1768;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf7d63b83b921267bff3903134f3b2f5a80e14f542a60790c243748f0aecdc8c35e4a80b11eb340fc25167811879e709e7f64bfccfab93;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0cd4538d4d834371ea511343264d24ddd2a8c98bd70b7279545d5934b203f032961ceb317d4a99fc08cf16ec5e27d54336b5523b99732;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da5e216f146c06cdb8056aaaf4d81becf42d974585f2bfe4f3a4001fdce71d4384a5d34a48539a2d91b0b227c4fa2cfb7608af238481ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78fecf87e89ed1e7389f752f6280ac815771ee048c4c2105e4be16aeb97e13c7f6ce4973cfde994b2c6597304f9652d06346896f2aed2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164bfeef0ec06aa68170fb8ec7f364a5aee54a59aae4f7591ac3b17637189345eeb9848f2669ff277163d70bf52d9b9014f09e49dfde2dd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19800225f323a132f196742e849e13ea4b5b89fca83d975a4ad58b9e498dbe7c959901419c7dd51afcf0c936f59f3a6c8decc6b136abebb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ff4c45426f07400658dc9203b0b3533292a15830571e7673f75d3db7db300059f998ca65050f8f2ff3e8876754b85fe8b11315936e0e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19323d0f70483d4b5c7a48a7fdfeb0e11ee42b03507c6949ec0992c0c6f0645318db8dd49be85b5de4e7fcf170219eaa17751316006086d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b199309e35a043d0a8b1fc979ff40c0971542607372626750eb8bd34ff9c97e868d9e4f1c935b038978bb547adb7e2c4140ced9c4337a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a50f9e564e6f70ad82cce885f065c5f96fad50644f449241dd9b628c6226c64023d793ced4ff2473519c30bc5de2633e88b0af784c4e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a412b1cfd00e9a03ab88c1885be11513b44e06f49b8d8b1e477a9d5b08888cd0a72b71084dca47dfd8a2acf8560381d37f4749696bd62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9c18c4a5531a2713aa7865fbbd97870d2d7e32156b81d353ea9009b31bf16ab98ec55fce449ff94b94605fd29ff3ca2ebc144396c8a4e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b2622f663f88fde206da30cdcba663a4de7941a9028ac0c24284f0c5038b56ca9871642f1cb83bb880c80343a5555248c9d0aa2b60131;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf92fb3c3ff2e5000602ce08c3c9dde83b6d4fe914af5d075cd5cd8ca6ef3c12a1f9c332e96ccff258aaef163c86a486d130f11d32dc7a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ab3be93bd9ff5b967de4f2635b475e0fa6dc2921c8840508efc3d667740697fde5e9d53d637584014e9619bf6ded91487cedc9677f4b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e7ba8d0bc11a8779abe6799a7545bba89209cc1ccf5acc90a17dadcb6e3b0f650b0c5e916129cdd39fa5be0f97d791843f940555df084;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138c992146afc6b1c8ae5c900f5b0454b044cc237b97f5355c1e9f6596470d3079f5aea2ec3fc6493f22e82ed4f503ec969b777f6422cd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf5e9e11fc8c13056983ced9f333e018f2bf7acee6172877665838b5f9c5b3e77e4d3e786d80925300147beed751fffcb09df417cab7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1607e096e48dd2805c76256a78b7045e0f70a8fbcea1c8a821571b9e6d24d8e667f501dab5423d5da2ec0f7c04b0e84c5fae5bc0df35044;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19125b3577a3a88fa15cae37d55fc8f91ed57bd51400e5524b100318688fc8d0f7206f8591b870ef561661efbb5dc6af5c881cd234b9bad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hefdea6b4d86ddcf719c5cd7f7f76e5d42272db2c053e903233952148747ffdfaebee5fae00b58e2e7956a3016262c8aae6afd8ec945301;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hccfa18bcc59ca129044a6927349f6c2a1e6896321e715f637576d2d252380707ac11b4b34d029a75ed12596274c71e666cc0aff9e35dd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6273672e29e27814f1481675aff41e780e5902d87f8490e84fd33a1fa372a7d801f0679fd8edc57fb520919b06a44c98c97ef926b386c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h632899237c10ee270c89bf022ce89246a5e486fce9ad7a23ee5d20c281bd41271e49205fe3a8081bf464384b28ff22e43e002fe03b39e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h750bbd25955f29a35e4b95c9cc128eef65d708bba8b3fe1fc416adf4122c1a9c0b946a76422b3597d82ec5ce5b4d2b44d5566bc1d8ae27;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1512a41db82924c214a4575a089f4784197752103c8ae73d0e1feb192a27d59b04a62fde617dfbcf69302af61c9bfc26f0fb9b91956c752;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8e5340b293f47d44dca9724e9e50f523f53e42e9f3219533ed162a0e6b2c961a7098d70934be2798ae42949baa552208fab57e1c9a5c8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h578aed071cf4e673620394559e2af5dcd86b252c6d2ad8e0d6a70ce626a4d5d4b96099af27e50901c80399b0f77509df079661b0803b97;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128adee8326a95b2c03c13e666a58b8db1b251f727662e9305bb645c0b9330aeb12588263849e4a7294c3c777c99cdffca51cb21537bc5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171d050317925ffa979c33fe55232ffd5e97d84cda0c8e1d04a8ac16424c42ecad6730117b687dd47037c64865a180d558ea3153899dd69;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc69922e2e6ece8c99fc93908b8ca17da8a1568bc317a39282ab98e466bd405c9baa143bcd6ff5d9fe6dcb645fb7ec2ceacf4480a6f063;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103bf481cb77e4cdccd98e4f4a794a5de43933872eb41e3542d69e041e4f639cda1ced1918cc71b01606f96c7544cde980a14d13194ff9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179e8dc724d02a991846d180a71a83df3ee191c731a43d4e3ddc660c6d9fe04ad4e65cd62ba14f7a02a39f313e9edbeaa014298c387150;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc8b101e073d501a59876312fd7ef86f107c982b0f5bb21b84d9cdc3b7d6ca67f2454ea28a4a8a783ea72dae443a772a489ed1c2b27238;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3e782a526fb8336676c582545c668e257a03337fef84d4425caa23cff321a2ea808f344987acaeb94b4d52827192d1004dbba024da289;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf96e3ca41c231811d4850eea3406ef496ebad4a2f6e08bf5cd1eddbe4e5393c7a3b978422587b003f4f313a8c63e8c76227d0a367a189f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7851f344085a8c1ea293cf3c5e0fc68b2e971e47a2b86d42c2d537a694f950285968592a9e3c910b522ce7b7a79d268bef39463cb8220d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd546ab2223759f14af11d663c75dc358f0b82d0e0a4ff23ef8ddab63880ae91a1eb71c1b9e26805aaab539aa011492ee8f9b0686c3536;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41985a4be287adf92a6c4447407f89dd9ec365ab05f3617a9752dcfbfdb115d56b5b7ff137cfb5e2f9508fadd3a012bcc9b9f8f854acc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h118124c648b19add937b6a942ef4895f6268ad2e9d5759a0b11f52e266ee8dc92508c2e579f4e819d5dc5d982e93892d3cd2bcc1f7bd2fe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae168624708774b48e1557cd83d49a6a2e49a8bd5ac3535d76b2dd68149a637019e1d00b298a64100993ef3e67205512607d9830684a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f9ec97b5064658ff68042360ba8ca6451e8ec52b7a3acc81fd18c383778c5f03e6fc2823b577ece54f46c4588f270d9b5036661f68c53;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6064a2300e7c03bfe3d02a68b8e7080f83ad5fabaa54956498c62d42547f2f6a9b12d4990b7d80a3b4518b8316757ac3a069293fdad7b6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h463a8446766bc47f8d096345aa65d2e427271c2051619153a371c4f7ff7cf30e90e0a06f355927d949033dcd1dbd2c09a2e8ba0882a98b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15eba739164d9d10b40ff2f1a1c6c845c847963c98889ac8127ddc48f57af78603b0467f443d729a2cd27e38409cfaa40ad6acc526ac024;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11519def9ef8f4763d7c51b1e520f48921bb3db23e366e7bc78de95bb3a51d49fb88e9b70b854b830e05a29cae50d0b1b8f9ec530012e4f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a5799c312f94d859d2e024278985a691161b3bae59bccaa03a99497d900664f45e443336606d1242c12bf7bb02398d8c371d74b362dce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a7063482f76176bed544110590b48c17853959bf7690ded3a3f8d3438457e721ab62f6435127bbb206801be07cd4dfcc473e08d200b03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a57d645d3829481e260bda33692c2af1edc1ea1b20c6c79b2321e54127c00fb38642f803dfb9854e2efdf5f5440ad7e819bccf1df1203;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15348192ebfa60e39df63bab098f8ff9436a8080b5fb8e0bebc6d196779b46b0010a25b02ab73bf1d0e1650b3779c66e8a2f4171b4468;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ba9f14a9db804dcfbb88a8779d867e872df14bfc2b228d0b16b1de260ca3f258ccc43b674dd2efdfbd5dae6c659cea23d73b6db0c2c88;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bab7b267844314964311ee2d1c35ed9fa7c987b7150e8f62397086c7a3ef1472b3651fa43fa5169c0fb5ca489dc53516af5e6088e8d25e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf6dcc34e95ef52a262e141f89bd1cde3c2e8ee5b29cd3348f02e75e2deafa11d14937ddeeb2a54ef45121c585170662457373baa33c0f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca6c43a5b8007c01a09fec27e861e4febe78bf072cb7546ee08924c521a342b5971f5dcba411b7c621a8235f82fe1ef42baf9e14665830;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf898e40aec47723601ef879977294b4442001fa99ed372891c1ef643a9ff0a7771bdc9268629f4aeafe3959fca29b420511bf55c383424;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e7ffebf0b93944612b48e5fb130922aa7bf93bf7e62fdb037f338af67ce9e99a7b1d8f24642d183211c3f5087fdc9a7e52f05d7b91577;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77b659d6a50b8e1f3c46062bdf5955fcf52edf26d46039e77e3747c7db382b6a687757cb5316c7f7b98434248ad0feb449b1e6431c0c5e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164b4a31f481bf0c41fa9ce6047082b25a6a7f5d5a4cf520df02c498590e96471101ce05bb103175d3addb30028692bfe0e19c9413ddcd6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af77dfb4c8701bcafb795baea16ff3cb4258fafc83241d5944dffb76759c3758c1d238563897b9a6118c03ba242525aa7eecb3926e5802;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e4ef5b19e0c2eed6f264f11d8e95c6e4103e7f66c1d9bdd563dc18e7730823ab56a9c2ee2986d84bf903990c081787bc872f679507f89;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e9b2511bc03e88ef35262f6c0882a7f030f6f33a6e3abcf3ac7fba8867d7116dc031f16db52293564cc0601d1a2fcb2081fec44d4dd1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fefc0b69dbdd815faeb7ef48006e0c083359a155c7e7d73caa5225cca79619cccaa3d2ff1af6c119a61b67192b56a92ff02ab0205370f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80cdbbb110d2827e31480a55d0ccfb61ef23537dd98c3151a26dc1ee6043da1fad4dea996e9300312cee00408903e7c57dd886ee87526f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd2ae4a7da89533cb27272321bedfc2515f0ce54045caf37a4c5065453f1129b80accb67e3f3ef34cad43c7c55db9c14d1e7215e40d965;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb660fc79a8fc905d96cbd6a8f294be2b51e382898e8c794fc16963d689374d6a63c2a1e94d907e2cc5f83d8ef61e04129a8e8bcea07b0c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8814f24c69331711db8da86868dd3ce753fc83fc0b463545dad475db7e83cc049eaa8ec2ee6bbc7f292e7426b738c489e26cb867b0b5fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190dadc5ab2c34ce705f07b439a895b630e74fbef711ef75985a94ca7a0afc78263dc3abd6f17eb64882e567dd710af6a231c43de575af;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ff95be02fb73f64065f39c024cfdade2c8f119b1b81bc07477f33916f467612d3dd8bc1003f82218b1c9f5afd9fe5c75398546cbc548e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105289223563e012eecb1b988fcde8b3181351034db220da1cacee4a45e67893b357209b9147e863f86dd87dfba5b1e17d47889da19fe98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h295b128311059506e6bc49d3eedd6aeebe3c6f5fe25c9ca17533d165b0bd452b2b3cc8d59adadae987b61d634043e08211e488840bbef6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c009ffc76ae46b0feae4856c5310e17f0e8983a2195251266c796476fd3e0bb14cc9a00b7717d7bd536fb668e72ae0a494b3297579946;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f19dd7b5087b0b142d9a2733ae43db7f09cf3bbed46f7f1fedb2a4e2c25ba8a53b5894de0e3ee11db61bf31335134618d2ace712e4c7e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d800cb7f01bba171e08a3bf7832493ce28dd3b73aa79911227ce931568dfcc554659273c6bc45930ea91cbfd9c6d03f0336fb0dba75566;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7ddb490e915eeb46c2dd78a90d856c9c77792aae3bcf12812514b878f9374677e57e8c81035e987a6ccaf495b41cf1b5f5febc995e169;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9651f41fb31cbd4a4a1ed872b1ecee4543c393c9fe0d0e106b9638bfacbb30a7e307639190de4b333df46441de25b35cc006aba0890a75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80d0a9a6d007efdff293bca332e22d61d8b8fd5efe70aa9a5a5ca931b7cb057557032df7910537861658f58a8f883ef957fb4d6589355b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d049085edfbbda4be0580873811a715840060d75140ff11f0fab23daa005a5c4b9a29ac194109b24fa337b269c27961e4471337e727da7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aada99a6d6ed8e277a47ca38fbcec45bffffa62fc03756e615795a1c0f8b97eb3295c4a37cc646554a50c06d934b722fa1c607034e496a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f8500b6be2ddabaab191935d38f0484c08099ca4a4ecbe34c0f161e2486e652c20fafe9f0ef49c1a3b8b12ea5070770f92b77214edec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27fafda8743b116798efb695748f1cc5bc8582b658991d5ed12e8932335b63847354f384a07a8d5dc265dcb5e17d5e787c555fa85a153c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bbaba9e06352b2116bb03ccba54436c7e9d59ec8174f32374f4dbb2efe80e5e9df3105195377db9a88cb46b65806965d6cfb31cbb6e07;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5fe95dde08452c3d15209e8353e898a9a6f4288867d3715a992b474e84bdb811bd51671a4d56c2d1e5b6a1bb4473d80abdf713b09815f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb253266fdf7aa0fd6b024c1a9fb23f24dca40d19fd7b9166f577ab3f0549cf18bc5d8a013a3a01b404d97d5452f16b2fcdeba4ec74279;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a460995e287b0683fe204bd6b97bd9ce1022b99af2eb050f06c64680a610b660011944bc80b327dd48d63ef6252644d76cf2482bf3f6ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95f6e1f29427870ca2e65705a9077b2b6c9aeb9b01161bb7b1c2da377ae3ccb2f068a8f823f1267cb8bb1a456197acfabb052db97aa570;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe7ff429a4d714c7e167a84a218ff2f475802e091f4b5bf6b7ab746679f2d4f19a74af9982a6d996e7e5803fe908737d41e205761ab194;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33b02b68764ea046c6517869323be8bb292f05a9acaf5e97b91df6e8489464e56b9b84c72456eec4523eae22d02eb87bd35d06eef6fcf6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1707a44a011ff4ad4cadd0c505615622d9da446be11b9cff738272a996fa9a2d96cb422f8aea1690541ebb544f60869b26b5695636c1633;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0a2a19b98b46b80308cf0233007b026e304e665c54e9b1113ca419b1c80f3def6d507247c5a8154d0ab6ef36fc4e00593b58996576062;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5146e12018208425f19a3c74cb5b283aefb9354b94c7018a07696386e6b0202fac91aaee3853223c41a3293e561e3359e06a0b129665a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2a1d4663e8bcd3d0fdea1fbe2273c6d16ded114f83ea4e9aa2ceffd2cb58bcc91f8c2ebd448616cf09d8e4bebc65e0b92a93e62b2d4e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3da701d41fa8d3048231f19af9543ba827320b9919235f3355701d7440848e47b51f3239e1f19c9642cbc3c8128d99dce9137d6407fa05;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1301351fb712e62546607348b675f9564a915fb31972c6c8868516e55897b37793ded7461a10a38a45d3e1799f3bffa54775bf28da2cd84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d532483db04a387dd5f9fbf5b21df5f6d8ef50b2262c834a4e6798ea2cfff1a558da9672634b35eac43b4e229f05ad1ccc59eda46024c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h131851f5c5efdd7d703bed2742b4fa9c78da960095fb69768954f87ef284f8085d94ba56435cc88054c3514773f2530a6aee5848d373203;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf99e16480aa0a188edb3a06fe6e19bcfea3851fb4df20942c7adfcc1927e8bc7fc73ddfb10928643e01359a56ee4d09aa6a852ea574f4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d3ed70535536a3764a4df4cad45f37cb1c5477d0a428ea6f14e8b0c2ec62d0857885f1bd5032054e4ebdd8f2329bf6c6654d57663d89b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dce68f27b52d0e1277884f2fb6caf531555d5dabd0b9b3183c7451c47e9c5ab580935c51b511222edc83beafa08dc72c7571bd41b1be55;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde0a3e72aaeb1b6f593e98c25b4a2a9a44f2a1787e7dfc0cd7e9494b6361b0d511247e58e1ab86afa01282de59239574792a22fbd7c761;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14548e16f1de57d965e4888c98e262fa9e22a9ad90f1022f9431c1e43d91b7d259f484ff69f3c14b7b9f7a13c1ea355773925e6483c2505;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f7320ccb30c6a242389a2f6ca64cb6bad0dd591ebdd002bbd9bbb69c9f3198224348fb1d6b21eb1b63a2d617900cc8b765fffa6123a09;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113b93cb88b9f164a031f1785ace9de07aab86a193c39f00eb92ff8bca73f7720ba3c30a730e384682d3468e77b76b298f20123e122bac8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e5c1565d95e93c3931a0c3b998d2ff4d39153e9a6474c4daaf12889674cc98dd49beb0011fca27af9685e7fe9c2ad75688601d2c9ddb3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha441df7e9f74ca7f57048b00ddb47de0072a2ce47dba6b4b7033b1dbb0acb0431ecf515786c9562e5da5b1b28e5b7c06963b8732343da3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b2452f9d1b637e84e2a9dea9a8d112c2af88c5ea4a4ae7b310e2ab469d610b1a3f74ed8d134ba9f4c1ffa76b22e66d7d1ebf334dc5909;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afb81a0fd93d725b4ec4055ab1cf8f7ad81cdf0d525467c44e27a32ecba8f1de63b8305d2e3852d57916e00cd94dfcb44f5294b7d723d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h565f5f0b753af2034932fefd19951094ec80bbcbb708f4969a2dd216ae92edf2c050052dffe8d7062b5057db26c7c88418aa44821f64b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h321d6643d73c8145fa4851cd87ad0d9a8ad24d9ee1d00ad7aeda990144e728e4b4863b57af1d00134bf8ed890a816fa8dc67b1fcb67724;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3c95269e5d7aa83d5c6579474d7830c9173c5af2dfbea93ade2576b5466d9290aee1a1a564ca548b1e94021fa99260eb32dcf31b0bef71;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a66704ff87ac358e795837f52cc9ea67986898086ab2fb9e89b1ca2804f3b5809b0dadfa92161ae761b3c254332a2107fb5e5b2788e476;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f78ae21cd04f6913f28db5e24460c79af2dd0d2bca615161eb9695d15ee998ad60e1e1a14717d505899e699846ec76b557892bf967705;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54d212c7a08e2d32831d4a4425bb1d6af283e11cb7593bf584fbc02d3d822461c1565744566167a037776e659dea675a42be916f9bae4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca9d8924c9975a27f17534e6850430bfa855e5e5968c9addf0f772567092efd4e5d322428b0b0134779433f2685a35695c0b43c337fdc0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15fc76b6702a3dc45fd0783485c8cba833d6396ca1b1b4b1898647e031885e3ec24b04825d8359f65b7f66bdf96e8671e0a7638d2b12658;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6707492618eeb4f692657f998909934f4ee88118251b02f92a7dc7e5dabd23943d20c8047116810a4a2cdc23931b97a1f17df4edb00326;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8f6cbb3d3b2ee659d521e726a65f319b7667ced7c959a8a53afe2e02b46c53e4c2530687f29eea8a91686f80d89ceff3c73730181f827;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d4e158684a27e5dbacf5cec45c033b06d67fce1597a9bca0203bbd834c0d403452a608399cd6a64fc55d74077defd914cb6d3bf3af71a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30a7b6a9348013e9d7b7bd06c16c832f4be5747335a107e482c4cb618cd3c96294655c8476061dc30ed8c27c3dfae1ea87b772f15fe69b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14eb537ff3e53232742597d81cf07b725f865eadccf1be57bd86080920032af2a4df8eecde7bc4e2b79bcf45084add1760a3444095df0fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he741c500efdb49edfdc84b34b539885abfa80666532c103c88bb283cb11ac6844b914decfb10223c6403118f50f02390f8c0e7e97d0af1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c01992647ed70edd948b2fd0bf44b04119d7374ae14ee443e9cad05e66c17ea4ba36ac8d02e101defaeebd7aec927b4f12f9f4c382e980;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e3a1942a3d989d83b719d505e1967509faaf54cc6250647246b24e01acfe32ccfcdcf36ba9df99cc3e19e235445308a6868a7518828968;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a33e4769c0c942973dce058c7dc072357e4b7ef9c6ed625ff1dfca86c0d17efd6de62003c7dbc2ff5d73f6ecd210924faefdbba8a352e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc88102143a15bc99f0867e73aae540cb7ca5abd2f720cd6194e085c02555fcdb2405fc4a8516b6d1d2b35c330658ee558ef540cdb6fcdc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h891d922d4dcf5d700f13e06253cbc1652633f21cabcc72cd36f4f87e4175e53a3ed5f5b10873ad01ec4dc0fd7a4f76dece8d6378bae322;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bf2c971632a6ffedf2b5a8c9bddfb33c4a6e2b4c4c78ff4fcfa57a8e56cfd991b6dd15eb3ebe21fc2fa2c88ab43dbfc48313422649aad5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8389cb67d2f961784d6c5c995730106d02609a04442de1dcee5b7c38fc81e0e1d9059d711d1b192fde9e3ddba1ffc01370a2e932434ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198018612164f55f6641acfb0f93267fbe0913beb69894b810250960a8ad34b6b2a34d8495cc9e6f381dd50874d5c55186856a3aac85f9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0d4ea343366fb07a28a676cb54277706a84df5aefe51df5d3bebcc46620c301253778baf3f47457fd46881ee67985eb69f929b269dcc6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b704d35e17403370637aa6c605fb46e1c629dfe86dd00c0a2de664a76ef30fb0528386a5b77d37ea8a568923c0896638262c37ef9e04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba05f2b0e2b1000285f5574bd4e76b1a529db4b9cad06fa090a74160065e80848b0ba64e78bc15996bd9e08a333c6670c6dd523d96ae3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153ff87d04f7f1e53c7aab55e4e19fff832c41b98693a0c564dcd4799a4ba1fc5b14be02b9ac82cf72bc42ddacf052ac828ce33f60d8f85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e573f788aebdac1c289193eca59605151ed213d2be39d60494c98ee220e930e1c1a4c0d6ee44337509bf5a52dd94278d20773478eb43a4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c66770091ee9923857b3f836aff7180520d61196c84e484ecbd5972779d412074cbe11092e77a41e9d9e764dbcba623c2c0205f11707c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d19a1e8d0e3653400b3ad5bc0084c1eca6e9e98b5be4586fe8fd11a50bccd151231816c95e2c79aa485ecd95c0fa24c64ad7f0ad9e74e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2a28dd5fb0a43dff2761eeeae41400689e9538368bd45f54889b04c3062ba8b5219eaa982aca8ee2e567f45cc6cf5fe945dbdf41841f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h40ddc62b7eed59f76d313c182a698891a332b83d087e90b8312125ffea054ff3b7306d0500109db77881296bd844ec1fa2749519a9931a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc62dfccfe4b29c474b993251a1ccea444e7fba0ef855da77f6f85f6ae8b7bbdab845509a9ef4fac65cdb877937abb7e4fa34116f013ebf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d9f160109305d6780d65965fc16948fdfcb7ddcd9d73fcb9a514111b819f6863608aed6fea20495ca3cab5b78ebb42580f2de44245df0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ffc03c2e9376c2032d3b5f5b8f93843a8e1242d09c633fd53444878d9045501b99a39bf9f1f1dc308ce413224dbba8b44694d780d6fdb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b50c12e67b562c0eb0b095486c3e346523caf015061d19ae412c1607194bfe9da2efde4ecd9992cb54669a1f2c0188bed24bd93469315;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b41c411f4e50ed6fce160f87b9ce8cb8873fa28a248203ce22ddbbb43e5cebc27f5134fbe4d275c2322239c15969c13bfe575ed0478fb1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afc3e9034c01bc3e7c8221a2cb1726c83819b80f6afe27132ad809996959207e04442513a665488a77e2e54e21b23b76d047dbcf0e6302;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddb547e5cbb50cad2eaec7512864d8fce8c6070585a539abf2ad0ad24c707cbd7402b4a0fb21254708f914c719792343da1e87eef77c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h699fdfe69d66880307db585f0524ccfe2f395114cfee2905c282111a9c75e6149d4c439a0aa2ed884a244628abf632f7152e6ea15c09d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18bd573c66d080c2a04b1af334bc31d0a66b28faed79f0700c4e47eca51056b4b38eb687f82270b853fd8d415a550c55289f812314a4d20;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae688b6d46c181b2867df5d27e285210c9e1675aa5acb255004bb40743511f473478acb53d1228e3fb9841e577e5aa4eada6ffc1311f52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5cc6e901b49b319d29df90cbbc9c25b1631f197a39e4c1ffcb4dcc488a6eb13630be39964e58159d6c0ca187f66ab1bf0481fd3462b78f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf94fa70096ebde55e05565b5b75084652b9fe30e4de64d1a89b5d6e34c0fde28dc4317b1160a91489d5c5133258e2647b8329f7954858e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe16c6d8f5ec43f979ade3f87f99beb8ecda91628700220b57759a93bfd707a6fc21c00d16c986acbafeab4a6631640f48f5e87a18fd17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1877e1cb44e1777ba7331ece0a63b6e41653e02f2558efafec03d0997102ec79e37c30bab27d99f39fd217b66af31f3bd74ffdec7271f7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a6e096303e5d3d2e5e0b105b4e7d30c7578a585c7cb8b2208834611e6dcf98f2cc4a28385615e4ba8a0ac7a4172c0e04ed3654c40e15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he74bee671145efb1d65268b68d51efecfdf0cedd7ba9944bcf6e364f1f85b24c5db64a37e906f277b2f8bb7ff5cf9356813e60f1a1dac2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17dbd3b83573b3f1bf624d4c2f986914889e758545945b54b99640b7836b4b61a9ea216e2b93c5bea088e7c3aae1c117303725708049f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h337cab529dd2fd47a7a3410da91bc03eb6839ad31ce587294e3b3d8cca653f2cb252e1d4cbd8fd6101687835a0fe25127f1f34848815ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41e9deb05a4ef4b0aa60e3c060e95289c25a204be8560b5064bdb9e3d34f1de42759b767ec1f63ab63485ef231e4b345a135b964e0ec66;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd168306667172a7126263ae085fc2cb1d0a2af5d3323ef15a52bf00c62a4659761b5d5b4aa39c079e7847bd373cbca570b5d4055785b33;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14bc957a260a431ba3264b766f1afbd2fcc8161726c063e1419e1c72f21edbc66dcbdb4bd064084b88381a8e96e26c1ddaa0745e746cda1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h37db105946cd422d6cbd1d33403b378a5a3d10a96364fd719a87606f24dd8b8217aa793e509547e5f1815df57b0c41fba29561c55d4a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d10d055a6d10c2addddc8ee43a43853a6dc44d2517a6a5680964e3413a8d99986bfeddc57b4e1fad5d80c90c2c2a340b411d2c49b24e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145c5c02cadfe1ad83729f1021e15ebbe3fa359195e6f5807c384b7371d9525a44d6908f0b0893048b15c9842ae921dd4dc4c07f5e37511;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4066730ade65e5ee686e8812c51c80e8d5d6996fa281c5ead6c9cddf8d88c2d91f233351b4d3cfb68229d89cea4717fa096d2d53556d5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77cdc644d6130121b8e8c5bd9e4df86b0b5e7827a3831fcc438fc6ad911d39aa8cacc251f5a2e9913545a3748dada0757c62c3a7eedb0e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e190a1af226cb2f3cb5521a580f366e4ff280423e98159feb2b6f4b452a81eaf3533b0af04aa865782d5c39b7334eb544a09c377a69c65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d148c064e6413eabfd45db820124d6eb75d2d0691e610eca5570583091a06cfe538c9ff6c6cc938c1c2a5b803945940a7b2c976676ecb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cdf05d4ce98f255f4614ad6dc912734e229d2661ca3674531b40d0e56eab5659e4ce742e18d5cd29f6be28fb828919378efbec743b939;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14aaf4edf63a958335ee927ea8eee4f717e3ec07dd86b5e808b69c0485e427c87a80a9e4c6eda09b21f5eac5cd0a4e23aad847c03e35c3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heb4e5201dbf019456f3c29ae10d4f4c14ff43bf72c75fe48d7a1d953c902a742844ccb48c0c780bbb5f9777704754d31534b197d5b20ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea525c86c427a85afa370a83f05992f0ebd0dc564d92f3b1433e4e80a7d35e684f92871b767aba0ec2edc50412024256a20c47ff1f5b9c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f6e737164d0fbba8f0229c8542b9b74e09bab7a1d1422f867e87d93488c14e5ab4b63f7fa15191ecb010242655c07609953ca4ec30067;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16cbbef628d34a2a1f9a844d0b798691f6a33a5df461e62cf94c1e37fbf174de9d95725b50d79f605f233e5f5ddaec4d7a737e05ad76522;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd497d1f6e48b6c8a1f6ea04911493e3d46aea5754fe0cee203b75b1be43a9ed7daab20b74549a00ddeca47f66eaa65f58303c35b225c74;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c220857eb9e9b0fe4303b7caae151d2013035ffc651b08563fb6ce2e46286e7036a3404d3da26f7442b109700c93fa33d26122c29ff656;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e466614742cb6b3de01aef2cb16e64f709fbdf33a7e02e7880014bad4af11ead206709bd8b1fd621e79c0818d578c76d95e9eb4c148ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6bae914bff4512778edd5531297ce17c2b7697d71921f1dd40a683f742d02837e59d9903df437460d2aa9493040d3d11a24651a7c6de2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdab35b303a6b0a566fa56ab1fd7395f309a08ed7dd53ee58c0e5eb87121e5a15758dd328836e4935bd420d5c224793cd242eaa4ef6de2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h695c71dc2c71559ad1c1b7844e1a9e4df415ffedff2302fc3b47b327baea56063e9eaeb08f4f732dfd90124907be9a0bd5a4d5ebaf4b65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h655cdebc0289c45ea0a264a38dfbabd897859f453b81f894e961198b7cd3ed095b262780db6d579f1b38c7bfeb8e5b479bfc8ee64df1be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1191001d91d3ec689a33170983c021f8a3247664ba032e1c52b1d8090ea4725c7ea3e97d558506d939c73bc47a5e8b2a215bd23675209c9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0e2e5c44d3eaf35fc119bfd137fcf2328f9526e66f630de37daeac4465ef3a2eff51cda703d4833978432891b4c24140134cf3542b5ee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7cd90602f1a68d79e17ec7edc732d87fbba5142b1b52630ac180a4c1d882ef2ac6f8389e0b1069093bc5c6437ed596ec48425b2f6319b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161d8223ae952fad85b492b31f8eddb8603c0072061b5105e446b5cf4f2328e606f383377979dc80940829ebe697453d9c07719d08ddadc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a17b71d059eb60c3daadd76baed23d0590c17afc6bde5dcdef2be84c1669c8a68db4e8bdaf7a1dded2038e867bf155ff81405e0ff0b59;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb0c4a0d520a5db800dfefc4f38c5bb0649a72a32f28db386c7d6015379f178c90b23f6f04d6c74e6e61216b4cff4f3c60bdba57bb9b02;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b65f0202a7e0c08f6a95edf33295616bed4a76588daba1f1a9bdea850134d41ceae870dc7163c2c42113306caa3e6b6ef811c0de7657f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d0eb465601d9922556d9de2e9aea0c779595e41a88e4f81976a52b0fdd654b4f6891eb72d1e81bd8835823e272580918a376e0a0b615a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b93895626b5dc2cd541c8d98920c7c26398795a251dc1b1c59e8a76fc063fc6f05fa7a38994f292e2fde108d42d3fb5099fc5545f21d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1358b8096b7f1398fcce7d0069db0f50f8ec427a6693cdfa485b89573023d63cedc13bfff91d2d7316028cae05f67ecd3672c42d9e27cfc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9b4050f64d2615cac55dc9e6cf3d263dab748367b608c311d7db22282eed85bda44448cdd2a7be17f5fbce2df55c1f432e7bcc1183f51;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9af291007563624cc14f97fdbe8ddd4aa476fbbf041ed6d98b078c531214efcc0c85afd8bdc9adf550604244e4503c31e7ea463b0b635;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7187686bfb64f0569dca140b80a0cf99715191c0e92da21ab45ab45a5481b402ee09b22a5180048b8ee37e499f202631fd458f00404844;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3197c8218f422ba5a330f71826661de3c052941cbedc59adffa7272422066d2a7bd9c66de2ef45cc7f0d8bd00df719349c9d8a4ccf1a17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e963ffa9b5da2e5b9e66d68281cd351990675c662d7d8dc6a64bee78d85d6b257bd9cc90864207ddae85e3245a5860ef7aba3e03325c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c26c47a1a6d20f59311beff5b5e14e5dfddba354f758d01a1fc2e305a9b7e48bbbda76871d7193c1a9161a209b813171a8c90e31df692e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2dcd1cad9e23d2c4445790af9792b09e4d90f8a822690dd5fb82cbadd92845d210ee6ced62cab49434cef835cf99236b495c0703dd7e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c03b8fddb14a85447fb8d32826af3009cf556c9cc62900268946b7e6122270c455736b540bc2acad5f3d870d17cd2591783fc100dee141;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96ad2a91234c2efccfa40e04dcb81b20e81fe65368760a56a7f0c41e96c477db03df7b6e601ad78b8d7a0cb4b9975602bcff335ebbe366;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c31e375d830ebc110ce55bf0b0d2e08df430910bb9167d0d297cdcbab0574c4075fd1386f05588682d3297254c233578f7af9ba9cace0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13fd7948ee661d70fe74c83e1c165ee497c3646c8fb85f541f5fd8a3a690f0802f69344685fa23d612dbc4e267920bae6f331b791612f6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1557a66c393eb666838f1db186796f1fa241828609ba8555765e0d904726280773d8ab16929017f48295b5bd2997c1b295a3b49a3ae83a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f4e30480f8d62762fe178743d5c12b43dd656b8bc7f6d3dbafff836755f2ca64edc265594168967434c7266c9749483299f00f59fc9fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1698ef321405f857d0da56e45ff41bda60e835b57f1fbddd82e2ac0947b0e36ecd47c1a04ee39e4bd0722c2dd7058a63bd472e89fb52a42;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd24d0ec1d4bce4b6a48b7144a004d2c693f4407ed6e4f2cea396aacd11b350a33a93de82c11f527e7cc07967824bf8cc174d4a2fe9d62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1178036afae5da35262b73e2edfebaff93812b6f6e92b8203d846aacf7291130f3f8620e8e6279ee5ca6d3fb8f7b0fd4e446fd29c397e60;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1686e291af70ade1356ad83192bd45428a5c013c7e707ddede90fcf79749bb9750caf5d880fa995620b5d41849de6d833bc03859d1e4b63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcf22a6964e5fca6b5e0aac27c5d8890cbfc617afc5ef6122f4016df73f67cb321f9b83dcce38afcb13d52cc8dce21cdfc284e93d09de75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3b806690762388a6813f99adc889183b9f994da4513540e8672eb5af8138e122dab60df6d849e9ed41061e07e587fdc0e5be212ba2262;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf36de8bfff00b386fe25817f7687a8c5923edde093ceb082e98152f65d65de1287acb3c65ddc25a71cc12b9050769e850ecc9e191f073;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcafdfcea0f8b0643f177e51bf1507ac1c469dd259d229c666453bfa436c5e28fdf597b0d3b15b3ce80adf82de348304c7543a9f1a9ec0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15cad222f98faf5054bf4bfba2e2a12e108fb7e266e2aa76be9e00ff7c4770c001a46ecd3bb15ef6f8ce3bdee6d33bbc4b43fbbac8e6f87;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17526050becf4a82c993f796b93efd63743a05349b39566d9b2639b8b391c714cc4cac3dfdba12a66d0b8297efb6cffebc0c10af0a2751d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1283de8d8bfecab91376ac073c9434fd9cbb6b5b272b68271af97a92693e7be0f881dbddf9b1b8481414127331d1110b19849e6a0822b74;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104c786e0df4380ef4e39f648bb031562b4e160a94b95fd0730bb7028ba939125cc9f1e763fb9c94d1bec37c5a3f0bb27cff93a72567a75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a42a04fb2f940948cd5ee724694f5d6651e0e2c5e376e4b05cd788189bb75db1f242d02a45cfd889275ee0df0594d226223a6e4b02b1da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0120b42d7e4c698202e523dae1e4cd5cbddfeb4700bd457d32cc1b36e638fc8cf7b7670f9d6a5f61fc09acc63988b982bc73811c14650;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d2891404e29f837b28ee7fa3f1769702d428e107d8e70da206d1251ec5db8ee6635b5024247f07bd108bc76e9e57e912314c513671d2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128ef81445e06eee6726bcecb9c7ea4c1009a3eb4c861fc6cfa72d861f594cba7d986ac499589e3484f41b910910296ac22fb98274ec26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180db721ac8a8da2c07595a9bc3bcfb53294a42aa4b76b687f11fd05df9b5c22ef5627f8179e086f0dc06316e71f776e6e988245924e900;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbcc3891f8f438531c4b7398bf131043806cd6af816a60836a0d755fdeb5763184d9698b27fd223edef04136c6a38bad208c0f9a22e83d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f35bd46466d5dd35a76e2d3ecb48049faffefb1dceca9c44654667a6172d61a53c3f52d7c55d38627206ba6df8c26c156d102a6ed4687;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d49d62b54f42a13cc050451a226cdcf956dbbd4abcf98d8453a1b494f3586b058f96935c0e16454811f1c5134a734daad51881d4eaf550;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc593d66be26e7cd407c115a3c99b5d9f6379160e9d9069ffe8a5c0f3625df67f5b4ee2f4c65ff262df28440cd916085d62ede52e298da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1fde7aee7af84757f3992749efe053192378487e6a0ae4fa0521695a0bb18647966197dbce42b9ffe13199ed0aed772f5d1fb639b034e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35b3ff17d3b8485aa57bbbdd8d08772b24f7e2cbde850052dca88bca54e8db06854c1bc531243679c64e3dbc0de3c34ca49339efc698da;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1074df8f53cdaf3ef2455a36cf6d1ac2e7f55b0e74f99f5d85b5139d69415c900df50d7c482c092a09746b91e23c54596d52e33c714dfce;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aa4b7d23bd27c1e5e4ecccf5e34d7c8b068e790ebc19780c818a53e9ae3ce64820dafb0c9b994b709e74e89083f15e9f6224e5b58ad479;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16785e611e3d2bbc6d17372f36ca97a5dd436b99ec43bda596de8d9ae5aa7f93a1737fa746af234ca98f75ae2ecc95d2f87bfbcbd6e177;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbbdbb877f11816a3945ecea8aa7b4b1e9fb214ca94475acb2aa8a5fbfa380805d22499323a8da877e82c55fce070ad5870b7ecda6767ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1041082cffaf716b645ee5745bf884159ec62f1d22d081cbfa1ef656159f007f44c58aca0b4531fb7e3d38cfecabf609bf0a61723b6af67;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c40fdac3d3a14299a0a47af20583dd6278b671682659c72e71214eb67ca13c8d5f929cb1d160141dfd87da04064228a365468a010a6d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1507c0b87eca6fc1faef7bc2790ddd8447e9235bcc74659589c45054d18544651ecf1f505082daa71c087dbd6c3af35cb950ae30ac6256b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf141366e249bc5b555b39a3d074421d184a8959a7b30d23283f773a14f3deeb12951ec4e7c65a1e7c4faed42d4987c043dab7cd95a8399;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe8490e005094a3b00e48d70ed350fff7257c8c3394d7bfe24e6c4494e56a1491c198a9d7e5a264aa7faaeced5e3ae40f624563a4e83bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ccf131629610d0285389bb2e0017d3a0ae031ceb41d908c74292d480c8ea2a64e4e3a371af9d95e7fbd052bbf46a197da02b3ac934d30;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1291f0dfae2a4542a91fb85e11ab08584b6bf55c3d4dddac7444fcccf1105e118a1a116910ba37daae8982728c7d8a6bab2a2b741032602;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ed4457c1cad7da592c0f66f44360c917d2f853744374caf051d23fda385f3c9ffcbd0acc52469ff8b171d4a5202c54b1f76430c32004b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd4385dd279319aeb8f2fac9d7a56a37bb619a16cd305aff6bf882d54cda01e6481b15fd90b01693b2774e5b971deae5a1b458b8de8061;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1149c9e89687bcba2dcc748f688d0a4c4bdb03edabf0ebb4166d8b74f7551f19b83f9044832fc93b3932164b02987149d36ec3082da71d3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c25fdee99f4e46ba07f39bff016483e8ae437346a5c80f14db025da9cde9e0c9e6a08dea22ed22069394d1666caa26f09fe1f4547b02c0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16191cfeffa839b3c2ac89bcdde3ca02b13e82b0eaef121ba6ae74a8586d6bde591455be280beafe8dd0cc39a4ddb3373a791f523b7a490;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ece9b521065c07fde84472209d7cc44c82201136216f6efdf1c1243fcb6ecc5bdd8abea359894fdf379645e50bde0fcce55deebac0776;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17713fd96de20c8e5c479b97fc4a498990aa2aea0652022b808945a0d8a8b52110edaf30b23cec2872aeb6358dd8d78d7608c70c41e610e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb46fdf34ef4a4d6f10a0d90865d5fbd1aac059745531bfe0510755cd2d0e84a0882f7a18906d54cfe7800635a49e2f640e236094e75539;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0258c0d8376b8391e74e5bb51302d97cb18d0cbe3aa811210ad9d3e288991979bbac930a670e6dbca835696e6add7cee0a73dadf72f15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha574c1419ecc80f0d895f3884ace1f0b0c9dbfed59b1e6722a58a9ef739849c07fc74e1863cc9b2499c528f7b4815de0a0e1368f1980e0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9bf0fc3c78f0bcd5ba24e2696ed193747e193a46a64f0e2b56f7aab579db250c854713d57f755bf3e647c62f95effe2dbbeaca568a11b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b96280269c2c60f8c96a8708c75176a3a03c81175f1d609dc37ad88a80fbe986317ebac0362d4723d93be8ca63e10469c10c8ef683198;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad98aeee72e205630f6930611cc2b2970f1807282214dba7b713956b5a5384074e7b06aa7b4d1e00793ba481c886c9723648e6be3e1bc6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13db63276a3c77efd8b80c8e7e2f1f0b4193e1bf2dc983f8958859bbe50c8996fdd1401f80f22b7176b5bc2e6854c54628d8db8a5070985;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d2b569b0785822570da623033b9a7857c776a143bddc0d4ddc0ebe35e01cd81b9ec8d155548f811f23622309c7fba514f7f44c86ba695;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2e79ca2178d95d59e00fbd5b63b05f104d33c4622ac7037dd65719de9ef3f6d16d6c0d37401960f3293da1d0cfe702c97d2cba326f6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h154b710eabb75ab2c7c465eb68ffa6430aca310bfd39f34eb44f9c3364f1f616e06a0ef26b87c32db41c33c80b2a6b1b95b2b77617e6c62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcb5219666bdf9632deea638cd12a841e22508ef2377b9be281392fee001e7ac93d91c9cc186a713f5c2b0bfc0c737a9862ca2bc169882;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79e48aa2004f257745e806feae4e336908dd07697419b94855ebc39443bfffa3b9491ea17f5e4250cbbfafb2aca6947a0981067c046079;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1b9fbe34fd691822be70ef8ccfe87f49eaeebe9a766b5a792bb8ba1e3e48a025ecbe44baa33e372363fdd60ac0448f1c3ca6565288c2f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e0a020b737a15e56c90f862ce7867eb6ad03713a45be10a240fe8af2f6be80ae165ff76ef227f3fe819353ad3f5f8005f2dff5c34a5cd9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5fde90ad6792915d1d9466aac1fbef19d60178dcc924f35c93d997a72642b2bd33afea47865c0ecda48279849f94369e192c4299a91d94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139ce00562ef0cc2fa97786d7fca6e1d4cf08bef8390d8c9fd212c0290d9b61047cd59415c1b99ac0ede44b39b8e2619c88b29b3b83cd2a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13de2e2a446fecb819d6f1c2d6d2b444058e5c1f51ad350fdd07c4de38194e2c9c9c8ad662c262303eea09920f190aa0565621366e7f5b7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bebaf1756d9b962d8e436878aef99f24e4cc0e75bd78111d8b5e65b13c078b3d91b4375a9a1afa137d66e2e8942e2882c09d2f66d2dd7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18648524d4242e73d2dab69a02e371ddea7e800d0854d2f0a9b25493b5353a7233c0765a37b09b3625a341708434903d4b9525ee5ad6c9f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f86e49ff8c048c7e1bb3830f1fce004470c34aa588e85ce6aecfc7ec34b5e1326702253fac8d41b8071cfa3847c41ff4f1435b2aa51c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1360b29b9b814e8f54dddd7a0795a63853f36ed811cc8e1eed043b4fcd6c9b7f1f20ce91490b917dc8e77c5934f93cbf4fdbc80438a2be8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b8dabd4da5d8d107672ea42367066d523f75d4a384ab2575bdaaa3fa8cc3376948fe97d493a1b0856e24a9a0331ca7a4b4d855a29ba48;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa5a5b298760403bf0818fe4735d5e9cb6ae2cf4a9cc506abdcb0c0e6a6fac09f43d38f28a6a53c0e7283926e2176e3cd9450005dd95f1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2409af08c60f7b891c467c85476bf6ff241e3b7cc780ac35c6232fd413d756296e4723f5e9f9672cf4157bb5753962196fa8a66a3661f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb004028af5866528423632be51e367fc62ad323f6fc683e225e06f606f435426a949f03929fdceb16ce45eec8bd19b3cec331de5381965;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a440f6d52e7f52b2069a8b087076fc0d489cfe41e6ae87794429711f0bd47551260836e6edf51ce6ce22103db845b053f3fb49fb7eda2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49c190a231101c69ac519763fbcbf268a90b121c574c84e93df25759ec37ead0e8abaee0865da741848e188a7c545b71011a292ef10aee;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a7c44f7aed758b947d0560d742f5904cc102369a12a77d9e24bdedaf6ddb01bcef1f68452cb8ae298fa6d877d6b28e71083491fa3de63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1539700f95c2d3c08d6d08e8ff26f76ac74aeca5aa16e34c573034bcc0b94ae24158f27f7cbe10927f0ef841e81406e856fbf7ca81ae091;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe05998639bb3317e86cb44f1de196f5554ff1227b0912ba09819288e5f0f6434c1193a7ac701374b237795c37d60cda3b3b3383788ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ab2cef10f48e64dba5289acb5d44f0d076118947513bb62ae178f8c2c98e4acc602427cb6fafdbdabda50217809348379e9263ba8d557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a5a472d07284057712424f4149b60f28657e3ed354b232493adee5f257a60e356494ad1cf9df4661ab30658269f26cc1ec5cb12a0109;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70dce6518214cb8ae1cf8a9ab712820bffd9832f7ef093b839c5d9d7b696fc9f1c58dea8d51ca7d85e1cc2336606edd37c55391601da6f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1efa1fda0b84b4b76f2c26316210794c1bd6170f3ce2e883043a1a4e8cfc6eb8d77f7b85bc9a416e15ea8985642fb3f89637f2b1f95e937;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf9b22a8412925641b10ec407338583178066a04d6c8f0478ccf29006f29e1ba6931abf975e917eae05a39edf0f499b8d743ced9819ef3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fcc9babfd6addf12fad0fac42cae7ec6910a6c2e2bb2813e6d0fa59c7b989dcb5586d9352a1ab0f26cdb3f865817da6418115f8f2b82b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc84abc34cf0f736f63c2c2ca9bf4dda92a5e585d274ccb54ec1d9ec4294b2d9917018600f26ee0a2b1e644ccb9714d7190ad8b4163314;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d9bc86feef7348c278bba5bdf4d0bf2bbace2c3bff53cd12c3c5a803a1c4dbf925ba1ce3ab1b118df255a33bddceb5fc972ae565e505c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hebf417198622a7f235b92705e758e81aa317d5c75cb553b46bc1a13042cff2a9927ffe5c9076d4914848166416748e8e1d3185ba2f53db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb54b2eccdb4a27ce78fd6518cfa7b64f54f43de6aa87f68ccdce10b47c6b662fd2de4aa8edd217c222d993743e8de7a3861a0a2d4acd4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108908435a9dc036e2c170b95764b5887e74783b38d87f3c5237d3def0d2d4111068dc3d4f2a58ca461bfc5a8d4a6bf184d6420fa12eb28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1246ce62afbcf49474ccf1a4a625402532025ec36434576bff7367a257b78f924ee6a49cf3c5938d8412a98873c16f0db3de9427af1a09a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddb8fadb66dfe85bba8488d2a2c20eb378278ac1094ef6166cdf46badf28d431bf8c917a5f63661f5a5d22145ee3569a932cb9d71778c4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11de446f7f970d5429e25987a38d92c61cd12118e0e1768ccad399c75b1aabb32ee72c461de55bce9f2231c97b840148475f4f37e361b72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ec5326fcc12129af7944dc8ce127fbc8255fad67dbd3e0c78d33588aafbaa67921e40ba3052e92c097dbcc15fa49e242e7bbd5454a423;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde29500f7e9a8332f06c1ead724a52a5539f49efdbb745ec5101bc68918ff8a7642372c5207a21045083a9d2237c2a80ff9bbb09d218a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15eee5668316e70de6f0e578d33941545b1f9f80f64cfd1d85d1899f98e57286857e9335978aae748b83ec3b0107b826c7d25a98a80c17f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbb2d9f7fa5e10e397630a38ab4bfb7aba7a0850bd6c684f6ce2c0f3a6d21af2b0e9e407a65d9961941c07be43ac1264d6d3f7f0db20ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1812e5f52e43c5370237e8807bf61654853521440aafecd27b8dcc0f8d3e23cbc5093aff648f17e97fd135bbd994f3f304a7a6f53e87a00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6a3322d8c66fbea7b08db5f90ebf571810cfeb84fcc4bea1764db451e67d1abba400815ae71c9fc64100c2793bd0bdacc098e05be4473;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c948bac82776b82079699230d76caea806b29036c33ba6b28c50160f503a114a13fbda1e54ac999afd144ce982e468e31cd0a5b793e13b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1988447835130344ffcf91e8ad75fe2ff3465f8ec380153cf32458d05b33540ad9c3fbcc97e9e1f0b6f9bfb7a90b538bf6cb375addd28d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58ff9510a74db78cee298207ad483fbc86b09fee635f0e968b6fabde20490ee666cef037d741f7c6159ef49abfe2ead058e1b443d9fd6c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3cefbea65b29fa74c4d4112d6b5b48b57ca1ecd4901dc1d9358a8226bcda33c3ee0c1b78c4babe45ba70626da94f7b3e3542ce9cf6f94;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66a0b0afd084c3b78ea719e33773a3ef18d21bd863d0caecebd288143f8df075dd32254c09d24aee6a30030c2d392ad5e3ac668999b071;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10bc8bf29966f9f5ac8f03ed988c6ddf326907c842048f621f88c9eb9b4456e813aad717c6fc3753ca88263b07e8df2008a51fed8170b5e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2c76ac2be091a7cf17fd1cc2ae76e6c402450bd3e39e0c9b9cf4649f7ac03c46a54fb8aefdcbb6e8a090bc3c69117d6eb28f62e086cbd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99ad659581cd0e798458a2b88d4156e3800f7d8b1b95006f9ae2fad5ca3986a43dd80eecc461b66f8c7ea4068e1b40953ea4d4d8c95b18;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1301237a0d122e22451e4678431cf5a7e8be1a408c59f8139b21ab03b156ba28680322ca8cb7a94c4a0ed51439454f4f18ee8bb26c61776;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he787400ae5bc9314c157ffbee035e726b1ed22066331665168ebab5368f3f04a7771fef1bea4f6e3e99d0522479cf0c8016defd145cd62;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1816b3bf99aaf977795db4752b44476b69a8c4fdc7cf01aec210e3af9e8b43940f042137b3ebb7cebbbdab4c56b7c1c8b418d3ac208419f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h64dd344bbb96ed4db1982a4d65528af43b156d4aec3fcaa7663377add347542149c3cd3a3e20776ec22126b2be03bc3dd6573016a1a552;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179f594be432f1d8a6f38f08b1f739269bbab4fe0856f9f5311d0d4f3b140f2023f67d964941b4ad4db8db9581d5d2353512fd4725721aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee8a4dd1e55e5c01b0224ac3c453d5b43fb0423fdc1500529beab50b9449c0994260039bd1421750b0ad691bb725b55934c84657062f49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cfce60aa5bd905105fc45304008c8b15e6eccf14fb7f395b42abd4ea163e0421371cb3d8cd0e1014f8f63d2e698bd652ef65cd230bcb08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec2fda303652fc0dbc174bdf27529ed0fa99bc5f696923275990d4651985101c4ff5e16bd54f38fee8d50860d913521d7bc33a4c1266ea;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa6cbbef53988f8abb7685ed1eb1b7446679fe8dfba96d5ad308c2301d85d5d64d2bc8693a69cd4e56770dfbc7039ed863ec75134b6cc9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1549bedb0fab773fba61e9d57a33a6b86190a8450c6c6b641b53f534a43db3a151fd4cd00c553d4abccd14c874c32c2d54228978c1f8e6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2b820fa16b7fb5ed27d032ddef4251b49a5ca48e615da8db52b665f9631d44959570a4de7c7dc4febb73daf79339145870d73fe47e57e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2efb47669060bb59e7639062111eb9c76774c0f05bb5aec0167a2895631e9115685e1290d2e046bf6fdfcd4e5b8455dd48916fde80ebab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14caef7d14969985ddc02959887f743ebfdbe257b157d179810642e443496fa369f9c1cd6264c7e930cd74be62cd3f04cd818ae5fe3e4a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8722d9d58b6b1076803ece870d1cdfd01eb695cb8ea99ae9417f0c6f172ec7233923eafe322f6c24b007f6fef5728fedf15b587beb7d52;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b98b66033d9e4acde7abcde7a24ecaa5f63d8b8bb51db7862e074bbdcaebb7784e50372c1f9263ddc3bdcb4e1c71de35808abd098bda7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17796bee754f1dfc93c174aae07d624a7ac4ef2c579a5b686dd7db2c02376736be4c1db83907e9fa69fcbd6dc5eed2b30b63bfe463ea0b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c3325fb431ab0453881d7ebaa689152c0eb7ebfb84d91ecc95d3060f759e0c705ae62e74cd7456dfde3ad8d2e6612cfa3bdde686f67cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f6cee76f4846cfde4266bcecee1bc945053da05f655043d518eedd4b7b5dcd38eec14005c8d022fa47a4441b010bf6cde3ad06a5edee2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58c86aba462565782110a594b653f68a45a31811199a7a14fac7753fc27e34aca48ac4d523fc1bcb256e4dda679037c78755b90d904664;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6951cd0ae0b57febdc834922e40389f0f5f7d88819b20a353cb6313beb7bd3fb79c9834196758a8a90d135b82a34c68a0f7e278c8a4e46;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a250f2505670705977f6a307870d7534af3e48417f2ea9d07095eb4ddb768f6773fe1743184c440576e366b1e1f325badfaa0c4ed924e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be6c2003e73bdab6d8b164b8f56d03c20e9e0765695747c4f0c3dd80b2919b289c7b68bebd7671fa72b85dd035697784e71159850b2edb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8e57a6ea9d7c978772c746f47d0172f9ac3fb3280d3427ecf48110b8752b496cdf76856ea1666bad16dcfa925cad91a4027c8016dcff2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1198314f8c0b7f824015960a5e84788e938d6cf28b35b255ada6b46872248da4c0ffe888f728d67452489c61c8730e4e456506ae4a2493f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2748196a39a175430dc30157fde90182474882162f3d1f807f6049a765a6f24beebfdafa291553e32f862c98a4b24b4619790c5fa4c04;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2bef986b7ae91f7349a528e32b511bd05b759d6eed00c9cd2be903110ae3693995f4bb0f493121fb9bb67075a2cc3e51b36c14077ba0d8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h691d58b4eede542e23bbc7a724c743397bf8844cbe302adaccea2fae2b6631076f99c16a0266b06a48e93359b527921cb6415694102ba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182de3db1be2b9aadad048159ed20bc924119656645f34e7ea2700ec4b4dafb0614a1d8795f3757336537602d8a530fd107ce25367dfe20;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a42f62b3b96bd74abeea3c9d0ee4de455cf8415c88dd7514aaa556bab2a143f660b31a44c0dcb05aab2965efa04e97904607e723a80ad6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5e28fc88c16a9e7346b0fedc1c308259b4a5aef364ad1a97fe46ec87d735a54aaee7902b69b5dfa1a22e836f02231946bb606d1f73ec4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a51e272d335cc1df7789b407fe17f4e45a6317094dfd5f20504043bc146bcf869d0f69e872fcff2b8298198377b734f4fbb54fa70327d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd49d9bd6c32995fd07bdc90580df296cd955fafabbdd43505eeb2eaad2ecb221b0975bf1b685f7633b7796ff58087b87420b2482c7fcd0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd01896083701f5f367b1f765307932a7a95d7c6bcdc79e362b6af9dcf010b54ef67687334f9777b32161b93b692f16263a72f8a022560;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1a1c0bd06054d0a801b4a57db51d459c5c4f20e49c7df31148ed22a111251b42fcb7236e56e9211311201cd94846ccfd8acc051944803;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3ce29ef2fd0090d0ef84b9a7f6db762478a05d4c049781726b60ac61de41d8578de5edccea5a86ec34ed55a3dad7f5bcc0621110c2e17e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194b5561814317577b05baef6bd14eb1a92c782a8bb632a663b432b8b4c79747e9c19f7c7176a5f67c37a0d8fc401b54f5e9d8300c9b59e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fe6636d1e1b572249d0b0e90ec69772c55881eb9ebcd07183500ab747a7a243db43b710998c3387ce627d3c0e8cc9af37f4db59ba14ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h165a44af0e99709743eb10f87433b460776e32ff2e8f4bed6be1660137cd7d2b432971588a3476a6845b0ae41bd374434d00593ceddf1fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91593bfedc9250dbad6bf77eb3780cd576b3a992d18f48e119240f10206148622c0b048c4f48d271be1094ae9de94a8c5e93bfc3b6a5ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1caa1774faa90ef009f240cdc70446b1a35c13ce4301cd780f6b1a05de22f129848942290f24887802e2fea2d78c9a9f4cc4df9b234b228;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175b00315f67aaef8b0531c9aed2a8d203f1f71707bd0f738606c1f959e6822305c9e5f02b367dfec7a3a76ca1950a79172908ea17a221d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112068285c06bfa3e41eee50ac643c2af9f9075e1fd6500b066d569891872c5d1bcfe433ad60723117d38989fc3825c9e54878701b3b2e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d5c66bb4930881e5924702b32dd5eef968d314b22e8aeb733c70925f98b07933cd4029bebd522f4df1e7b32cdf0cf7ab02d7122a10b8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7664fcce814a2690ebf72df0bc00f01adf449af8bb58a391dc978dea3364f094e9d480f275462a771bcf35827b0acdbb21b44382e192f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1066cad2b210a282f6b28d666d5e9573ca2fb846b4ac3c46b153d0502bf1db49de38e79ccd23a7c724365a2cd90d41c3e7216faeb409ec3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h61a8a6bad380a45011cb165135d579b5214909669f9bcd39ebca2ffcb33380dda076c8f5d6ffe95cf0e34f67a44e033c510eba13b0179f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13613c1bea78bccbe479cbd90e2208cae9da94fc48fb033b9e9290275e80299074e1dd55c6fc6a5c3c3ef7fe33c3e738ade982117229b85;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f03b149ad9e62e5e980e39a6dd501757a3633765f2b70c46b02897d66d17cbd4773b0e9afe42a06c4c4f46d7e6b7cad0e46bb61824e307;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc59304566fc622b93ba426a1cab08bf4396429807abd9147ed6b308d442a5386285ec1381349fbf45a1f29e02b0e4c341adadf114a013;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e69ce6965fd40029e50b8731d456877dc7d8a151c4e625e6dcbcb58fc319b14f99cec53ab9d23729ed62eb15b669e42319f166572ae4c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188708207e88b62f07f0702bfce111ecb175132b834ca5172e77d9a0c087fe1cd79434c21739a59876069fde07d18e9be13c80a449eef64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd3bf48352aa1685e417043dc65d40a81749529031a0c3f5b60390ee2f539f760315072876a2764dae0ec9ede8d5e92e8a1bfd9f8d0b9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f443aaab099e5f44c4f453fe80e188adb5cb689d8e29c6a0b56a63ed5ef99c6788e20b8930e92009adbe69590b42b7dfe49e13798c4d0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26291200baf5041a5a78f3fa2c78e8d8a29fedb5b19cb007f412e675de73d366b84c1c093923963fa9292956a1fb8eca72824341f66527;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a45f53fb97c306964f3514af2545179b76f7e5f3880f202533b85cbb790dda390dd40026f12e936c5cb0158f9549b001646673614c3952;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a32b6674ee9970e994de9113f6da3de371d05523d52ff010ad8077da7cdc8ace0291ba1cc40bc68e68d01c669a0da83bdb4bf3164deb6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7aaccce184c301e3798058fe1d83d21367c9b1370530837a3e0eb4b527cfdf4b9e0b27ac89c32ff8b6729547388d586636290ff5be452;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1909ecca585cfd27f6716169c36758b3d7c542ebd74a2759ce5d676e26652ae706e438e34c652a8c2d33463e1ce3b9b99aa63e7d0854212;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h35d9c7793b678c4d0e2e4a8bf12cf07a658cf75ff265f5af755b229978a17888fb9b171366e1be52f3937510828dcdae7ccfed904fdbbe;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb68a69ba8bc3a727414c55b985737ecb7993135fe9e613b7150d9460382a3007f2fc3d3b050c6ce27602fe7313d2e8fe57a077fb86078;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d4aefcd77a9d65c2548a6de6a8beddf0bf4220465cd1ec2deec6e4ba936e71042961ba09742890bbba163b5a8743195e472b0924a05018;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hacdfee969b21740a806c7197a57ea91a4baf478f58b2d9ef04a46856cb71f39922292946c8042be63caa574cc2dbf5aa643b320de24905;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a22b4acc283326913f141791b93fcb601177dab37a170b5cc19962c6c00f6a09610c015ce2fd001452eba9f0ee7c04c813ac7d9471db1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1005d4b363d241be53eb20e85d6b89743a0d7be0cb65e7a7ebfad2c10667da3cd84d274ae2ca5932e907067de36bc277ce1d612b8527512;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcda07511ea4a9d2da75027dc83a67b49799a323050ea37621857cd8b96da0c9f5ed791c93ff938490e8278ad167fcea370a7dcfc263137;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8713805f3ef8291163c0719cc37270004433d8319650d396f982ead77570c7ee60b8a1040d181970d279a1e47c4b1b7504e617d933b7a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155a6738cf07c4a52520a33d641398d8bf78ab4c9f41ae45b4bb75277c7a9b5f543db446ed22b58dab16d5b04f310376d3662cda0ba971e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff169f9878dd329251c09752bf3a322cdbed5f1eb4048ce0334bc8b58379ccede5e5d2f732f40a0523a99d48fd9c2c7f08360d71b88c86;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d4b2b11397ccb911b3c1c7fdf350ccc1377bb03bd854a42d1c6817b6aa0feac195813b81c1926ece5b26ee6e82bbb96fd63e59abdfe047;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151236f10c4cce4524ccc9b2d8d17e7495a90fbbca363bfaf0edbbd094f2e9118f15e9e1f00b0aa25fdffe33287e700d765446ebd43133f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef7278357616557d265f429e6f18e7fe42ca64c352e40b406e4d9b9d650ea835769d9a44c40277abfd2558f27c34a5753f2f1cd372b4d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65cc8ada46cf9f66e88c7a35cdd9340b8589f7adf3bacc40b5f1ec037f3325ef8d37d7c4df761874dc202e7c026710a67ab650163e0ae8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e8e41bb49795fa77a00059a4d2c3fb0b9579d739305be10d302554586c51230048655cdd6111ffd5e35fc2b667320d55cd230f833877f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a468cef12a585dff6c9557f65ea21f28f7025e602d5733f599656b2caf9c6588ea7b4f0bf702d3d877ace951f40c182d718ed04e9c7cc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188d712e5b6e027325271d274b400049b64bce1ade1f905409d3751f1c3284dbe11013f2fef044aa8dfbf8763aa8bf644af919e30451d3a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5dad94837b1f510b8a700d52a625b4983a01ee3fad615188199f32ab37378c064d14c696865e8b501e32abf6dc3bd6acc6f19dc673616a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d3b5ee0b0699e4b0aa111108cb631dda7e8b42272adaf9de7d8e2448a83337cd7b87560e2eaa5798146d647f98b3ea69a61381f3bbc65;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81d57b7c957b1a72470450f5182256562e6f97a9df3ffbd15bbe324e70ef104cae443f50804aa01fadbf53ae599744c5a4558e0129c6b5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8fdfe1b0ccc822e1849e5495a29a452f8ca0324534b96bbbbdf602b856f8254904c1201f8f7e853f2247974cd2b74ff4830f272ad296d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha357e1f4a2e2941e5de52ecce557e8aab5add608201e1318fa768c6380dbaa3e0e58490e62e4c8d077c584e750ae7c366c15c79a7fb40e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2dfd975e5ca8f133f5e7a6217a6b7e9d7e31e2e572329093a980a24aea59bc381f5466c9b6affae799154ec8a96df25fd511137edbc093;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178ed275d8efa53cae24fd418c6a8eece455022845a92d947d17ec434c184885c6b66e78306f7d9d6073040f67cf736100c7327724c2ce1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcab855850dc0df8626dbb5d5ae96489f286dc404e16e8ac94e37ec625742a7357e68eb167a85dae46b34998434518bc248f106fcfd746e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18cb6f884d459171746afb82219316605b9f3c670b0211bb7973a75655c635459dd8ece54db7835c24f09b4bc1a632132adb4995fe6c5f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h281504ec5991716fd213e956931075a8884326271a46a860067e384200f497c377efaf39459cd74a76fc8bf7e47d3e966d5d6eb3154dcb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h174dc9240288a731a51238fe0d9d68a86a1e46d0eb261db5e2f9d95a86e5d792ff75a362e27e2e382829a6c93cd27732616306d9517ebff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1046a97c547cd2705a8bdd1af132c1d14b0b0b69eff63b4d410094cb36819f121ace67f365dddd7082cd8535de45dcfe96f84417ee78f6e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdb0565f4d00e81f4c378ea151412dec2dc7be6d96cf841ec4a101e398f3fa79372b0abad051583b401cfc3e9f68dfeac5cc51795dc9f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b33220bc358831109fee898a2f3fe6700df42f16870fa1c0617ca34130fe04df291b67b59573dd363380f9b680b41668ca663aacadbe2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h813ccf061aa0244e83f47a61f708eaf18c83f0e70cc7dafb664e0606156bddd7657c60ec91bda9ccae4fe7d6040b62d3b057a393b3acf7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9ca928b0c5e61bf177b15bd9e8dfbb777e2fa25a140d04d1df3b33b13dc01c7370068ac50379048cd04ccd8caa8fade5e1a0edb572216;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h640d5b39c50fe19793fd5993723cf162c47740f0963c5ad0c4cbec5ab49af29f539f467cc66e8671e45a0ca1a97e403580a20a70c047ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he589c5c1663a0e34b9a9c6b2f48eb61d67363e6668c7b8a6e9ab71f4d56b1673538827769638fe44944ac5216bdafb93d079f16a01fd17;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15731024529b5b00716669af81db0decb6278314e6c30c1862df88d27915d784122c94c627bc67522d34bcf65428c33314c48a08a12afd0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haffcef80ade4855ed8e8745cac0f7bf72b5c96d98565eab53732df608be289d28f2708d90f26a0c55c71178970233137f1386f3fc706db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h604e6c25249d14245a685452d440e5252816f1c1a741f05aca8d660d4311eadeccebc81ce085e9ae710c6185a7f067317222620bfecb6b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3be025a4effe54c11abb2187667024b8753483e6e0c422ac645683fb5e9726cb99097a0573d3423c1a3093828c8e186319f47ddd2377ec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d3d3bad2cf7425aa3d24c089ef785b1591dc5614b712cf55cb2b91c3718c32caf0ee231a6c5476d885a68dae8bbd29a35bb194bbfc84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114adb7e7af9d42aed6bc1730d5494425abfefdbf89e2d38ffc8544340d8e8675505b01e0c05df04783e81f3f79809cb2a5339d768b5e7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h170f7b731467eab60846b9666f6157705458b048fb6135324ffa673d8b083a2a8715cb276bd1321bb898d749a1dcf9a831f01344c813215;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137f53ea15ce6daee6645e7e8c057e4d2ab59f98e2426658b4a92721b226f7352dd2f7aa922186eb141ad132ac5be91e55d40b291b89084;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4afb2e87f046e9190821b5aae20d8a17e61813e4841fc2653e86aa9a4e072c1e2287afeac1ab70a348a932817301fa8ecb0987433c15e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c9a5a784477b5070f9d4218547ae21d5b40105e6b2d0c075b974257bfdb3a1c25b69ed64eb2c4f3251f4b9840bd975d8ac9797f3ab038;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b9867b2cde3cbbe184165ad078ed7faba3e6adfb33e97ca5bb28c7e47e4df2621861db496699dd0e5da6bc9d3fdb92715e477d87c077a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h154d66ddd65376c7c5396e5c691c0f1d45c4824dd57ca3260399538b9db2db37f32ad4badea8d602b060a9d36e561122ded1288c4a79650;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7fc5b8f6d752a146896bf57e0418c036d026fc933c2c189f7fab4e4a8aec5d973e2f7c17e79c0a35bd99b1cd5e6bec8028cbc3c4a7255;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdaeb8a1be48fd9ef177cab54f39a8a8b1338b014612dc64b5a291fa0cdf2ebf85207899adcf92b3fc2bf2bf405d46a355f92544d68a9a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h184ce4041d52c750c7631eb5a3351043d56d7b2fd3583cfc1aca081d1bf77acad61056dd044943c7271b7fee7e43dddbb5bc1061d77a945;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadb57636b7e245019718889ebe9cda41f30afa10c874481de7b27abe758a90fdf9894bec9314e96a4484621433950ac9a5908983942ea2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1389ce72193f5f63d5df440b5c11fcbf6c9f523cf549588f516dcb8051f4b4f74bba2dec1e3b1bc7e3eb8dfb6fe1677eae95d1f951ba085;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d528c6a3be069a5b38fc14997811035b0239d9ae39f80db77e2c69a57ff7be7ebafffd0c10c688a5c6d93d1a71de8aa362a838fe85eb2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7f42bb1816f79ca835c78d60f6dea1008e87b5f586621d8c3e6f3f302271e92b9abbe0de09d5f2c827bf51f7df0b63f724261ec858eaf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71e3d2a8b8ee67ef90473a40f16a071cf21ef1d8cc521e2630c2fa76e56319f10a19e0b00ae3aa72631a88d5a39d35a2365a887a25e820;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179c6478177f9aff9b4393e4b30873afd6242db01ae43025bd5874caeae5e5600c36aac6981c1a5c47e9b2c7ca0e6e8bfac380090b750ef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f6994f87975b4f6e7cf982f878d4ecdfa9f2498dbd8df10688f1cd8fc314b1ae01c80db78da6a7b423389e67b92ab40f8dae58d6c58c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5da98b10513033ba479c4e554ab0943d884d5ab9b0fb8995b3a5985be5df9114cf90da9072cc31f2322b3e44a6bce8e8de67d6dad2d932;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9676932ac074673c1e898618d8244dcd5d78aa65f980882c7967402f3678ebd376c7c3b714a08a1a1832e8bad922665aebe84cd4b8521;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47716d65f6b1dc847f741d9189731f1ff3906301f6b8df0984fcfe615624cd18c8184b0edc2d2837a7099604f5f27ed0d635bd872ea05f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc334a365b6c77ff4a350f6a38aeb7bd5cf604e60bc894a83ce67171bb1665d145f8dc05b2513b78d894144cd496f8906a8970cbc788157;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b2f384e939fa6e1f778760bf0a9fd1d64c0e5d6cdcef636a537a26e12487d910281f21b46cd98b4fb67069586d53ad50f896996a5e328;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b430aa990ea65178626a82c94967d1b8d8ec7e856f221158334875c769e4abc70f3b3f080c01f879ab89231684e6d77e0c9495b93229d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140f1f1a540926ce1459c7c6fc9bdb56d2ed5a75bec30296c3c3f02023f7df148302bec6e3297ca0472c08ccd52ff25de388cf5377fb123;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h204ebd8419057fe2860bc78c8e29ef9e842cadcc105982575a83aca828465a5dec185f057f7871d7059578398a08527710686cd5004ab6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98e7496beef6c5750cfb523a2d2c8825a9229caf032d60a60942b6152c0161eeab502e4e9a540723a652fd6626f63509fbdf0fac9d88c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h585be71b5c8def908242402ab60adc45ef40d29959d62a8af5c2a1da654f57091a596e52924bab91dfb50ae832d01d153c054c4484c925;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd371fb21f93ffda5ba5b6b850537f247f479804dd59f50cbc21f0101c3c51979a9da2f439669cacd804c09f3ab71267a24005d6e468010;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2e7984ad10a81f38534b0bdce099a81e882f4ffe9a28b8ce299ef4acef16898e90f802e2cd0b9ca0c810ee4c11c9f8e78cf8aa08850a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16004f875c6f277b03c33d4d689efadaad8799797eb032cc0271e3341be3db3e7b7bd74c1de3b6d2ca9f82b7177570ca7a116a34e9cfaa4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bbe50cb1fe3be479a97569d4a7f9f2dd744473fac3ea15ceed8653e293eab31939e4e87ad481acdd71787b326b51f4f14eb4c459f58d4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0656611832297f597557fc10d7bb239a32a56992edb3f82f932ce80091a592012d51da199de28d4f3f12f9b1f20bd96197f29ceee2f8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd149bc46edd00f9365aa55053c0cf97fca1a117f7975dd2d7c225a072bfab21b29733f03ad90980786e2d7e26175ef318e4e74fc9021fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3030db9819a4b71b8226a3f1640ab505ead5cca4c77adbbcc69014e68d1910e4876ea5e5c1354f498a0b9f6823b60d5bf793faa17b3f49;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f67047c4f48678dff27109e4dcd3258e3d0ae6fc3b5de26e6889815f8de82d7279a4568c0a166575cf12caa9097061226378e50f900260;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163090afd1ef82231528fa59ee058086da53f6e0dac0a25329c869c100adda266f844f7d9c3abc81ecb0847597f2a91a5a2eac23c345ae9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ed953c71ae4e56dfc79f34f587a4fe33ab4ca5db95c3d1c698b7ba252bf13835950304cab0afc76fce10c22df2897d0c19978e82f47939;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb58e6ac567919e2b11062b31bec4bc92dce3f92560af754b95d74c89038ea858bdca5a91ea9904c1bf7ea6a1a70002f3103fe4f630800;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e2bcef3af342487a998bf6d94662bd66fd7533b4eea496d98b19d25a56bea25293b754467f115180800284f275fd2234a24b69f2bd061;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad20222a21fcf5999116a41966c4a21482e70836f163c7cd7c08bca16de35f01166f6e95776df6a4cefa855737aa46bbd6cc3eeb499451;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75bf9424b841e94a396a62315f1f1563018ef203c9d091380986a880042198894092698e719472bb2677127ba57c400cbff97a11982f53;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2225f070204dd25108591265b0e201e579d8b8f15c3dbd3588ac49cb8adcd905ad403868f9bec6a2d0e2b45c4e288f14e7046033ff895;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3d3be95d4971a67ce245f963106322b6c421709d798d7898c4bc79691e009d043e00f7478ea2ffb3b295b6049f8d297869158167e4625c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9d8025fdff498d622fa9958b97343cbf64bf6c9624a340aaa3d5dd557939e246da55aa5eb429d8f430c8e7136703f9b5ac860e4ba294d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha800fc80ea17e078d8766911b877b65425b1d49c73224ad59e2e7a2a52d91887e4dbd43e991281589b89724eeba28df228eafef46f3247;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b780b2bc984cf13bbe931e89c4736e5fb19235598dc6d9ba751db77dc2ab86adfe45df066fe4aeba832209b7bc2888168c1d7b53850808;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cc94e2781a5fc03649570e0a68ccbd6ce8444804d1db0ef2e42756f820a44a2de7eb7688a17fd8b3ababd4a790c0f78815bc8ab353a28;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26e3f84dbe9d2f72886790f49c8626f5bf1dd67123ad7de76df8e1433a76f285c93ab30702251ff74c3ec1f460dc0d18f1810e14b2fee0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h656b7f98a767e6808efe19aafcf4e60c3c63ce3e6ffe52bb5b353b5026a8d7fb9eee518dd5dd0eae67b9e20d795a982874f8c8ac58e899;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe4a9ec6c6747f1b1b20f584a0a8f9afcc6c4f8f6c267da8bf488a8bc37cb1dcbb359b67eb77a5d7c362a44f4404ea3bcd6dac232a5578;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4feca2f010308e2b078e12dfdd4eafd225112b9daf639777c405ce168149b45c8b8469cb13aa17cc89381629a49ba2042f32249f4cd29;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1000abdd48aa35e517ca060f1663e9c8409e0c7cd47ea3c2f375a9b73d66df3262e94971827926a8ec43115fb3607ee10f8e19a0e8be7a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd077e1800baf403ce6673e734c17b7a0c2fa47f4af40c8b09737ccdac7460e9bcf210e502d4302b06345e6da995090f771f9f1433f732;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ca68b3327369334ad471d8fec80ff7c51741ead50a148a12ea32f658eaec11b3a32bdb15282cf91254525cbece9df79bb20869bf6d6c1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he93f2724ca3800a8fa033be0452a8ebb9d704ea0a790cecb5c5621612bbe4fb0b53efe277ed88ee60452f3b7198773e6de3ca3e6ac6ba5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a96dcd930e611fef1b2be071c0717a775a5c33c3f96c71196c0ae1f74645551290e79e3625e0c43c98eb58fb0031a69f7f1f5fc55d808;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1186438cef64c51ac6a36bac0cff5526dfc370f766db2b679eced25f5baa549eccb9ac9781a30deefb47a4fd853f1ce6cf0cc603c60f088;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3546922554a76ad27b23c6493509f3208d357b14c8bdf7d7582e8d599488c42cf4fcec58faf01778da4fec6ab604b8132b95f488d810d9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0b7f10cb0bbf47194bf351a651f4fda2d1a461609caa8f72a1704239f33c129a4b62fe6eeecbd413d66f3f01cc8e0751a1fa7bd861125;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d85753a548bce6b989bd904305803434fbe55aeb2210337009dfb173df47c089f3e7a9e8944511b793c46cd9c0f6d11a8c7247383ac7e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1639e70c689ad2d4ffb2674b78e0bac99bfa79c2491423bf4d194b3b8a43045d453decc90839b7da577d9d98e836c8846e93405f569c08d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139d5f2787ccef8f92d48a3e7cc2ebfbbf860f6f6cc199b523b65d2db9f0139cd76842e48013640623f19e4d5a98ec49b4c2c4394e9c80c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fafbb4b04110994a84a4b02f7a56c05e9fd9fc0a970f253387cda232fb3df67e979108857e71f31b2084b25ed984b568ad0bb374fd4b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb8cd1fdad297161e24e9130bf4ce67797623ad2fac83c1b9b2d23af12c7938ae7fd92f0544e7a5f39470cd58a1cceccbabe7f15cbe09d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db8b8070a84a6f716a7a496a51276c87236131f89f536d412388f8edf3a1cdbb11e46460ca6816a03b71b7c483484b689287caffb90bcc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19367bb1e23c6effe88504372fe2b01f5c3cfe5818a588058a0e9da66385327aae410f4ce852732ec973c03e4e228a75af0eeb9281a9105;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a119efdbe259373177043cdcf32468ae67909ee2bb2b5cac4a376a6c249e304e1791edeb5c8f2dd86eed613fcb2312e2d4817856ab6776;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3de532a272bcc90c563462345f085b3328212256a33e0a48de0cf27312334e1a42dd1de3acf6c2e3f5fcc308f1e1bd4e9fbd6e8122ff9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb57255b9cbb509524c9045bd54e6252ec6129602da79d4ca5dc8930b25ec80466fe14077217b966e700e5b0dae728803864e19e8bb077a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3cc138424fc287ca5293a90c188bdcb31d7edcf91f543f61158d76db1bd9fecb87acb2ed6c2a57f9f2736a03bf62b533c8a7b6e262361;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c57ddd31cbd383d48d084908a9750d7c27afe4500aeb87ff026fe6f4744059afb39f80a0fec44aebc7f7db6e22893b52319464d57ad0b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac8a98c6dfa33156e7a3c702365eb7aff337b7a403eb938ca40040661e79bb512eae38120995cb8159b9cb5e5705daf8384fcbd6b1be30;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ba07ede473cb09d101f441c6c18196963b3ec710f731708ebe88e2731b198835e51d8af4da892f84d9a9b40389ece142c7adae311d04b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d97d73beeb6422b2e368b1a7a13dd3a67fd42db7746eb22b41c86381560803b4b8bb82374f19eaf812aa17972c74791ea311d1ffb6316;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1698e2c9804d1ab09d91ba0caa0665c70dca1a24476ef42839b1685661ed86d07333bbeeab49ce47fa82988cb7020ff41bec03759df8e95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15c5ef8bf6694396cea8721d4051e9c6837daecf9d3c8666d46d647714a9e597b9e81e80575838d35143ee3fc0c61153351c40a2659c7a0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d969d76d213d38b4bfc257de9630e3a2dacd36d81bc98a5c884c1ac8dce91c4c9e9dbcb9a461d6ef24e2b4bc0e193dff99045d9b5641f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9e5f747e19ec1d6c912eb136490d90d2a15fe696b16fb3ec6884feaf80c9cb5de8136be22ed59e1cbf4ec0473d390c0366643f84498f8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b91db67499714651d460a5d129fcb61751ae82e0f42fcb059b50c3b16975a0da897649a29a31e00901f0554ac85d637e8424a9915ece2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbcc4ecf41109825733c56011ad0a3f1d7f451bfa9b698244e1f330eca9c7d951ef7a51b821b90ca036fbfc35bb72e0985723e4a3c766c5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b74978d98578795bc379e848ba811d822b4662256966b1c3336ee1af956e3806beb8b50d34faf0e2fd039bcea671c6b08a8a0ad85a910;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152c4da8b0ee61856a81a443a812c10bcf2fd678d50c490e3d920265e33315a5c25c14e68ba49231f94f3535222b6bca41842b700e95b25;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3492ff867938288cdb05b9c5119050c8578a9e25cdfd231432fa314dcfa4f54496c0bee48f1780b0be523d5acc2fdd85aae447864de4e7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef29ecfc377400e268a83abf27c3c6a64b7e5bd32013edd8605fa114531d36cc90a8ad7cff10238fdcb93ce695b6c342d8d1988c5c8c6d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h498b977700af4a0a78e1b8c257d5d9186d0361696e9908e903c64a1e1afeecf1aeef265d1be6e7210679f4781fdd67ef0c8817c6251d5a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c94c6a05319ef0a81d8af68736456c232e5cd4c83d38e9b7f2afa3ab7d6402a53a641ab85bb17d0740523ba38f07f59c09e1a4e99be9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58a9cec99ff45f93f2cc08cc1bf887018a5db2fc3c81f9086b96c74c6dbc22ca1fe50fe7e8294307469d942d9b55f8ad44bb242af985b9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h786cad6e5f56c37d382de8c2556432159d72f51815a75ce730d46b2e216025d6c5386e58f243819245597cc56b9dc76e96b7be24f9e7fb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8c7fd338ee75c2195490e841fb7bdbb146822d448f82941ff5d91da1c8a72555dc9847972c2e8c36a3e572d90bd415f775b98cadc6f47;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e0f284c1c9aad4d727ee352dcad32c2984c2b63ff4968595afb8d2789a1cfdcf877654dc9a8c03609aa084d9e80cfa9b18a867fb5ec01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha16b92e6d03fb46bfce621bc54228d0adf70904ad00f9d567aa35ac24b6a8706664435bb9f31a22125bc3398f0f5ad3747f1b00860c32d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e35991632c4b55010c0dcc7c493adca714348b91f9d86c22e3a5cba16eba38cef1837839b72e4e204185bb89e02d2cc1840e88241675a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ad3c0d6fdbc552e631f573ec5ada8fcfa4d495dc8177ccbbbf75dfcd7ef0854ad9c9d0f49a87c8c375b71e803c92463e8ebdf7f002a6f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca1636d6d6a93b3cd8bb66d7818ab967b738ed3b37ddc109e5631514d216e0157ed6e8df0d97c69a6d915534f01eda2ca163d926dac517;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb485700dcac9eb339a0a81d6a1fb92f6b576a580fa8b62f408cf54edb5c8dd05406c05c099f57da4897a0fb31550a30d354b647ef99527;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a41df0b1abf7751feea7534223fb3df050734ee56b9d8cc05bbe9a2a6d6674671e0307ac17025bb85f7b4f2b4fa734675236048c55314e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47d41bdf6900834f388cabab51cc53621657a89f81e97dedd8261da31d2c3c3616682c42f4a24b0643bf9259fa34b7f72b708da1f2c136;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e167d7fa9019b07fb8aca9da47613db0016d95d41f7078cbbc6ef1bae4f94495532d4e6b59fdddc9744ad7cb2e2bb9eba1c2e00e9374ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b24b9edaadbb9cd2cba57018b50b9311289705cfc4c2b8a667bd142a0fe628524cfcf63a6d6f7180a9438a6d8773ceb7424a86487d978e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9cb6448c383104ecdcb902d80907d8c9e8598d066ace5d6e3805bcc3cf190511eb5db3e8b9ad1b8630c00a441f14612a8f250004e66c2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h269451a06a599799349513f06e2aad1dab3d686e2f5deeba2910324dbc0029374e9551b84092473b1343f015443e94bd1081197303b077;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b420b84da94abf11bb505ffe547728bce7bb562bbd039688a19d0ec5691afa3f865827ef99f872b72f5dfa6277e182c9286710cdbe454f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf39dce73dedd23ac0e343f652d8fa9d3d016f0d74f79f60f81b7431976a02eac266d95816bd39be566616ea198fca5a4dd4ea3a96c3bf6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3de114b23d765009a2c6ad91d71bcacd7b4f9bc06076afcba3dfccaeee9a066bbdee1d062b54dfda2db98b16807c1df934b51d656d352;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199e7389c2a8f6670292f974d74fee471624554157de2d36179cf2055d32e1dda15a1b36d982abc6d7625d660b093de7ea3e0019dd2cc7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ad5592b224eb327799954c6f183e4d135a0cfd72329319e304ceb460aca37b52a36b7335abbaaa4a1884ebf190709d4afacc6b2cd408d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff2b26ab5eb610c028b0437eeb1dabd4b202df027f0366511e5c268ff9087c78ede268589dac93dbb34f31cc9fbc25677810635362918e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13efb3e957dd590df5219803fd4b4c1985b94befc0e2e32f963bd1c33215dec2d2f850668d7eb03488090b5af822f1196d9bd02adbf6a64;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c5abba3a70b6feff8f7c4234b75ccbdb4c5844326d85c2f915972222a54a10adb0716c21d086be117af7370b5c577405cffdd7d2a9fdaa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106454d6fd442d85736b9a4e10e26be83bd42ea4f26f197bcb1cfb0e80a79f5db8a77cba2d42676e1f3cde53474baaea03cb8838dc1c3d5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc075f73a59a46fc29a179e5d3ba2833681476284a1480f530abc9d51c87034c507bdbecfecd21998c2766ca27b24d46502dddbcc04a8f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17f0debee1dd1c511fa40548f75394c292a9680b1963c93aa9ec9a27c2d50a38867a4660abf22cb4343bed5661eeaa569ff5fbcbd35260a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1696b7938d6272d6f2bdd4b3ba485f93d2e08c8a4d34f6aedc0aa6a2ee3145771f66b275ed3bec5b7f662e5c3cdb91a9fc86775df17605e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17935b5e4b08b3d23702804e4fc61fc16d2997e9242ebae19905bcb9e80ae52d6a3b64219e1647a952a5bcf5c896455d54f1a9c864f7da0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0fe558cbb07a0a64ff99065aa14b81dbec5652077be56b2bba2e519e15c7f0b880bdace4c674d21cfbf00ec59492edeb130fe28e5679f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3df52de878c65649c1cc80746313877f31ae22bac3b49123f88db65fcfe891ef9269ce12977c6957903d28a2ed9cfe589b9c5c194178f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he639cd9e5ce52256c74f98812f4c44e4b587dbad7d4ce47fa15811dc8a52a41063bde03ed84d381e5ae99eec8b2e7ebf09f4ff8c6e5ca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea24b8f2097e7eec7f62a821c70110351b865d8eaea440bf2f5dc1313d1c860c40a5eb366c59c00fca227bab8bbe54ea96183d8d07ea4a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afb732255335a8358dfdf93642ad799ef5c0a123e821ddb6f07f461dd186b7ae6c460a2a76166e0cf06934f7d7e16f8b11bcbaee8cb62e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161fbdeb7d14326f547a6b0ceee018252c7660276dbf0d220e98c0cc138405cb1663c6d4f30cd879c195f9d98d81d39c21ee163f887bbfa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d09e6a0fb717a5a2d39e294a600cb9b57faba4cb7f19e850bc2779ff24ad3668f722aab57be88df619b4de6092e8c56497208ba5dc2de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63ca0be4f1e2d8c0c6cae59d5ae1c8ee5ae3694c4af6abdd84e289dbeecb3af93a7fb977931fa8ea13143d103047ca2570019616459e7d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1578c92ee3da89075e0d9a8bf6d37e51a163eba8c5f671214c0498047ce7476981705a2abdf22aa7a0fefa2c81d7beba846d38b39c546cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h176bfbdc11377b9b6e84806428a17daaa91204de4c370f71c7de85e9b56071257fcd64d89860cef30e5097be5acbae35c51dc8cbed136d0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1457c12377c15619bfde70725c6b9c2dfc6824f4f6a7b664cea9ed4545fc7b6fcec0fcb736d74b98d571cda716aaa9cc313533fde1cabf7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6b176df9faeac40ce4cd442337bb1654554c848f4255f68e73f211f311c5b4e6e68737a223610b43081c85c4284834b83a1d1d0912dbb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had799ce089f6885df4700d919859f4ada08807b9c47875678ade72f17b9947466d3b0b98ba26cbfcfc133c91815891cd0dad5b5e8e3ccf;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f394502e0b151b98bcffbf6ba6ad174671124648a0dfdd4b3ffb7456f15db6f5bae32ed9e55580d5e08e6da3d5dad13b54e370630114a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf76e52168de15af45d041ac72548087ddd5538ba7795548a4a3e254b49b334eaad1274e6ddce8c435d510d672d0d50fe47efa17b97d0a9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71c9f1484b8566fdcb6114ef87bf65d4bfd6b8296475e4ebe0382d94c42b81fe671fd8f2ed166142778243936afab75d8da2cc542fe729;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f34c7bfd7ea0cd7ee36f45ad6fb8e4b04ecf7bd1b36f6d057051d5b8ec1fe9d14011c2b3a0741cdab686dfde7827330752f4f992243f3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb94ffb86f11b8fcca3d4a2cc9e99cd77ac02ccffbcd5806fc28d29cc398c6f7cf2c8e7111d9ce778f58389cbc95fe36db6a7d68570cf0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc79215b12706fddde8f5bad7f434e2f55bbc532d2328883035f8edba75d5241f282bbebdaf85d512e6b6ac0d9d1bb08cf1540d02f94a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11846895af3615cd417d592722d3b7099fcddd9534c91a1fab51885838c0645d23c07117187e8953610337c1329a7ec942b5dcf14ee3086;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea5ef5177b1aa6c81a71f36e7fcdb51a4a2b7b2cf731ff2c90f98f215caead5ac390af7720b38cb2f8677326a14561f0316b85c890e96e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3e004b7c2993db3b18b22072e1f38079d1f89a1cc590ee3a61450d0ab32377fb9707e67b88d782b9788851fb0ee878de2bb6355e370e08;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fce2f1d541a000c318f5444390e375fc320b8f0d4d6d22579c425b69f860e500855e5553a0a936e98d2f52e7990279659ebcc51e23557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1f50a83d5f9fb4235ca274674b9bb4a4e60452fac61faa93a9c116946f0fc6a9e245306b5b07bc8b687029fe107e7442b4b066a240cf5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d01415d55ed7a98256d31f120723813d83592ad6f543b17591dad053ee97f4faf586c4f460b61fc6032ab1040da2fe5d2c2f2a985eca3e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e0530fa242eeb1f378d4029323571fdbd9e985eeea02bb590f9f057a8c74d2bae390a47f4bfac7555390724054c23ecc94cd1ac2abd15;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ad7b1b10d03729cc8963014c548dadece201a0e51ea7f2c645c1fbda374120691a81719d63bd74c1f78573e2544c137dd26b9e05c1209;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd62486699543012a10d9288bfecb3f629e602452072adc07d72cedbe224a8aed8ad72c914c5b4c795b2b655a5ada1fcfa309aec0437fc1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1fdc2ae8944a4de89d7e9902e88ab634495b522a7f9d1867060531217667743b3a3a12490edf79c41bfdc764ac2ba3704714b76c9bee9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1389e93214b06a8575b32f4c74998081a48e001c42c26f81bae6a0d5b88ea05f7f50a58fb454d33ee25cd78c766ebc8d0dc544782787e5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h706908cba99889745cf3096a57ac6164b125ba02d3f5e151f376b9c3d15f9032c0bb9d9eeea578abc4bf077875fc035d1ddeb10d75245d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h835d5fef3637e2a3c387b94f20ec2b8de25e8e54a30f10960c4596c3571030cae2a5b85458098a815f7f1d916df608f45dc9baf047b859;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157274750c4bedd240f230447a79469522a5066eebc8739b0a10653ac367df52ddca16e0723dcea0ed61fbb2636a1066a87d61cb4a6b4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha6833f86dcc86eab14a79b914c6116be5f3d0cfc4fab0bc94446573b7def236238e1c9525d54c771bc52aef199c6bbbef35b3a323efcc0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127777c86cebf9576d3d5d28fa86768bc65b3c3eb8fc3b3ff671f05f433144477f4e374613d4378582add5f7ab7cf63ccf9951143ce11de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a71527d544828ce1ebdd41615a2e9bce8b04ab949a4750e486863233c893f1f5634384e048a4c7cc7702271c25f807275bede2037f12;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1816197d9cc25743fd91485c2400d4491e4271334235ab8288171d4ed80322454394cf5614f4aced92b46459fb7a79a4705d58a487fc1f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194830785c72b6d39c88783331644b7db9f60635867501611d0a079cf4c18b729fea0d7201d91e2f4593a81c72ac3f35d9bd4ebf8f2b874;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43f2f76cb9d5e319c4acd8d5aa022d4d4a19bc26f053c8397724119dbbf05c6046ef664181b29f2a72432e210839deac056f059b118e98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec152644f55e6e6974e451311da206ff1efcef24f8ab26d878c043902559d1799d6b3cb11f601adc784af9a45cda3a9b5f43d91f922f9d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2eb35bbe5692176cbc6f02541d643c35e8c55e62204e1448a1b7c5ea73796e2215c0740252efceaaf1099fcbbecdcd636f149484a5cca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b7514574c3cc30fa98e8f4fc6a789e6ad97c30ce2a569cabf0d5ca6c022671ed96719479f00efea875a84234b5aba5277863000413fc4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49fa67d2305f94898058318fa0fc0d69b04778c7ed9104a5be05709fb5cfe04f76c0d62f47ba9ccd37d269eea149f586861b30998929f5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb6f736f47f1ab208a567fc800862caca3b994ffd7a7899b5e538251973fc524ab1932197673034c1eec87443e2aa2da3f80f9fa7cf5f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ac897dd3d175e88cbb708f3b6f8a364a45a0ebcfc2671db7da8178ec55f6bfa4dd96661db2ee0fad7572de91f0ff5c25b973c819ed063;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27c1f7cd374090485dc784b75d17f22a895c0c631c1c1d16a9de02cdb636573c8539dc26d22a43ce5f2057e153dc4b0656fe3f53106287;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1574fe6adc40c281675a5902bd9bb8d878540cedb90ffcc04a3db0b38389baf287e5791adfe4914d998fdc3760aba9dc68093de1b89e37f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129c6c6e6a6a7512eba4ee536b7e1ed0a0a97726e30064cbf3a07050d5ce616ab211c878dd42e29d5f035d595cb80737ffc25c3f16a0c4d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d62c3790da0dd8b07416c96e7d7dcfd99489f15bf951138b393d8204c48d6e578f475cae6cb35507827eb20bccefc648b85471aff3fd0a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af564825734cd81a424757c566bccf483ea5e38ef97f2f880103d0ae187eec1667b3c2ff64e98387254a95252e02ca274aceff067cc484;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d867dad3ec20554d8456790b879e8db52e7b1e80feeec22500cefa9cac961a9ca2194a379c21f6616e60f42cc44d57abfa3b4d0135765;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d4403ad55aeba46d3f4a3ddef596ed3b5aa622c8c4fd9188c13fd7a4cedb97f9a460ecfaf280ab1a7cdb2f064348c9349b615521bb02e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f9fcb46ed111f9eb7c3cf9945645212f10b62939b45082559fbb9adcf2e1195de04ec176a283c37921815d4fce8d66ea5b45ef7e144ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc98f81c1e22496e641f800b0deffcddf3b949eddef3c61ed92dcd326a380069ec9780a10199ac0e957a1ce36129aaa75b8d23c18c93d22;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b8edefe3e5c1a196e1f6602f14e8ff133ebabf2dba86035410881dd4027ae9513ee8c1d928a63af4dafe8a6c30ff96c98929df02ac09a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde0be675766fbd74fd76962bf9239cc5cd5776df05232bdac75361c7df78d37dca3afc3e084a7268a63f916bbf9ae10a7f6ab585010501;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1173beb99e3948f415c36db834addf70488b01a121fcdfbd90d32231a77f46ec851219a84168133b8f8486abc4de74bfa7771b4086a6ea1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24248bf9941616d289780e9b52e0d0f0d26e47a87e743df213b9f1acc180f6abf37bfac497b938a575add292df6cf242ce22182118dc58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0c7894954f858a1314a911534044f0349ce6d2524ee5a1d3068d096b7e44908de21c0c7a18f03f229e34bc727e0692cdd7fd4b0861475;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9974224538a3cc9ac77d418f1f761ad568a54cb334f65cedac1c910734a540e508b1d9a4a3a357a9d1632cc198e4f441cc7bfe45093255;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h128bb1b8abdb304afb7257d5ddae9aba067d90890ed43c296b0d95f184926e235e6e2d36732b0af805b94bb04430450ea51d8076dff0256;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1e65366ec0d41569be72678168bd951c801c6083705d81c3d0295a12dc88a522cea0d2945f8b28772e7e310c3c653efe799c57f56b75c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6f3f601ac7f4fa428df39f0740e1794bcaaf1091c498a7b44713f9f0f2cb0756b6b9b827716d4fbfa511bbe80d91dd52f46cd8d6ff4bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d333e02bbec6ac87179f68928a05769e37dca170eedf0bb376c91bd614c3c368cdd8634c48a2311debc08be75ef7827b5640b424faa3f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10ea9f077ab0592e87a5bc87fe6a960a15e877270fbf0b9b1bd0e225a3e2899422634421bb967acd155f3ef28f3c25112a01c85806480f0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109487bcdffa982e5a7561bf857409f47a6371d0e61545887f189bd1cf30e168a18036374bd4868654b26ff38b78b7ccd6ab678bf0aa6b0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1042cc7cdaef2d6770f703135703e9352fcf7e37344c638e5b3c72d11a143225f31e82397f187e3ad7337e224a00569718986498a46bf0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113e5f2e685576d046824619af9307241f6364d2bd6c26bc3399348a5d94fdc312a2725d8a9314ebeff268b662b524c77b2f5ba77d9aa92;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d706d5e17905619830f1f5e1ac48c7d194564861ecf065b336ed7e541a620a9b57670d3c82eae94f4096481ae518bd3289d4115499dbb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1299b16251bcb0eb1b9d29fc98db9e240151993600313fbde8afa0bbb874659b9fb20d5d29b367272164e6360d439249cd160c44345b96e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e567e25ac3b40d12a44f9c6f362e4207cf6a72cccd2ff2b6f8c2f36dddd561887ecb217bc713877e9edc254043852099c1e3d793f1c86c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f16dca8085d2dddf6c9f69c27221ae705cefe759030d2e66d4e504106c0113bffc981627735cee8dfa2cac46c7cc957317d45da6a3b8c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ff239bfc9401c84a63afc3dfc7433e7ed49a9b12651e5ad7039b884899c7f457e9ac9eb667243d8a947478ac29ff1df980584f9eae3cc8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15fda057f8634a0ade6c81a33c4dd7fca51f774b6e598decb4bd260c6ef3981a69332be2bebf358f815ae307c0c2726087daf7720d523e1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c21c81b133c388307904421b7a8a66c2df56cf212396d95e008264bbbb1e912c7473c6452f818ecafafa732169c2686bfe4a24f720c014;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5eeb053a914e6cf9aa78097fa708430094aefa742233157ceb78356e4430ea966674d6ec672e4e5acb87a4575f80fabe48d4894021aeca;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18be06c827faf95e97017e21ff0bb3ff171bc0ce78ba8c0f8bf25f26794823fc79e120ccb80d40af8d38ed7e2e211737376858b8133dc1c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf6cea287e04c925f4e705a13cf4791b5c98ad12cf55449dc212311f42aa05de54b719f34089333476ca97c5f14d3d1c539a6f08141983;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20c9947ee921afb498631f6a06cbd76ae39d15c2080b1eef768d4bb0a21aec2bda9b9f4b1d97b6cc668d64684772f303745f0b15c59b26;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff1c4bad1c68d9ccf6c7d6217c2c3cbede897d3c54edc4a791edb084fea928ed3dc00161d4b9484ba68950bdc64754555037ed185b6915;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7c8be450e73989aaa2c5fa3b7b1fb83ff53cbc5622b7251ec6360def3bc68696c647ed21dd8c63ec117db76687ef3c5f252ccc8b04702;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190103e1ced87fb8a73934dbe78de4aacd18541eccb38ef982e2085cd957a8aabcfbaaf85c5190c04a49cb5577165598d1489b030758b73;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43bf6e224450f86fd9ffd5b9f3c519facaeff811a6e147f0286a42c6a800c80732d4abbec4b40a3a10d9d6cbc2184fc7e9fa565574af83;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b7ba0cf6869e840df6fe8f26cbfb186c051e4fd6c835c46d6eeff2b410b03d1caefb2456173c527b936a93c968f1537a94a5c0c607a4b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cc5789d68ac9d5bfaf81bc0929d3b4cfa53613ee1aafc90b1d7f90e32edb499ba6a58a2c9f2a04e3d7f330160f6e23a24bad07bf47433;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4eacd21fc4e5bab034997a66349c31495d15145396522b74c92999d7a40f71f1f494b9e0d3054caee197e91271bb7955ac3d88073f3498;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heabe0683012b7e0c69aa12e734fc20075537804181e46ac70ea5223ef51d8d532cdd7f213c5a3e1150ad476180beaf880975f17ac0ac58;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf600f88fb6fa833d65003da92ad203722bf3bf3e1397ba3934df387289d06edf51df23c211cc1aedbfcf16234a03994f788b49ea59d7d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f1d2fd5294ef991600b414ea04cdb28f023bcc882881748a3702ffbfd969f8c6cc6f6bcc0a1db262529d3004e301fcc55fd9e8f4654024;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cfcdf1922aa98134fe72f00c889e129d84ba6e68c8ca97960bb589aba7f9555a7a28e2dd1a9bd4b4324b99a484ac9aacaaa5c7edbf6ae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bef10c457e399c31fd9e21f39b0d3ce6803796d8df34973bcbff7a5ad08df02066f4b8339ae095c9c27bc7687e0a9bf4b5891ee23ff76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69a7cadf99235e8d9319dcabf150d9e7531437797a1768207d2ba9c544994a73ab69a34631bb7658eb6f02e173dcdd480cd42fd2de68d3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3450f70927c958490aaf28b742292053d26f75f4f3b046a26726bf9737b368f3094c1e8f4cf9f7fbb1ee4425c69e1a2846d96dd243668c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a4e3881958379999ca47d7954f15a5bba9a6b9eb6e4446e0be6d8a74ec30b874fadb82dafb8d0c455b1f0781b33aa6a03142aa57c81;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ebaf70ba688c132fb1fb520a431b17f00bbe6e75817a5cbe059ab8364add6bb6169593e6706389c9cfc677992bdfc83390219525029fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10873c52abba00b78753652991d178f8b17e11a2677b0d61cf32b78029b2eff7e673efff6907030c0b6fd804582d506f09a18430cd81ca6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a44e2d83b6c1634425233eae826402582f7bd378ef75a11bb681f831c821d885831da715cf3bf0a179c829da422c1dc5eb703b7c3b528d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf68dca0051f843a91ef8331aa9ecb4fcfbe8b9a4b6e5e70c01d8a606a4aea15aa6209e53ff30a8557b9d9d9ceccecfd6691776da876fd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf08ceb8c223bbf6d6251395c7fea5dc7a4cb041e7a7c7d9a936b8cb097b932635af26f6af10b7c0b6754d4aa02b2788682e996c95967d6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff696f8ef065b0d0bf0f055d7c0def391df976ccdfc03e162a320bad18231e28878403446a85e0c929d0d89eaecd22fa00d9eb942fb08e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h85b52cb47c49c9e565aed322433ede90d7c80bf6ff51ddad89bef941f61f78164f0ca334f8bc9e9c50c80740685861baf9c2916c063275;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h945818bd40cd2bedfba6a90338406db0519e0aec1969b9ec95ca3307737b3e962fe50479a65cdbd4d3f5ce59d47b6f4322fbab3573dad6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1536f4e555d81855375511f84fbfd5adb32e27bf823f6abd66d13984c219600f9285463fa6b3d55f94b959090938070844da63935b89391;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd40a20b66d972aeea8bf3ff439c59fec64dd5be37cd1ec2fe044643f72b47e5b76bdb87cd0300d802e02b0a3c1d816509de6c108956fe5;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he13402fb8455cefcc9533f9f333a952bea083ba77d24c26457b275aa863daae4f73464c244b3001580046e9faba5ecdd122d80f580e205;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129fb9c0b13a327e9af1f877bd9a87560c7e21ba7fcee6f14f53b52970f90067d2822299f5a803b003fa111724acaa28773e2da5634b06e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3e67f203f6dde9d510edfc64fde4aff8d210b168c79d278de4952befc9a0c78ba6eebc568560a4256a0aa6b13727b918d04ee334fe7f2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1358a720c8358c7d311a2d9447386f867a2d1c0624fd1de23c0242d91b5ba466c239e4d7f3c6028acf0c7004dd3ba44c359d094af8323d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1def05be5cd047f156c16370e8136969dc90256ddd314d616f255daebed98e646a53778ddb1d3fe1442e47421c6186af21230e805512590;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11951dc45915c50f550b294d9323d0ec55808e43b4133b0ad088c41fedb45d104ca366415d30e6676ed29cec1234e8aa13e04a112573d5f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65672e5a3fdaf24b7b7bc393bbc1d3fd4b94adeebe3930e0d247fb22181c2f9b59daaf4eb3b521086bb4056baf413553e15ba1dfa49ce7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a2961084269c4687bce59520d72ad7ed69e552864dd7915f11ba9fa3f0c620294dbe0b7c5150ec3b1ebb0df1d05be81b0b59df49066034;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he81c725bd620114bf0fe0e34159888a484c3f907676c5d25533187bdc14b0e3042c06cb4b72d556b9dbcdc11bd24159e38afb1785d2e77;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hacce4cca38d0a8b2fa9dac46a00ae236dad12aae48c4fd93587a2c80528ec951ef4d16c3ab0bb8537cbd6a0895e15e26f85fca77af4cc9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce73407a125a87aa28a7cf835157e7c3fa9f7ffdb13ae98bf87cad3a7f71ed79cd1d95848fbf7e87c99485ea6b2a4ee3aa096ea345a7de;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e3e030b065c010d708677a24ff32b11755e671ed82dbcaf0835ffe5631f574c48b84e2f15105f77b02dea30297cc101043329bf69dbf2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4699392db25d2212184564d75cbad13a39140e868a4c9bc8a63335ee22c62a6b1428e565ee7dd9eee15639f8682060945983a727a81a10;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec8bba39c93bb5c28ae65f1f7d401f5520796e3e09ad6caf8f2b2c5a472514782281d800392ec56b0ffe9c4fe5b7b17a97579561a1642b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h785a8ded7dbfbb229dfc776a4d3a39bac8486195e752bbb90a74b1efab0fd6a4f4dd37bf41ddc80bfa93d8cd18741c732e9099566f10db;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183c067a6f557ae96ef5384cd8d8a8050bc520b6ac0c427ae57653991e652805eb1a4e258a7810d07c3dda442915e594e3507c6755d040d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149f6ce2f96ec91f4f0193ae51183880171f36b6d0eb20268f678751776be5512bbacf6d6d553a5bacfa8ca2cae89d58156719c56471cfb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4390fc6fb06279a8985e3c81e9903d5b184b635075d36334e355fedfe59a11aafe6f6148e53862bf7e7fa50ab9bd200d5a891d2857e2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1187d2a3649a0c95f22597ae1805fdb493957c311c51fd3c83168b01133353b1a771407e90b50b22a1af36bdbf4ea146ba1ebde45c0b41;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e3a1e352579b858b98de0b8da6a36126a999f8953f05061fec497080aae37c7339eae13ec65b488eefcb85cd8ac6c3f46720a9a461815;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h144e55f7f615201c77c76d2ed1154e70406247bfde8ba6a7fd4dad15fbee831ecc15105ebae58d8a4772da09956996bfaef6666154b01d7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha00a56b6687e37cdd963ea4619880f9eaf5839e9c8282c422fad7c9722ae4d6d932fbbb2a7a3037b0cfada5bc5f4123fe31da43a3f863e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3051431199b2cce6da45cd8595d0be833f5ef93b3aae84da453b98511fc8bf8b39fde11e45c2e84d687d91bd641c462892f1d11648056;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha578c0faeaf81500abf7cfeda6863f8728d4c6fd35f9cbdfdf945409fa5074bc297af37b26424ba554a0492f8382e5d38a5e38b51c0f5b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173ba8c40497f8b307a413f5f24420295b5d290261443e54bce9f6765e17ba4c084be57e4b7158b9fbb50e81317fdab6ee30ad097a36945;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cad1786361a9910fd90791e5814913d3abdbe2bf04c1a16ffec448efe57532533d7013716ee47f734bf54dcc13c868677d525ba8c5ce20;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1657fd341291434d4261de7589aa88c4ace2b56f3cc3f981bb24ea78a189f91bcfade42982c54ad453604b9447a3e96e148a7e52ae29b01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b137f22fa56a4e2649b57fe361997c5e0d8f0c606dadf85854b50b474833e2d7532c0484e04c8b6d0ef92b9e26e538a588adb80f027fa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1840eb4246914e51823f7b8fd1dc97d9979c3dab8dce196978f11bd753d3c726bb360cfb87c01e62e914d964a503be2014963fa96bfce1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14305f9dc549d2698b8cd87eddde81eb6d7eff0b97df5a60be109175c65bd8127dceb8f6341b58a1d6d2ec53b1198c3269f0ab645c6e4e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133727148978c89e7ad8064d1755092d791c04aaa12ddecc6d8be279b987273a25e15035d9db0de07cb0afa86ce56c8c13931babdce5e95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d15fb87dae11a117a5886e7643e2ddb56a7eda522d5e6e04af950b7b5ce06f538d561769b4ffee3459dc99bacd8e4bcc42572393b9d8cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30768a6135f056b18027f929fef9408a37b1383b4cc3cf218ea3a69bada36302459c8f26f5dfb794a83793f7fb5c0a362c42e7572660c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dcdd012bb88c83de0dabe56ad75eb10a9f5ef9998486e89a7c9a97adac2320c2e2a842b16d405f0e1c36baf85d8f10e676f3164dc817a7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h933bbc50adef31944edddeaf36f9e7df9fb0008ade0a117c51c94ff9c5ca2336eb7ddebbec7f7c21123333ced7b9dc540c399738fc2df7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd8cd845bbc64e2394b15d8c3ad79dea7039b26758564373a86d8543c606bb08179a6c6e1fa0851d22a6c61abf3321ad80c44c22e3814c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb46c55c2856d8682e83968e2c7c71e51158df9add7e01ea4427169457033884f087d66e4f36463685f233be14d19948699cc996c43a75;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf8a9d882df6953c60043cdf106f5f85031686a6b9674ba2eca955576a4a9ddaefff5b27c3491ea28fddbad2ae27ae18d10f9f9a8218d25;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171aecf438615096649c694113bcab828fadf7cea1c7e4c29cbc7f37abde709c6f43c9ddc429c3b389fd4d385e86786002a549c8f7949ab;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2c2ba7183d27b96099565bcf35da4af7bf7607df097d0cd80e88d6a644cc8a641ed4d4ba51bf564a24ce8801cff4de6fc8219972da189;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h473090fc11bf020fe96019610fdd8131e7a6079abf7ac305e11fd90337bc25ec6333f68b1452281cd234c922405326feda30c643a52943;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1692b0a1dbea7511cb175f3e29c43e34f100211f7d1b5aafa438324d99a8408bb35ffb25a4d30924d9479dd1e00fd6706bb8e176285b491;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15616e5d9eaa5c0b1ccf7df35c512521e5d43316fa84b7363f5f6eadcccb65e02a7af2b6f09c1d3f33c7e766132c330559840697d6c1d61;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5596f6f9bf948d62fdb6f73ff9b2785bdebb7eebc9a3e567e661f3e52ace62a182eff603da7d5e984e40d7b9ad817a632be3e9683ad95e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187d71fb4ab9008e2a13096d7af49df0001c65ec4d72cc9e6aeed71dbf1f42118e4338eb2c0a296145ff8bd8d9a454ceaf4ab5a22bdd891;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d339229edb3a2ab9837ad356bf936cb6b6ca69b1dae05bc0055cce06be78491ed68eae2e4214c0bd94803117dec78cc15ac3575791f72;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heecdde7fde9892d81807dfacb957a0d290bcfd79fe02d4030c7da0644ad6f5779c98a37ae83cf8c9037e9de7ca3b37306f5bd4deb0450e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h127cf2a8c96d6346907a1a176e575470d48911c12873e48b8586c68e952d76365756b64873b3658f45f41c3647a3f97406e764c01afa654;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d951e42ddff4b3111cc600ba0edd3d18e63a8d91928b34ed1c1f8f834cdd805d29c1f659afeb3d5fe53c90dd56031fe83c87c8c51b8e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h89e4d9335827382232dfafa701983aa57cb743a6d6c8f6f0051ac75fec0ccc45db4f89c64834ceec6eb2037cabbad85adfd93ff8dc6ef6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47e3f981d37d0c564f2a5561236a018a809ce603d0e0851c018478445464e471f60de70b6e9d4ea8af47f6ff7f300ea752d3445b8410a6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f66f1a7bfcf6b3752b27c28f2dc308538cee292ce6318a5bb3dbbc2b95940cb9acbbe0bea29980626e25dc726b6a5392890861874ca00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb11fc3a3808bf4882fae98ac42c3a2025872df0e0a81122dffd7648bfa1590756e1edabdfa3c8074fc4f9b83475cb8b8420c16da5f310c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc02aa1724a3bc23544e4b1316ae82f0b0b9bfaa693c71507a6342fa856f971badf5df0e17cc00ffb0c696db4c856dd8d3738ad103de176;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e40829ee556dadd5728dd576988fdb57df694d3eeb5fc2fc109706c198377f44dfbb17ecf693da083959ee2d6f504af6c4b7b5c8bb5887;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e286da8f7beee33b47948c600159f7cc5e397d2dd8b1ca1c0d412985600b5f6e528e646197affcf307d86581a36486718fe8835c4de69;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88a904e9fbf043d5c869492b57e9d686127c4803cf22233120f239b29f86acd90596aff8a0c64291e95476867e71a0639a630c322e85ac;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3842f3ae19f02eccb2d59a2b916e4329df6d0030de6ebdf6c8506e52a704e2e91e08c269cfa4d1b1fab4f07fe61c8f2d88954e50bd969;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfc7c2c341b47956b91cdaffdf91f2858521ad8c22fc04e91fe6c8e6f7a23082abe9a799e2348d99aed754fa4a23670e3a87e6bf129e85c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3e137c37029605d8a56581afb41ecf750a5fddc14e72da23c90da70697f059322fb31129e167d92965db71290a2dcf38ba2bbdc6c7191;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e5e86125e291903c696cbafa0d1cf6484a26cd45fc7f13981e261d64908e3350c8b2a8945b6e9e4c3962835b302bc0016f7835b66d549;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcda2b1809eded87a17687aaee7bf0fe6dd7d5c280cce90e0ec11d03ded6da49501bb9c032bc41b23554b017b2fa4fe857e8e6c9f8eeba;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c8f1ea8d7ab6c2e5d2a667f35609c30c4d72cc82c7b78356eb98316acbd7b9124f01b1f60b23b97671a5b1dfd9ec52bd11d971c701a9b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c54ee8ef9d311e38739222a4fe1ee51c308584d55db1b213f109dd07e3fe0a341ad1b42ec6f4e24da0e5bf6009a16bc4eb3d7bf941735;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1514e2f0e7088ecf95ea43d64aef18aea5a1712c8d6904adc0f16f7489b1ae7fb3f7b36effb7a522006795c5b7da2e3b9cee271cd11c431;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ff0821b417067fe77b26c2d1caac0a5b6329a9215ddc6d759fca4369a6692c022b44d03d20f46138cd1669e6eb2bc15559cf62051333bc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175c04cb9184660ac4d688ef8d61ded844060cb0953bebb51ce9b49f6c3ba7d91cc37f43bcb66abc9443c8a3016d0a4060635c652a02b31;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f767fd3b9b5bc9a27ec959a4685783a1a3852458035c240ea8775b5a8f333c3c58620dc777566c63343f7af8148d9abc5f2d42ead1ed8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h417c67c54c7ab4767f6b7c1a62d7e668efd96c13ff8fae907c97b2a6bc2ca718287bdbe83d71eece0e5970dd0857d07ebf5aad89c663e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h84419c2a8af14ed32b1c6b5eafb35240050347570133439d956fb027d5c5d6ab26ba1048390d17f9b154320329e4b9b10fe49a91229463;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10573655c346118b041712b6ee600a94e8787a472403a0b5d7830be284f234d465f7ffa893826542bba91194a335fd0366becda2afaaafb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ddcdd92e49c61472988b7ca184d51cb91fc681ac545a39f464deb8da27055657f6c4fa6ab5049c187fbe76bc3cf0edeebae9e9e9000e1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb50490308ef79bd06df9a1c820dcbc216802c263f94e09583cf50e3d291e39279bd01c95405a94d1915a2a75010e57ec0ee00e90b857b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14024642807f36731d62349d397f138569331cfc489269846a0ed382793f4ffbaf16b9f7177ad1abfb6823cefd0777da19785e6e7ee6698;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hccbdf1b60427dbbdf8268e7e03d1e53b5873eedaa3f63c52c0d3eb21e1b58d3fc16869771bba59e491c7f321429b94d0b90b20125f51a1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104ed0900805af15bbdaea3994347be5bf7a0569ca2a83bf599aff2956d6e99ca88092479ade2ee1a41b5ff61de9664895013bb16d80579;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f14846f38a97adeff42e6f80cfb8253bb3b429a002597817307e7059aa5de9430597d0620648ebb92ac91e2888b4833f2ecebcc964953a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146a6f7f042750546f87a963646ff8166e12c676916302a9f484b956348175e23c9470020f5833ff6052f897303502460896d48616c7f7c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce4c0dcd6e81f98896c13766f0c146fc5b02fbb4519a41a77b9d584193c31c92a08b4cc8d16359b702e7144db36a30843f2e2576bfeae;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e0b5dba46ac683c3be436647681baf59bff37365313c190637e8b8eae0d154fd50732bb2c74ea9089044e88bf2d9e6a2b74f9e044719c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130317c659671bef3c1128a1eb5e41119a48641e47119f6e08cf72f0d433ffb488b8cb8b1b0a369eadf1f72218d48be0c96b7e543fbb897;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc378fb4b45c74b263c0af3669b0a07a5a11a78082d46921dfa4f6ad4d87083df6e0042fd04b3bafdde30ad92508af1ca4802b7e693c950;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130ca9a026750c7718e7bd47e932070d90932bc3df3cf96c5fbce3e1f632b8904b2fbff3d67709a06fe5192692288f81282e7d86bb12b24;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h818a9e179a111e66bc8e8b5fffffcf7ccda75856505d8f78394bac5d7fe079d5983f50e23795e7d652b097543ef6313eb235690c94d203;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1795fcc3af185aabc7a0b2697953232bf5aac535030b3bdf117f75634b0e0e73948f538c1b003c610eb1e1da92308138a6449252a1ec955;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1508dfcfa548981fc1c8a7b854568089d9a3ff21f4a6473571a83ddae8d5a8edfd980bbd4401c61c7df2791d518ad1eed0a6254197ef9ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha25c171fc3748dde25ddb4ab9a7e944fb633a9ae822381c721ae73f704cb195262671a7c730797bc1786fecd9659835a6aa93f4d2308d1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f7ced9f7c5c0a2d5981387fa57b0f3c5361948c13f7494d411bdc9f8d90b191ffe1ff622343de72d01b16d183807e0cf829e6ae340304;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f84ee9e0993dccf38d5d08d994e24cffe995b2c323147589f057884a36a9b854aafff96a3015e02030b102dfa384806d77609a31189f9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87b6434dc49bd14736cdaa22e71a678681f29b32a9496f15417ee37cb1a85292a465b61e6b0784892c156f2eb2fb45dbaa627e3ad597e8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e3da4a9896a22d54bf29e2958184dff56f12c2e4c931fd87f9fae66303b67009a58db49b34aed6cca7f3c5c5d905d6723f09c4b269118;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e20849b645f238d23278f1e50f87b69ddfd10c52c6cabefa4ea8a5715ae365911663b881c56683471ad4effbb65cafe1b52838d707fde9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dcfa8b97efbccb9f41b856f506af33fb9f22ea65be5156e4ac081cd9d69ee662de841967a209a7a4ad18b7d51409f04d110bd3861061df;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc596e622b3138763ab71d9b077ecfd50324d502f7ea59e56d80d42045d6832843d8f7998c66ff55c13f885913e8191b6c7846a29bb968;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3c1540e63c9df95ff60bbc13af2128d0d70e079189a21a47bd54d660e77c41d7ee2a46c05277a3b9d9c136f83fffde2391cdcde59a08e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c6d5f64f8ffe42ddcf4d26432dbe17eb1aa4bb499fcac417fa7616775f0df6c2c42180bc77aae7566d5d95988c2dfa4c650b3a1b24eef;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcee4066308cdd495fa389061f3fd8f3e7ef823a08ccbbce1d07c4106cbc348b765d0d3d9d027d2ae9e34808f447510f9faf6eefa474f43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14128572ba3c3816d45f4ba35cd2f33bc7412c5cb2b2f63cacee19f90af4ae707c40b50562b3468d22bc92838bce59b122fd9f4a3c691ad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166bc820d494a13bb865570d673107489356857a5b7f59ff854fe5f97d8f66423d81eaed647206375d5f7554701209423c2d0d4d9eebe84;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1874530138958e564d83b5cff780012698a5a3a4d34f4b186e1fddd6f7d0faba34586d3953737596989df8983190ea20ca150769ab37e3c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b35284cb7c526927f7d1b8dc27ca080095a92086c09e48b38649885e2fab4eb583d41a76420cb8bccf2d8102430e13449a6b9e69ed00;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157a05eac04fd211a398abf698cd2679bd8561a11c11d0d8ad5ff5163e542c8104035083a221e95711bb9b7496e72b6a6defb04b091e54e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba620335a5a4a452c9178e5e27cdd4e4e5e769e380a83754b5adb6fdd804360164a76472d2dae2bfd90d710cf8f11b263d9e1a2fb3384c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66d07a0ce70271a7d9d6fa50b99b962c280dbc4e6e7c1627d0786136fb80fd635a56a9828653262ec7be807199ba41e6f93e97defde8ed;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he69c6224727ef48824ed60d32967cceb833768ce5ba9a3eabcab8d3b1df37b1211f72cbf84df3b80fb5af3d6d21bbda4dc058a2b6ec0bb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aee1a64ce50f489967e3040d8951bc9e38505a1c21452b56083d19608223082074d6a9e3c69cb488b7166cbb6000a31b9f9cd714e0af43;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2f648f2b9fc71f8e46d3f55d2731af354547c18e52133991c2386ed8d8390ca5cd95a27495f736f3e8e6c705d7c8fa05fc58414ad9949;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17485959c0ff74e4ab45f4971d072a75ec960ff4b7ff3cf84190c66d61662c2b6dc9ae338081b7fde383e5ba96ddccd786630f7c6557864;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h671e14d03fcf1159a6e9c6e2ae950e7da5578950ab5ca78b17b1c4ec713731f731be033646c9ab42d8496dbcd988f81fb6e13c93a4f560;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he97a8f86decb2ce0e8a594bd19c41c6b20b11c18ae00f9a945ffac22a4f49278598994ed55aa0a016c28b9ab1ecdf8db032aee07b8b7cd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10be3ea7573e6bf86598d4e71cfebfe144ecb1c25f41632eba6fe7588009a66467e1b6d8bda12eb4f1c4c1b0b01aa745036208d97869078;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h68a976b66f19f8bbd7fd8d86df5c9c9c595f2307187becab70499b6859fdad10d8c04a50dd134ff699f0209d6b7d45ce856c608a313670;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd92ff108c8e40c70db25af780c89913987f0453af31b89ff4104579129d90b36d88a43a9c0f971fa110fa1d7732d25a3f727e714a3fcec;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19788941b213ca51b1967bf498660a2f4dd563eeb4d3f54195b510984995e817563692f61cec8bd50feaec2d6d6fb941e3d89baefa058e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d57103a87a141f8b869e1f1a91d17f772655c274183f41a755f7b8fc2a05fde786372ee02a9224a692189b92437f9440285d396aaac343;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d370b6e8d756ebdb8a397f2d8c0e1706dbd4bb162ae405b1f504c5d9e5a5b511f2ca606b8d0ba3e2165bafd5aecefd38505b4005a6a98;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3de74261688fee31cebd7b388fae42cad9ed29821b7e8271ab1c2c7b69dba9e1c3e7d26b8ecab8e52b34dc0763545a58d3fe0abf1076c3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd51ca78176935c027b84c91c0dc33a78ef28ad859c6e4f76b0e3daa8e3c1a2cb448a9d22f29a43f96a7fd1f43702742139c628ab6e078;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8734ba82cf00a26f0925c84b9e7a90c7cbe694d7b42f3b96f116849edad090b8184a423ea31514d1e4e8247b8f87523a28782cc8dd657d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbfdc16d79ef03efd322c02800ad8ee1ade99c3e3300c392e111fd73e8baff1b98cc80ca366eaf889409e40e51a42651348b0098c1d8a2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdfab5f4508d1b8b7f89b29505b6a5b5d74ba4ed2cb3dcd783ee997db2891ee63529394b451f144bd2ff394acdc7371819ca20c8c53bcf7;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2bb113b63b5487940e6eda4ae874d8c70d3e7add48be5d0a9569a6f785997b2261408591681d18bae7646bca0f7555936636d84f30be8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4577978d84da25c57fa2324379c091a0fc46a4071f575cd91e064b3e9e793d917bde56860be6d37c68df188b21632a116db17726c586a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59633c12c69977335b35014d3662503d21c76751a6e944b61a42bd2b9c5b11faf8f66125e0aaf952e6809c98cbfda85f2e86ff0da97a16;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ae6bd5c30d3b0ab7dbeaea91900ced3714188bfd7419c4dfe5982c6e3e946b5272d4b9d765cbc4e11f251c758e6488e540be49579beff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1945b86afaff7394733ea04bd9f85b14f2aa0d085621ea5fbdbbcb714087215de3fd265115d5a6318f6f0f8695969a83af1f326442fd79;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e6b079049072f9d32a84eec6a047dfa898dbb343d1d24db2b026884b62a682f4a898a27af3847d9110b6fa9e9c50f6bc58b09c268d332;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e6cc2910fb64ec657c0dda784f3331d3e561f1383cb14b6be81762133e9273d4cc4bea3b1cf6419b8d37d331e8aedfa01b0a61aadd572;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e659ddcb2f9fc161970477ef92e2298f4b68ed5bf350a658227ed2f9d8ba91abd00c3048897e3b8032127f4a1c507d876340e88207f325;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181e92185878899ece423e1a425dff8be84575cc134c349db4e81cd426454ec9a0eafa572c3919525af5e5319b4c2429691268eb14e7b7f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfadaba06d80665f2a7c3c329e9c6902ee2821b35b7c017f3feca35da27f0b329d0657ad501aed8e9ce9cb21ed575c8e878cdf80bd96014;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10c28cce15d5b39db71769e0c419593be69b57a69258048d6d330ade6f910e631b4bab164b96b44faea8d1d59ed4f18aca908f184fbb081;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f38639c384099667bf33f7fc858f93994a4045ff15aaa275e2a9161c43cc3ca6f211ae0d31874e34d066c8baff6ed770e5f345004d1c1e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7cbfe86a9c6c5c1c00a62e0e7397a63e32a39a04f0c15eb67b6a2c628101ada672d642f632598c85649d6b345a2f63b2ea79a9ca8569e9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168c90a12c89e116543df641d308f0e0024715e9f712f3c8a6b48f01aa96a76bff10b2737c9e321489fc2e26e268b99f308ff23a8c3e551;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he24451450d7a58fa6cd595a0519f124bc211337024452644804ab478f6d47bf10b4577c6a303008386c61284a15e36d1dc2c189af7401c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce0331b76ac86dfc357b0732338ac09a1a84120e18c56af3869096ebb17ca671c8ac6a24cf6666cd1ad92c91259655c7339a6f72182db6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117fedf046cbb1aa464d0392d468faff573e7c6b526401be68ec1c2ee0fde6936a80c4641e89b178e10c5576b44b0f5b77316b9853ab7fc;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf2822005defb85b702f15d6d2ed45b98aa2c59cc1b8a164d64e8050ba9ffbce9905be79855aaf32042e3674b1eacae01efe29480f8d62e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5baa7d0a6c7b5b1d15e44db1807eddb88cebcdc20f0e9c7f7c1d59d4cdd5faa564c272e3d293e272528fd2f5d6f2fca943ed4a522bee1;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15c9c98ef5b49717671b49b8c84f126c4acb005566b2e66cd78a3b3a206532297ba4303ab7c98ab1b293ce6c2ac786e595e96cba7696316;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73b685b6ece73113ada64747e6697bf881a518a40022a57dfa58f5435a3e6ed5b00371c7b88025536ce7a57471b79c42e58e255749665c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5eb4600030f442a1da311435a29e8622d414ed0bfa91efc5abb32b72c2bc11b9dd87a658cc3de5e3bbd44d36a9f451cf3186f668bbabd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha0a09b6a2922a66ca05a05b998b95ae2960738688daf44e40dd58720c7d376a734f00dcf33ecdaf446ffce546184885e06b309007a6945;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182cf55d3df6d83e22679eeab3b5dbf0222e5b53bb2a114abdd2f5c1a2169e3b64e261ad3ccebafc4a4930af24bc7fc88a04520a5511a03;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h616da0b12419a65b595066da9e42fcf3eda51c42cc602c3869fea6f3c3db3958a4c364b2117f319e2b01cb1cdebce30f04619dfac55aa;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1372c7689fa0044111330a43525f0a9df4374753c08dec81dc601e7160bf3d0890e91cca7f7a5d95e9a9eceb1011ac402051138094d7f8b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h174d933586b14d3999e83a4249773e54d42a7bbc235134eac88fb0ab523a33520952942dc4e2f076f334a901543bea60c328f456cd53dd2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h489180c3fd408ba39aaeb47638a9312751666bd45a4cadc30f9f22307898c7a76c7ffbce63fba77b50a26185cb0587e6f87fcbadbc6438;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc9fb03ceb55ce26913681678777b71c0c43464e0969b2c5c1db8ea5fbec7bda00af7ef4489d7bb46e65a58d7243cc8ad14204122ff470;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbfc56f2b516bb33c48c609d54f8d59f56b81c84baf05f47f17f5266f3e601d2d44286442421e659f3f9e2f582deff50cc4a8d78f23d8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114a57616696541c853d2becb6e252cef83c19233462dddde21662b0df000edaa053c7122b5768f0f722ed7d3257ddc5a860a82254900ff;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161f6d347b1fef65a502ee15c9a7619398aa42299bba45a4f292d7ebdc83e096afec669ec4f882f59f5b9836a820d777f88d3835889f1b2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d4776487f0f66d558d7d5c0f0e8dfe73309c3cac493d6b3a4236a3ab19464228cd74ddbd73624c78316a3192314055b28839070f66cad;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f2993d08ce26d381c7905a8778b560297dbe0189628a9dc851e341a170c2bdcf6f550faedf2977025476e71ed8502addc0b5240e5351d;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126ccd455945318641ba828b3909188eac960c8198501d55a5e4c0f77a3745c79af39bcfeb9d6286278ed133eac1a030ccb8c9b07698b38;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e833517fe9004428b4592c485660c6d24dc73e09dd69a9bab44cd3ff427765e98aa3c8f4ac02fd93ecf051bbacf45d263489ec29ba2f42;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h295877eb8d44c163aea1cb969e9e95ea1f405d547cc4b41abea574b4d99380e1cccc532b58d421aa992c9cd1a76922b0c911876417b7f9;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b06d0139984f608804e493d66bc6d6379691fff8073ab273d3ab4a166adc72a1c67398632ac94a853e5a9777232fa334567ad24170c76;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1eb3083c35585d977d7120e9df259fd5bb2772b2b1098e8b05ce890a0192ae9663ed93f0a3a02ffc47ba1638f717a50318d626e6709be;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha44ed21dac5aebd5d990f6947f05b7f1210364cb1144e6e3c63aedd91b471a7d6d19161742a9d0a6375765a5bc0db637783b2259fde3d2;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e93a6a07e3aad22df0e86e08cc42406d515e6f9220244f79bb3686458703276df6d41bdcbed01d5c71355235f303b2e287f3004717b557;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bd4f395de9089cf8d6c680cf8aa5bde79da258f9a6d18b9fcde4f7cd6cbf37d970b5956d1689ec1e386f7a6934daf1a80c4a3dc4849e3;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2548df1c58a2c9393740909b6dbf6f4bc88c5a64b1a3947402143407fe94ba407dc4c4048ccd76e12b268eb9a92b0a75c9d3d9d224541;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf40eca3a95dc93c952ded4d90f5a2c90de7cdd8e8ef860f9d8f87abec0893864fa4558a29ab2ffd4fcf89b285731d17a167df04d077bfd;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4937716a34d73c45112ae0c76afd514edcad4e408ba1553e7c732523dccc21027191dcb0793eb5dfebf1d8c7f660596494c1654b1916f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc31facd1b4a9c84838ef3717cd84ff18387279a862c4b6aadf29b9531d36d772dac89a265fae3c5460e54065ee451b3f7dde4467d515f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc73ccbc1d6f8d0a9fa0a827f05d59d4b768be81026730dd9f7efd63cbefaa668f83c3c82ec4d6f09a9d1557eb3bda20f9f613b55f36cf8;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8e0da86007a4a3985262dac046596b7dfc693070d1ceed7f836dd2ec6ca0ddff6e119f0b2b63528142951b65927066a8444285266ea8a;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f55f9312729d2bee56483d831b6a8c6e24ef67de8d3dcf86c52c3b3d12e365cc9551a12dd7d98bc57a6da0d42a817a21afb9b904cf182;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11141e896928797503026102fe17c6d556bd80123992a3d10cca4ade693cbfb12d7e9d0190f447b42a905413009bdfb7c211da90dee7b23;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1636a4e58a8e08893b0f1fd4142c8ebe87b37d30a20779c300aba5da394d78738b8f2fe4e9acd5185c357dd51a93f0c1a04b058ee08eb5c;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc38e4e31edec53b8b4e60fd6c897af97f9d0251b7ef16890945f3586eadd6c35c761bfa421afb6ea7d91db34d3a013f39b582f7a1df86f;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e7720e6c0a886791f7d9d3778d249788c5fd1ab1557ff6da070219fd067ccd57d8419517992ccdd4119209391c917018348a4093e38e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2e1f8d036179143dfc32d604e71d6e4abe61b2c738cdc4a41561e8f9b47e7feddb6a4fa1d17c28a0c6ae1e459b152888f5f394cd20c63;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc91f4b07768888b49a52d3960c85ac315b0c203667fdac4635560287a6229d03a009cb0f7961e50e59cc0cb1094ed668901f930098cc51;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h119a39ae65d01655f56c2d09254073280e7c2efaa9fdcd88fb812539b96d10703327e65cc4cf6d70e5633f1b49035daddb5e868f2e5f4e4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h468cd005e48461a6c2c4fc498edc5c33e7881ac2e2c2987001418d0b4695e2350c343920195b3ec82e564d93a6b8b4d507bf23daccaacb;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb24b3a2300fb4c5ad12db3835b6a64c8e7454d3364fb7b3315b38804ea4fdee74b76f2c797ccbed669a798230fd4cb5e8be2d977c7be0;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f64d72054f6b50c1ffbbb03aed1b52bb5357c98200ce7f7562b44e8a60b4e6a1d8e858ddd83875b2289b6f457a4250aa73a320ea967d7b;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1f08e348d397435da5c5689e55a17f66ea86e39442e3e25ee066a200d6ed2342f8d2ff43c5b194880082653512c9cb6d0e16596901c01;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ceb8cb2b72f26f247e49ff985e6ffe63d93d853615ec444e915a1480110761154e3862be963624f1ec9677b43483cf51889905d6d1573;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3497d0e667721d057f22b27563a36b2bb8277e433b1af74c16755d678605a33c71b4ef8b355c0acf6dd74edea7ad8b75a5f44db0b4b836;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb1229b7cbfbb3b40385acc43b81019f843d88e6c1592936e86e46cc6e8f552e13aed4613350a11156d155b7eabb83cb94b31326eca739;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab226e3b08e3fe3b5cd76ed436adb0b36d5e451f8a9af90d846c0026049f1f6fd302b56882a80437f75152039f9c51b0718669daaecf95;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3513c838abef287dd0a7ad0ba71389a70e2e6c1393f52ef8d534f0881785030aadc42f087bcdc4ca5595960a18a7f725781231e2392621;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1642a987891e397cc9243c690f3aae1fcce7604bc52e8e032e01817208fa47acc12cc85aa83cf570bbad260af548484854f136cebb84540;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdff9d63ca16ae0e9a53a03de1f09f4ef808b8e648df302335eea2b2f422d0d5c578031375679742e685d2dd960510880da010b2ec3e79e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a10e88ae772511f9debb3c91164ec1037d5cf9808ce949a966e1b46e9402453d94b447292cba6593144006530259d8eb7f18d2b0035854;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b0de1db6f86fc5d5babedf268f13ba7831e9b8a6c00fd6c4da9f865b0f9784f45a44429c700c417d2cdddf1f07094e29671b8e8009ae4;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b26d75bec25f3928bfb35dcfc210d7a09cf6927d25d6a0c365c5cb29048ba69c6f3f1653be8d120dbb2560f59907b5c63d24d986e1b57;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17512bdb54e88e222ea22772eb1c67f57600af9092e25747723f36f7d38f42eda1791c1527a2edc73c243b902a539ff65c1e38c09644820;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0eae370a703f240e5aa2a49e56502ff4988063e981933ec18d7ba8bab41cb0bfd743c63bd14522ac2531c12175fafb4d65b4414880b9e;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f975d62050cdf4013318dcd748a2cf78d2ac6e2ba1bc667083ea98c0a1f1bb313a5ebc661b02eec780170e6dee4711170a945d7f5d9f6;
        #1
        {src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19055a8bb5814316c785a5007923251fa1ca16633db436e5597c183549e02e95a80ddbca8cafbabc8066b412b3edb1d1a8b3bb958bd87a8;
        #1
        $finish();
    end
endmodule
