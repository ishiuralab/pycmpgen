module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17);
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    compressor_CLA64_12 compressor_CLA64_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17));
    initial begin
        src0 <= 64'h0;
        src1 <= 64'h0;
        src2 <= 64'h0;
        src3 <= 64'h0;
        src4 <= 64'h0;
        src5 <= 64'h0;
        src6 <= 64'h0;
        src7 <= 64'h0;
        src8 <= 64'h0;
        src9 <= 64'h0;
        src10 <= 64'h0;
        src11 <= 64'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA64_12(
    input [63:0]src0,
    input [63:0]src1,
    input [63:0]src2,
    input [63:0]src3,
    input [63:0]src4,
    input [63:0]src5,
    input [63:0]src6,
    input [63:0]src7,
    input [63:0]src8,
    input [63:0]src9,
    input [63:0]src10,
    input [63:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [63:0] src0,
      input wire [63:0] src1,
      input wire [63:0] src2,
      input wire [63:0] src3,
      input wire [63:0] src4,
      input wire [63:0] src5,
      input wire [63:0] src6,
      input wire [63:0] src7,
      input wire [63:0] src8,
      input wire [63:0] src9,
      input wire [63:0] src10,
      input wire [63:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17);

   wire [63:0] stage0_0;
   wire [63:0] stage0_1;
   wire [63:0] stage0_2;
   wire [63:0] stage0_3;
   wire [63:0] stage0_4;
   wire [63:0] stage0_5;
   wire [63:0] stage0_6;
   wire [63:0] stage0_7;
   wire [63:0] stage0_8;
   wire [63:0] stage0_9;
   wire [63:0] stage0_10;
   wire [63:0] stage0_11;
   wire [11:0] stage1_0;
   wire [19:0] stage1_1;
   wire [23:0] stage1_2;
   wire [24:0] stage1_3;
   wire [27:0] stage1_4;
   wire [30:0] stage1_5;
   wire [23:0] stage1_6;
   wire [21:0] stage1_7;
   wire [28:0] stage1_8;
   wire [30:0] stage1_9;
   wire [25:0] stage1_10;
   wire [21:0] stage1_11;
   wire [18:0] stage1_12;
   wire [11:0] stage1_13;
   wire [3:0] stage2_0;
   wire [4:0] stage2_1;
   wire [7:0] stage2_2;
   wire [9:0] stage2_3;
   wire [11:0] stage2_4;
   wire [11:0] stage2_5;
   wire [12:0] stage2_6;
   wire [9:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [10:0] stage2_11;
   wire [9:0] stage2_12;
   wire [5:0] stage2_13;
   wire [5:0] stage2_14;
   wire [1:0] stage2_15;
   wire [3:0] stage3_0;
   wire [4:0] stage3_1;
   wire [7:0] stage3_2;
   wire [1:0] stage3_3;
   wire [3:0] stage3_4;
   wire [3:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[3]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[4]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[5]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_1[6]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[7]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[0],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[8]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[1],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_1[9]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[2],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[10]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[3],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc615_5 gpc9 (
      {stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[11]},
      {stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34]},
      {stage1_4[4],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc615_5 gpc10 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[12]},
      {stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40]},
      {stage1_4[5],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[6],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[7],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[8],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[9],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[10],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[11],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[41]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[12],stage1_3[17],stage1_2[17],stage1_1[17]}
   );
   gpc615_5 gpc18 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58]},
      {stage0_2[42]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[13],stage1_3[18],stage1_2[18],stage1_1[18]}
   );
   gpc615_5 gpc19 (
      {stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63]},
      {stage0_2[43]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[8],stage1_4[14],stage1_3[19],stage1_2[19],stage1_1[19]}
   );
   gpc615_5 gpc20 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage0_3[54]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[9],stage1_4[15],stage1_3[20],stage1_2[20]}
   );
   gpc615_5 gpc21 (
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage0_3[55]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[10],stage1_4[16],stage1_3[21],stage1_2[21]}
   );
   gpc615_5 gpc22 (
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58]},
      {stage0_3[56]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[11],stage1_4[17],stage1_3[22],stage1_2[22]}
   );
   gpc615_5 gpc23 (
      {stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage0_3[57]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[12],stage1_4[18],stage1_3[23],stage1_2[23]}
   );
   gpc606_5 gpc24 (
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[13],stage1_4[19],stage1_3[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28]},
      {stage0_5[6]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[5],stage1_5[14],stage1_4[20]}
   );
   gpc615_5 gpc26 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33]},
      {stage0_5[7]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[6],stage1_5[15],stage1_4[21]}
   );
   gpc615_5 gpc27 (
      {stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_5[8]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[7],stage1_5[16],stage1_4[22]}
   );
   gpc615_5 gpc28 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[9]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[8],stage1_5[17],stage1_4[23]}
   );
   gpc615_5 gpc29 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_5[10]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[9],stage1_5[18],stage1_4[24]}
   );
   gpc615_5 gpc30 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[11]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[10],stage1_5[19],stage1_4[25]}
   );
   gpc615_5 gpc31 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_5[12]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[11],stage1_5[20],stage1_4[26]}
   );
   gpc615_5 gpc32 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63]},
      {stage0_5[13]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[12],stage1_5[21],stage1_4[27]}
   );
   gpc606_5 gpc33 (
      {stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc34 (
      {stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[14],stage1_5[23]}
   );
   gpc606_5 gpc35 (
      {stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[15],stage1_5[24]}
   );
   gpc606_5 gpc36 (
      {stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[16],stage1_5[25]}
   );
   gpc606_5 gpc37 (
      {stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[17],stage1_5[26]}
   );
   gpc615_5 gpc38 (
      {stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_6[48]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[18],stage1_5[27]}
   );
   gpc615_5 gpc39 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[49]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[19],stage1_5[28]}
   );
   gpc615_5 gpc40 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58]},
      {stage0_6[50]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[20],stage1_5[29]}
   );
   gpc615_5 gpc41 (
      {stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63]},
      {stage0_6[51]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[16],stage1_7[17],stage1_6[21],stage1_5[30]}
   );
   gpc606_5 gpc42 (
      {stage0_6[52], stage0_6[53], stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[17],stage1_7[18],stage1_6[22]}
   );
   gpc606_5 gpc43 (
      {stage0_6[58], stage0_6[59], stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[18],stage1_7[19],stage1_6[23]}
   );
   gpc2135_5 gpc44 (
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58]},
      {stage0_8[12], stage0_8[13], stage0_8[14]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1]},
      {stage1_11[0],stage1_10[2],stage1_9[11],stage1_8[19],stage1_7[20]}
   );
   gpc615_5 gpc45 (
      {stage0_7[59], stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63]},
      {stage0_8[15]},
      {stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage1_11[1],stage1_10[3],stage1_9[12],stage1_8[20],stage1_7[21]}
   );
   gpc207_4 gpc46 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_10[2], stage0_10[3]},
      {stage1_11[2],stage1_10[4],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc47 (
      {stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9]},
      {stage1_12[0],stage1_11[3],stage1_10[5],stage1_9[14],stage1_8[22]}
   );
   gpc606_5 gpc48 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34]},
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage1_12[1],stage1_11[4],stage1_10[6],stage1_9[15],stage1_8[23]}
   );
   gpc606_5 gpc49 (
      {stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40]},
      {stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage1_12[2],stage1_11[5],stage1_10[7],stage1_9[16],stage1_8[24]}
   );
   gpc606_5 gpc50 (
      {stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46]},
      {stage0_10[22], stage0_10[23], stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27]},
      {stage1_12[3],stage1_11[6],stage1_10[8],stage1_9[17],stage1_8[25]}
   );
   gpc606_5 gpc51 (
      {stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52]},
      {stage0_10[28], stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage1_12[4],stage1_11[7],stage1_10[9],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc52 (
      {stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58]},
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39]},
      {stage1_12[5],stage1_11[8],stage1_10[10],stage1_9[19],stage1_8[27]}
   );
   gpc615_5 gpc53 (
      {stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_9[7]},
      {stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45]},
      {stage1_12[6],stage1_11[9],stage1_10[11],stage1_9[20],stage1_8[28]}
   );
   gpc606_5 gpc54 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[7],stage1_11[10],stage1_10[12],stage1_9[21]}
   );
   gpc606_5 gpc55 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[8],stage1_11[11],stage1_10[13],stage1_9[22]}
   );
   gpc606_5 gpc56 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[9],stage1_11[12],stage1_10[14],stage1_9[23]}
   );
   gpc606_5 gpc57 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[10],stage1_11[13],stage1_10[15],stage1_9[24]}
   );
   gpc606_5 gpc58 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[11],stage1_11[14],stage1_10[16],stage1_9[25]}
   );
   gpc606_5 gpc59 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[12],stage1_11[15],stage1_10[17],stage1_9[26]}
   );
   gpc615_5 gpc60 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[46]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[13],stage1_11[16],stage1_10[18],stage1_9[27]}
   );
   gpc615_5 gpc61 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[47]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[14],stage1_11[17],stage1_10[19],stage1_9[28]}
   );
   gpc615_5 gpc62 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58]},
      {stage0_10[48]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[15],stage1_11[18],stage1_10[20],stage1_9[29]}
   );
   gpc615_5 gpc63 (
      {stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_10[49]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[16],stage1_11[19],stage1_10[21],stage1_9[30]}
   );
   gpc135_4 gpc64 (
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54]},
      {stage0_11[60], stage0_11[61], stage0_11[62]},
      {1'b0},
      {stage1_13[10],stage1_12[17],stage1_11[20],stage1_10[22]}
   );
   gpc117_4 gpc65 (
      {stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60], stage0_10[61]},
      {stage0_11[63]},
      {1'b0},
      {stage1_13[11],stage1_12[18],stage1_11[21],stage1_10[23]}
   );
   gpc1_1 gpc66 (
      {stage0_0[63]},
      {stage1_0[11]}
   );
   gpc1_1 gpc67 (
      {stage0_10[62]},
      {stage1_10[24]}
   );
   gpc1_1 gpc68 (
      {stage0_10[63]},
      {stage1_10[25]}
   );
   gpc2135_5 gpc69 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc70 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc71 (
      {stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage1_3[2]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc2135_5 gpc72 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[3]},
      {stage1_4[2], stage1_4[3]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1406_5 gpc73 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[4]},
      {stage2_5[2],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc74 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[8]},
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10]},
      {stage2_6[0],stage2_5[3],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc75 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_3[9]},
      {stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16]},
      {stage2_6[1],stage2_5[4],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc76 (
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage1_4[17]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[2],stage2_5[5],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc77 (
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage1_4[18]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[3],stage2_5[6],stage2_4[8],stage2_3[8]}
   );
   gpc615_5 gpc78 (
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage1_4[19]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[4],stage2_5[7],stage2_4[9],stage2_3[9]}
   );
   gpc7_3 gpc79 (
      {stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage2_6[5],stage2_5[8],stage2_4[10]}
   );
   gpc615_5 gpc80 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[0],stage2_7[3],stage2_6[6],stage2_5[9]}
   );
   gpc615_5 gpc81 (
      {stage1_5[23], stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27]},
      {stage1_6[1]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[1],stage2_7[4],stage2_6[7],stage2_5[10]}
   );
   gpc623_5 gpc82 (
      {stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage1_6[2], stage1_6[3]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[2],stage2_7[5],stage2_6[8],stage2_5[11]}
   );
   gpc615_5 gpc83 (
      {stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7], stage1_6[8]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[3],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc84 (
      {stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12], stage1_6[13]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[4],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc85 (
      {stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[5],stage2_7[8],stage2_6[11]}
   );
   gpc615_5 gpc86 (
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[6],stage2_7[9],stage2_6[12]}
   );
   gpc135_4 gpc87 (
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28]},
      {stage1_9[0], stage1_9[1], stage1_9[2]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[4],stage2_9[7],stage2_8[7]}
   );
   gpc117_4 gpc88 (
      {stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[1]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[1],stage2_10[5],stage2_9[8]}
   );
   gpc117_4 gpc89 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16]},
      {stage1_10[2]},
      {stage1_11[1]},
      {stage2_12[1],stage2_11[2],stage2_10[6],stage2_9[9]}
   );
   gpc117_4 gpc90 (
      {stage1_9[17], stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_10[3]},
      {stage1_11[2]},
      {stage2_12[2],stage2_11[3],stage2_10[7],stage2_9[10]}
   );
   gpc117_4 gpc91 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[4]},
      {stage1_11[3]},
      {stage2_12[3],stage2_11[4],stage2_10[8],stage2_9[11]}
   );
   gpc1163_5 gpc92 (
      {stage1_10[5], stage1_10[6], stage1_10[7]},
      {stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[0],stage2_12[4],stage2_11[5],stage2_10[9]}
   );
   gpc606_5 gpc93 (
      {stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12], stage1_10[13]},
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage2_14[1],stage2_13[1],stage2_12[5],stage2_11[6],stage2_10[10]}
   );
   gpc606_5 gpc94 (
      {stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19]},
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage2_14[2],stage2_13[2],stage2_12[6],stage2_11[7],stage2_10[11]}
   );
   gpc606_5 gpc95 (
      {stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage2_14[3],stage2_13[3],stage2_12[7],stage2_11[8],stage2_10[12]}
   );
   gpc606_5 gpc96 (
      {stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15]},
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage2_15[0],stage2_14[4],stage2_13[4],stage2_12[8],stage2_11[9]}
   );
   gpc606_5 gpc97 (
      {stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], 1'b0},
      {stage2_15[1],stage2_14[5],stage2_13[5],stage2_12[9],stage2_11[10]}
   );
   gpc1_1 gpc98 (
      {stage1_0[10]},
      {stage2_0[2]}
   );
   gpc1_1 gpc99 (
      {stage1_0[11]},
      {stage2_0[3]}
   );
   gpc1_1 gpc100 (
      {stage1_2[23]},
      {stage2_2[7]}
   );
   gpc1_1 gpc101 (
      {stage1_4[27]},
      {stage2_4[11]}
   );
   gpc1415_5 gpc102 (
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[0],stage3_3[0]}
   );
   gpc615_5 gpc103 (
      {stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage2_4[1]},
      {stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc104 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[10]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc105 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[11]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc106 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[4]}
   );
   gpc615_5 gpc107 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[5]}
   );
   gpc606_5 gpc108 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc109 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc135_4 gpc110 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[0]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc606_5 gpc111 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], 1'b0},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[5]}
   );
   gpc606_5 gpc112 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc116 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc117 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc118 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc119 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc120 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc121 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc122 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc123 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc124 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc125 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc126 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc127 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc128 (
      {stage2_2[6]},
      {stage3_2[6]}
   );
   gpc1_1 gpc129 (
      {stage2_2[7]},
      {stage3_2[7]}
   );
   gpc1_1 gpc130 (
      {stage2_12[9]},
      {stage3_12[5]}
   );
   gpc1_1 gpc131 (
      {stage2_15[0]},
      {stage3_15[2]}
   );
   gpc1_1 gpc132 (
      {stage2_15[1]},
      {stage3_15[3]}
   );
   gpc1343_5 gpc133 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3]},
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1415_5 gpc134 (
      {stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc135 (
      {stage3_5[1], stage3_5[2], stage3_5[3]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc136 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc137 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc138 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc117_4 gpc139 (
      {stage3_15[1], stage3_15[2], stage3_15[3], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage3_16[0]},
      {1'b0},
      {stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1_1 gpc140 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc141 (
      {stage3_1[4]},
      {stage4_1[1]}
   );
endmodule

module testbench();
    reg [63:0] src0;
    reg [63:0] src1;
    reg [63:0] src2;
    reg [63:0] src3;
    reg [63:0] src4;
    reg [63:0] src5;
    reg [63:0] src6;
    reg [63:0] src7;
    reg [63:0] src8;
    reg [63:0] src9;
    reg [63:0] src10;
    reg [63:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor_CLA64_12 compressor_CLA64_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h18dcf1b617481de782cd7001e30d2e3dc040c186334bd799c0ac079188b66f7d985c946d2ede23affc7b8c6cbce6e9db84b8e6eb9dbc0f3c9b6c866c1f84c0370476d12a22f13635076665c5ec5c8cb2efbcdd612ccccc89a0d468df4e72e759;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf14f6c94cf6438fb3cfd7f579791a565a443574a45ed3dc6e3971dbabb0aa94341fceecb0b1fcb759403ecd5fb4046f7471090abe05aa2550d54fd03937f57cf921f620146a610ddeaf50397798a87c2e0a0d2b4271b956dbad0cc96026091fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hedf1db15abc10824d028717d7698ada07ef6f377f5b5ffcde7490b2c557948c356fe120fbc5dc57b40f09dcff700e9de2b21943bf8ed641ee3741c1f084a6aec6c067edd79b7f89d69cf8b4033ac6869b764a67a19bd6afc0cf45b5136cf546e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha7e81c23d949561548ba378ffeb5bcd718528154bc0c3d52ef4899d25bc1df4c5fbd398b75d6911650228057a38359febfe0aec8c450dd04c816c6dfaa0004601cb42ff45b3dfbb2283a6cd854ef5a79da632308bc554de9d27a06d95ed0c835;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h8d8507639f78780f8f32d7c7dc3fea91cea3219bfe09e1197917b9537140a664cae13de249f64b5c7a4286a1585d27036bec50f7f5dc2460acf926ad7dd8c8df01aaf928e6d2cbdc5682a5e150e50d36f5be788a660bcacbc92352128f95d651;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he8d0e3d5f6f65008d70952315c8c71308f4dc3020eeae086925b22a955484c6dbb5164b630596d827851bd77fea5eb54306416a3b3b993cb7c475353fc9da1f36a271a306f8b4450a64002f782182588db016e9ecf61048cdd63494bc65c9c8c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4558eb0b58460d4452ad0608af4268f7976307f0dbe915be8925cffcf3a175b2e6aba730ca6808cfeeb280861711518b287e4cbde9fe55a1223d219415facd229700648ced8f0ab551bc0160e80e59cd523893196a0ec13ad56a95a9b3de30e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7c354f279161ba786f4da25da24235466dd9c6d120cbe972925208839788fb0c368378489e8ea944ec3e32cfcd60cb04654d8b9a7d30091ede6d339bb458852fbdfc8d0359b70c47cb8064a803227c961bc3aabdb69fb64eca32a9a997b03fa9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfc257b0822bbc7e8c47b19a40bb9cfe80a143ec221f52154a8c94ac2a73b7b638abc78025ddbbed0a3ed82ed112411a88d4caedb1771b6c58be9884748af02616cf21bfe19ec73e4190163c7fe47e83cf3188dd52b53bc27528ac1db9a1714fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h823bf21af2ee9927efd3a0e9375fb01e118ec465faf2ba1300dceb4fbfa0f6bf45a8917f1f94bccf2711c4956bff2920688423095ac26cba590756410723be86428e50343c0f1e07b14a4e20b11ff7b0a94d6a097c8a8c502685432bcc8d4b91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hadd7d4c46dfb3f5b03b58a738ea68cadf4d7ae59cb1b32d69df19af61b8d889d45e297d623598b577f262534e5812fb09c34c8dac1a099d77288c5a0b78fa55726c24b2d82ec2b456f1c10e74af10c046fd157cc244cf2e032e2e972bd62f9d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h93c602e9b2fa10e6f7369d2cb422e949af40ca7ebb4da19d7fb83fa7673a0e694616c42bd2a2d1921a185c88db17d50d56e3bb5ee8ce6bce706a676b7bf2ec50a93b05fb1b9c1ba497b0fcbaa9fc0f18b2ca4e5f960e345009156ec0e9c9c8d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h6cebe5f1697849b11a83159de89905bd4d215bcd47600a22d29ce86f177e385e6c49ea2912640eb6d8e01e796a2468ef3378063c2f29357260425c3fffe97833b7bed13e48bf1fcb65a0f6a07dfbee37b2399f539eff2cef3140eaa816a04211;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7dd1db58ae5049f6a1b4935a3eda61fe0aeb9ef943ab982b98e51084c462ca1a055c1fa3a701146e1a1622ec63123eca6fc549a61c236b3082df75e47915376a0526c7c35a0f54776f89c2643b15bbd079bd6fb0affa56b7dcbd597db8c16951;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h47fdfdbe40b8c27445fdc3f1c1d1ed4e38c3ea19b0571d0e12d14352d20bd508c1503856d17e865f2f9116981d98a473fba7c424091c49fc40b7224d536441afa56dc40ea05f3c98f6c6c979340924f5e5330e7279afebce00cccf4d9c177872;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb1626a5d1594437c56277f71539f29fe952f140f5dcc35ddc8dabbcfcbdea64459a4c9f31fc716200a138a3c3674d619b4aca555c5d21a2cecd6ba09860d1a111d9911314b3d991117760108f7c7acb6d613484662ad8ff6a1ffa42a22a07331;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h57e64cb676644b63c67f3f0aae6f7ea8dc9761dc6b548dc507076770495830a8346b205f17476c66ff9f7a0ae8bcd42b1e4c4be9931665a5708772dd28fe3404228e0531ea4a34468ced4ccab67ef1d8942f2964fe4c4997dc17f97a20272977;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hb9c6bac64a2506b45ad4e41b3a72df77664121f1d915d247aa37bd73fe803abe590cae92cc59a81a959840bfdf46d389ad2ebc801af46e6ef73bd0fc7d608b312f6fd42267796a8702ac04d8e6cc4e2e1e979f06b559de47493d84e3d5571083;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd4c8644de575abeb916a456754109c09dea38066740949d0ba0363da9e6afba03407b02f2e96b818bada1991b331f20ca4ad5fcc201b1a3362be1ee889f67b0c39b6cef527d354e53e0c6016cb2c1c7cdf5f1a98356c47a839bcacfce01d0070;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc71baf542a6d1c32dc5532e15e004eb4c12a568ac24366a33189e2990998fa6050e3325f46005e1266562c5a25d3f7e6e28e10ee374ac17ebc4acdd1b9d213786187aa15939e4fcab7a4dc37f48669257f1b2aa980ed18a562f10b0474140994;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h1772517b16483f2cf9a044dbb095a5dbb498f05aeb8684217e536ebe3c74f63dc7005d93356ff31f976a89b853d54f0aa20ed91d09e6c9f86c4eab63c40a405071ef8d07c0f0d61e31ad680f51ff57e2bd06ae4685d9cb366aba6d8d1a6e24be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hcd164db79797119644370ecebe91b7bf6c85bd82fba8babeae4730cdd722514b8dc51250c65c52abdd3822d5dbacf5beb48e23b7948c23351be181d2f78233ebe7dc161e3fb697236d23d3bc6dbf29a041ce8fc1ce188fe1f6b09272d06e827a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'heec10ffe590d2d5a03ddfe778368ebf01eee425d0f4c7a84fdc65964acd4f9ae344afa2820c4201faf1e1b0fea96a79b9aa27338b74a4503d7a1db1c1dd0542f2d9322a20639274cf130ee90f75978dcf7c2c0c45c07a1b5f07144b2239cdcad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3f054442c443714d022604d55083adf83fba4a83e1c397b94cd5b069f9f472a60803142121ac220391d0de33e3852ad2d9a08db7aa8c09a3a98b6d216763a8847027aaced5dcabc43deb025244b6870b7fe897291a643a11d29acd31513cd45c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h18522d6f2b34e2d8a3ac862661eb7b66c7c2012d244f5b8d6f31c761aab907cddd8a29f9918ee3c8f8dbf8d27c2ccd624e188729a47b6909de6976df4460718c831fef5250c961eb3be5063d4ee290c959524c372eda56b33f8cb4a707e4db66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h23225a3952f5e05118427de2f5b7ecfa48c78a6c87dc6ef804a2cfa0db1641c2bea46d450fccd6277197f1c337eb048685233d6c8212e228930ee56025621a24dc2a00147cb9b7acede9b86a6d3fd100251e6cf9cd910e3938c81f8db2b05cea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd7dc27778cfa233c9e699891032ad481ac14d0d3eed147abb456a0b6027302e90b74c21845f209b3016d16f273a54fed5dc762fe3dc99798e8d4acc7bac133a4b8f55b4fc3060dc5c8358aaf23b9460de38d56457daf59e4f6bd815351bda8ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2a3dd48b7ec3bfb9e785b084b311df8961c2c71c792de8094ddf455b7159f7f042127b2fc2ce90a1bdce936393b411df7bbf0d0599993bd94fd64939dc3cef7e0044fa180add705e58cd9c3d5c09d06eb4233954af49b7a7ef194c831d719d1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h10503bd64286c9ba61c681f0e1a36a25d1f01b73c08ed03e406267f50f050f11030301f8be41609a348f34463fd5ca1ef321eebf17031175681dea5ccd6f9d529a9470fd459187b59f9ab21b55aaecd840093d0c4cb2a34d6c291ec98cc843a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf719113d3acbc6fb3ae9c4a781b6973d5d2cd4e1085cb95966b76a9c1f343f75b52b1aa21b2c1f61e05800bac2abe43bd9f1c2bff118309ef92d06f3dd2726e9ea9c2bb18714c91ebd666fbae3b6711656fb1fa01fe9f36a6f572b9723e27881;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h657e36e485eb19a4e4f16f78dee3e5dcfa6255033b62e01e1fc2cb85815bf67326d929825bd741cae84a854ca1048708eed37a003b0d5e1c70f893964cbb31c9dc30bb143cc63b65f3e6e289343d6f497b71ad2f42c0ccd1d4663efc3d8f88bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha4552b1dbbff72851d04b9ecbf475f3ab712cb561ff723c16aa7ea70e2765314405dfa668098ba1cbc3bb9daf5df508f8f79c40f74da650217f0c0d83c52656e899374b4484df1fd81a43f6f60faf12076b10c49db5f6e653da2776cf73640ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h22ebdb30d11a8637a547faf2bc138317d43322202bd910a7370793cd2fec9f84c759444d7a18655fd955e4792a45e5c2e0b053177f6025cab5518c7c5d2a89293b3676167a6ccf9cd2147d5984f6a4776faedd7cbd3f81b7cfe442685abd5563;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h919f1c1d02ce42e7578e61f65bfc73688f11384de05f23b64cc01bab3dd601a685d6102c1ef26c56fd3773ec939bd370ed11e73ae1531babb214ee18d385b764b80e8e1d890a5a6136979e05da60f1f824f52fd2de3b04d736d7edbfb9ef402a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h78dfa18e427c67979e05b154f9bb61fb05872f8ed50f283d57345d0b55db477cfd10208c0d60b554908e92be5cd60f73da997c4d8fbded2fbfb39c496913838c397fa916b354e09f723b87951719eed726f99e3f2284b70ac04986771490035f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf8c6038b93ff43d37e013ceed7c17ee11f4658f0f14b43ee7bab1722c585c27c401662dbb3ca74d930c820b406701c4d5186773956bc52d90144e6f89295736b274cc7ca5302a38040287d908783da9406472d963c5f5c277393c460e0520e5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf2228c2d250e89d46e74a0fb9f7bb170f2f362a2f36e7caf7559cd49510c8dc3337aef30325fd1748224e56b2b6d2c46f948cccb13ba76fa31de373c07cfb0d13415e4631324ef7d1de39039f3ccb73918890b4e205b170d5d3656f0678b5bd1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hed3c2bc7e1f770c27219e5f5494c33e9e6b2aa855efe6cce53b65bab372d1d50e2905adcbc9d7a468f6c4c76f4376d7066da18c8e3808d6b3084f6fb64e694ce1f209a566b7bd75bfc3028bfac61b3a9c98c5c43895fae2a20fcd2266d4a48bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3758bd90c25f2364e55965f2f5951ebb40b966109b9209f3ed9d3d244a90f62730582c8d1c319cc6d22160896b50f6fc8951bcdb96eb461a27f3a1a16c53694cc6a8a03757f1303af09148e8a4e5eb271a9f1b5d9005873747f01d0531c60065;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3c496ef7745e5c661ad7fdc8c561e6d0b8806db33246c10f6f87353280166661d62d83c6cde0ae3c706a5593a2469414ee7a27ddcce5c8e7a19f94fc4e1cb6cceec3af8febce4f0e0062e9b28d86b91179b12ca4582e1d6d43076dc169eaeae3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd10c8b350e86d5d443e78222daba7a9a6f76c074f62c4e46a1cbefdd09aa38a9999aa2a42cd0fd03182d9224e7a2dc3d1f5f6e00f7b220198d3ac790a5a460e8770e573aab0cd498fd7edf1d474b959c6f17cd8b4b5d295458e85a101deea58a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3c0a37848c2a1960046b6b030c38bfc47afb8346de8b69b4c75d6f2eedf0f05976137646aea5b972ba6a80fdea5f620bd7444c2b33ef828b1ac19af26f15319a68775f9654206f8bc79743ed5d51b0a58fdcabb2cd2ed1e26857df397a004ad7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7bee78bdf8a5b5e25c256057dd4ca2eff888843173e60ad5c53fdaca37e79e9cbecde440f6c1a7575f7c412d7ba0715b0dd76e634d0c4ae31e98c08ebd05e549e2d5d80d1ba346a81d383952d5c4a0a1617ead3385b209a7ec12b82244e08e05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hee0fefe4b7b1dbabcaf13075caa1ecd925b15f7b8a964a6b6f6f255bc5705f76349c1db7134fc2786ea0000c16f56b80c8a9cae6a19b0e7a47950fd49b745abb1efb5306bbf15a7f0fb4118b7992fdfc9d6e630e72cc622729995838820a5a55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hdebd570db98b2e05d9349530de9b8bb7bd306298ad67f2136d0b4eff438582c0f9c9632289d18f2697d78b97986384d6404567aa76497f74dc82852d2037924aabee0be71ef34638ac6452d3a4be4ed994f2844876bdc37e5751621df6e3c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4212885ebb2ab0512ffd1798df1efb74c84b09c6a1616194226c62ca3cad9e48822a699272e290613dc0258e72098309a51775c1eddd7034eafc91680f7c444e65c24086a83285e56fba642d6265a61b7cd38fcc8f587e3b70646e79b901590e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc90660bd73b8ba41d7c3ba14620dd9f348dd56c7bc666026f6483bd081319c2c29ea7279eb2baa9b87c8541449079b60b32de336167253a8fe3907969cfee87eae20351199b48b9e9dedbb149f3a943a84eef65b056c92a5c4cd7b3e82f569b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'had707318f5ea32797cbcc8f1fe69eb1a0042636fe4cba95bb6264df8abc42e0f60cb773b6b8f01775a1d8439fc44807eec9981d97444f6e183c7790c33110efc2b4b5d2e26c19356b2e00d97465ffe741b4f14b8e5ce673d7bc765413bf6bc59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h728adf2bc40243e7d9aa9e2252d8f3b7f46b89615958b8f6e99528834f3d99601e39389323abebad61ad3b0b0adbc6ba7836ebd47fdc45c57e632e92e5ee41f2c8e2dd69a876287b12d437a9db881daa6b8fc1ce4fabf56c18a228ad365d0afd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h81913c5c317bd03436e17a218c37c5e78c698766b4836f30fe788953b28112e73799ea66f0da40fb86b58f5c674cc608cc4989ca9f0e5f4373816f9d9224a2c12a2c1d0d3290f52b023926257f93a7d5b7598b5ea07dbf30d1a94b234336b8c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfb5ef2bd6d076f62ad453eb3bb2c247ff5193f378d557de2544cc79fe79641c73e01b7a9559bb0871f59c05cb587cd642af4fd9dfbfab2f87307aa1d4efc82468a4f06d019aaf0c6d2009b9a24f9821af484cccceade9391309a1d2d29c8b8e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hcf3741ecc3a229f29353a7cd2082274ef8a8f04c3bfbd7021a232b9289573460142eeaecf082f0b51efc3987cad77c0f1efedec4b89f05406d5ebfe8f2b7bc1cb964386655811f06d2f693e58441ee4d6236440749d663a161ee7ed4aac8ed68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h43dc9094ef2b50588d64256475caeaf99cea2324936ea97763735d0fe85df4dbcc63e5fc7fb2a9fc40b945e142ae31a2a88106e5f448d78ac4a5a42d387c9b59a5ab798513b2dee7153367db3a19daa68736cd6d63d3c31e302baf79c8ff444c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h54fa6329b19941679b98f93d4b6271e9dca3550b92817b7ac58dcc3b1a35b55529a1acfbb1ff97bd3c92229be071684e6a16171b529f1cc6b81d398466a908071a84d24bc2663731cf2580d4802bf5ab6c37a8f2c40a64a563846c3b0ff97340;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h905dad5ce8424821d5c7922452f51a91e64dd6394546c59abf2381ebc177d0bcb5c50cff3527283acc306252806ff1a3b52a60888972f69f58576bba7f486bdef7abf48b20f33ff606cab6f8b1239f0b6ab7ca20645e5e2455c3ce6452d60993;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hec88e80204dc815b211c97a495f7578e5c9f06c25562f6c254c8505bf4074aa03913438c563aa8cdbe90a1a45cab4a93a5d39e947e9798fe9bca59d84b4d1b263593d36793d7a35797f87c2c800745844e10bfc796befd43b492b26736f01dd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hdc31b702bb089e81cf9faa588acbb05ece5cc15f24c759935ced970e76d71ebaf82d23c64c081542d6aa4a135410b02985d8e9b18a3bf8c1487790afb1c90ec55033ec060b461a0f490d83873f807007e8fafc733705ff3ba622da7a9c8d9dbe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4110be244e92cec771a8e9f176d2036f4a032e23e92d65b7093bc3ae867e5321edc29d3113c55406cfcc7dea8dd97bc341ddb152a0c517982273dfd4590ea43fec74bf9395de9e1e5dea3acbff9f26e1ce96ede9ee36b7f05b426eb1e93df79b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hab3654369a9768ec8e194198752055cd59c0141ce64d1e6c0920e7c6a937277c4c499f369a21f0e82ffa9c6cccff510ac0d626e76444665ef0d2b01f7f0f2a254a9e1fd22d954b8065d03adadbf6b065318fbc89bce7fabbad6b6e76a002573f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha2c934a7028b930a9694dfb35744548dfd1fb8d1311bfc99fec7fd1642352d7deb42234598426712c44dff1522bf9c90bbf7c0b5d2dcedfdcd442bc010441addbf87901e4dec6da2299629932b806e952b1b6d05a2645ec79a7db61b3ea778ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf04909ee1a4419cff4a4a55861375d589fdff208183baaaadc73979dd389b4052ae631d002e0cb3d57a39e3253f138c285a6bd9c6bed9c50f6ba8a660c894b0287fd4e16aefc910994eb7177f72a70db774a39774aaf7f6f0048949bd71774a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hc1344babf1f6eb3d4ed49511f83fa95c61fc020bc244fb757be06f7f67ed782b44ce99d617fda2071b22634b28a3e59b46abeb7b62d45b655cb48745d06550118a42c3ebb18b50f38fc845d0854f39469b43e4f76a7679e75d66046f148091e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hd8b905abf0b144bf4bdbcc669fda637850067707c7ce26f216c8ab18645a04721597b822bee38e393821676b3e4c7cea26039dcde9fcf20f02fbd80f82fb82c7b8ba9b6035029a2e8c88a6b6156b41d8c244712cc75d62de164a18b6896c9bf4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h9f6e1b265c05e19b11fb97c0d241d03707943e468bbd7baeb22444022444547976fdabf731980357f219aa928d37f8b402352f622d08ea6e6449ad954cd3db29ca9c013b0d63728d54624d51f7df17bc7a7a64086378e32196f20cd6445bd0a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h29559c581affb4dc92cf01b1bb7a696b815c04770da530da670d24f4141314f7cc3476fce64a62729abb302b3a8fde9aee8fb576585485eabff4d50cc0a5d5c0a17eb55b0a28861614d2c269c348a0adafef76090f5f36e431d19af586d2a9e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h82acecf3d5c5e46b52a01b2f676269193e9e3f906fb1b044c148ccfa0c21be035714939fa09abffc5105ad1cceeb914f1fe94af259397b976c7987dabd170704355a735983603fd9da87b3a6190d35146dac5261a5344280c17dc08a08b064d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h724454827c0075a972e513b3e26b6c91a7dcdd89adc84638b9122336926afaff78e8d3349a7db2409fe06fa6454e76991ed7f955f1efa6806b57bf9b9b98386ec60fabe6fb7e2187cee49fc3106c584dde3858a6ebd4211f40600e2b87397f7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf5d13e534b454d3326d65c19acbbbfe29df91ef9469b85175449277710a482bb51ec1f192365a421755c432afd74ca278759fec60789a05ececb84c81a494706c3f1e242ca6592a60464d1874131bcc5313ce918ba69489c1f32f04311bcf9dc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h2d5c5d15e25bbaacce576d1a3518415f2f72c5bd9a3df5f1c20eccd7b3748c00267a605b8483c7a0b4a6f381a8d8f02abf0ce66bf86072d9bbeb4b07ad9df55a81ba8f30bff5ebf97805f86714f115a69ee0d0be00a5bdb5f94422ce895a5e8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'he58c37150c1c68e0c52034f86975a591735ee39877837ce3dddaa335733f52621ddf4b06293c29e6daa46e98d6bb88305f097f7a30d9de0a970f1b372508effaf3e58cb18cc16af5a2ccba80e56ca7397fdc04566f68600e6f9efdf15bb27f67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbd1acf1c1d5727828c78a7ab7f1f9a28e9c75d7e8c9e3afe4ad1d7c1405a88591fe9a56009e1b1ebc01649401d1664d3e4b560d1bd48917dce2b59fa5c84f1baedb342451a8e3bfda2bd9f3cf745619d27d0dbf6ab06638b5eb02a069c30058a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h40f389271ef3cc2dcb2e30417901e46ee743802d93560afb31960c14b1a1a3c14cae9d7b3543804229d83b84e0cf51f89e7ead98b26aae48eb989f6a148081561ee8105ca68543cd91e830a8722fbe53d9f9501a6c5e22ea29ea3e5daf1f6dde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf09376232e641f81544b366b593aad7e1f2e48b5487e094701d0b3005fc358d25407d44f3634fccc34373c7e49034cfb1c74ab85e9ac00dd7553c2813484f476c798effcfb584054ed0dba7aa75aa790f8f99486bf2155a346006be0891c59e6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3bbb6efa68a31e1cd6d4928599023cd36ffd9a58e64451fedeeb434ae853ce9ab4b16ba19ec34e5b80b4c6773463e203ab494dbee56889db4325d82f9e3fbc474d8b2bcea9176bc1d5beae780a5fbc3a115d07e59c6bb5500e7b4b3de444d868;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h1a5f02b902d8b1af07b74835c906e87979a50d179dfa836478ff40bf9ad903ee5e4a3b25506ffca01aa9a53476132b057a1326ba4a96162f0b2d49d98228b6e74397a81b13e9771161a14c9e51591cc2172a3ecae73baf3c7e50f77a7801a09d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h85fca2a0a5955391f7af86d79a5fa97d7da1e1799e4b031ff1266002cc82d93223bafc9514617c6e35e538f359336b8c766e516ee210b06c2db9874702871c8c80b6e22afbd1c7db5f110018868c3536dab53e63f11d29cfa2f62995c22cdebd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha5cc391cf031154d666110e39aada67464d395e0082e3dba202b4a4926fb095f4a28b6073001745cc9fad56734481b0faccf2d26278c435d948b7c462fda606fc1a4257fef820ec87b8af72ea3dea5891dd272806cdfedc4cc8a0a1abf88d08f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h20d31fa9bbd4426e5509b137b925fbc98d2fab983177299a3b998304018895659b9a1394aad91d173aea96328ff0f9f4c1413b6d801698e2d89af5ecd3210549c29b55b59145e681a7d185add917702b141ecdd5f71a2b3d9d22140a62d91fc7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h40e3be9bf0edb987cb5ba52ac7cf476b092caf3e07c74d1441d5a138e04ba293c996a98ac4ad3822b04c2fe820c2774f5e090426cfae8f4065b7e958c19036deb9e64f58b5934e5e4145b1ce08416a4ccaceba50d541cc30d2a63de1835d7008;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h37a74d4f1bc572c0fa97cf4d11f47c3fa123fb7b03cd30411c89b9cac2a1f5350c2ea9ecb4f88dccc2cb2a57e448ffe87b65bc04717cdca54a1667cd82b4dbfe99ab02d51e266eb692c0d63668dfa411305c9d86fa74f8680849b5757da60a04;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h4c3ca52b027815d5c950cefe30d97384f9454b5c6104208a39442ec93eb43fc5e9cf4b60d995ecd0135092a030d36265687b6c0b62fc23c09669bd341e154d0b31e83b3280e9b469619baaf2fd0b77938978252d6d35ddd981602aba3da9d8c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hbefb72506658574f6a639fceaa09df0930069873f86c448ebb10c6d98e60dea9f421b7df45848bfb0f472ca51f2e428fe666b637f52416222c2717b4767665f2a8512195bfbd2da8d5d8ff4523dc3e5ffb31f6f1d8a68f47573a957e63ca76dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hff4311e35bf91a8281e29ed00c83261b7ec4df68c54f69c416f9f7300e62f566ab8a95fd4d0c5188bbaf7973279b7a0ce0cbd944e55ae8add3ece1dbf9c60b6b475f66cd6ae659b714147a5b0f284eb07bab5d7ad34fc04e8649593a833fc097;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hfd93b6412e2eca88c49592accaea58d621a9a80a30f250e49e4e7d97da66d4dc17aaa2fb0c5d7114130d15416ade58d218d5338750be223ffd644b4aaaba94f0971044afb7a16427fb4f541a7061e73af40e168e06be6c9d542b8e7d762f569e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hcf86533c8713bb211c451b35af8126976f2b4a018a73e64268e134c0627e42e2180c4293299395c7f9ae3061d1ad58d0cb422512664ff8b2c582e87d3375fa34bc7eaf6ed34bfbda4f9594441b5677c976433e87fb33d7236c4caa3d761f6410;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'hf53eaaaaa8e8fe6099fe3b6d3f9f15c7f511d43f7879ab9c6119714ac37cac137c7716c4e8516f1016511f7c34d46dbefb6f1f3a227f7dd4e8ae091e4f05cdba3dc5d81254840cf9e8e3827dc5ff3a94a473728f87c736cb0d78fbd214ba225c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha739202f2e2c7c68a8458cbaba4f0a0302b3e3795a2aed9af71d5532e14a7f208b330df8a47a24550158af28f34071bc781eea9d5531f2e3e56a857978d843264bb7c26684f9d362227953dbc816648533a07fdda27fcdcdaf35d832f0059c99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha14ec6a27fc73c169c976c1d500df03890fcbb01ac43a9e899474c92c47ef473cb7c54ad8ae466e3fa61352ef5446cf235fff4fcf1e1c8375416fa6d56c086901f1d36be8e079202a1f6ea738fceac6b2bebf84ace5072aac956aa5e1615a8ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h64efb128ddf4d0fe48c16889a267d41acd0de8a28e1dc1d9ca62bdc9e8b65288cfae447e5d19d29a8ddbca5f4708e0670d3583da6c4a261ad4162ae674f170dd620a4db3c106346789ee154c108119bef93fc8cdc213b6a221d8c32e062de9d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h847878c031de80ef80b7c745fd19b7f313ac2281ac2ba681e7bc52308a2508ea63eb4ccde01ecef85353c719aae9eb7530ea33af4638e29ebde4545faa713db4d604be8889aa86379054a85d15723e2a2427fa7b453e07a8cd98ff4115eed0a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h60ea3498713bfa2d2016b74a5ccc7a7b1049395aabea412997d95ad268e0a3aa9d0e6f497105f6a3d4555875091189120fa42bf8d5b837838e97e249e2039621b1e21d993d2a50a3e490d58e54aba927b81485391a8170ab2c3bbc4e467106a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h1181e0932de808f155288016022a794336932317e3377d236a06da2ea95ae7230ce39adc2a217569a7952fb8a0ee9e163fd2e294947d5d6fe06e1604bd6c889a5e9c770d7cd34a1562a41c2b48a203c534ccf033c3341d04cc4610a96e4ee661;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h7d9e1940f197d0ba3bbe2e236f6ba6872050ab0ca6c31dad575b0a9a56f33c89ccebaca6bbc3e18a5e411144cc676106df2aa5e239cb4324ea615d9450b6e34d9bc72f39c0f42417209d879ea53bf76187f98b0f0f312b0fb00c58e0cf61017;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h959c2623b99449ef31a55e1bd8171e5e69a01ac10805016c8c3ff445f3ab082fe8ab2ed368b15efee5cf681c53d8581e167823abd1701aae4ce708523d029d8a11d11c7d2de30bb1f6c0284fc01bfe7519071aa1355d1c9ba68ab676aa3902f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h507377a7c119e6ad549fc26950fe3a409ec76e6f658192292a8fb55b00094484922b5fa7146c7ed4d3a80085f19c81dfab7fe535cb9125824becf8806411aa3cea236d08c95e4bb2f0ebe055971baa6947bca76684883c42aea2db170ddd70ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h91de047615558994c91c7fe28e41d6217817414446695c34a974038950e27d856bbedec86db6a88cec95427fdbdf12fe6f44db3b565c3849a81ca46b67d1491cc9f6449932d1bbf9c09aca07bc8b5168f866ef82e2e614d7fd4dc1eaf0b25d82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3daed01bdc02d09183d815f932994b79af30af07645a59d8a9d839cae66c62d89d37cad1fd2e961b2a88bb792c8819d85813f88e91324d24d4f5fbdbfb3431ca0cfbad1503ba306acf21998bfb64a02de188ffe517d69932088ee1afeb052b5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h3f32e4c590147199ce0beb161c8c33a8884e8f9ff01b69b934bb722f7d3f628f5d0ec3b18a983d536eff181dc1688ce429ef4a2a6d604a397aded546b8191de18d3e7c39240808ed74cabbc42537ccdf4a3b6dbf517c4cc52ccb1cb98d3297d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'h97f1fee61980c376dcf615db471487f66bcd99de48f45d2fab3a53fc8bd1a4474ff18232c1856326370a38d83e28fb08ed3cec26d15c32370c0ee882b2c79eb357c53363f2c467c716b18290b843ab714437547c553b90525b3e0e122d7eb04d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 768'ha45ef9bd0844138a4b8120771bfb2acf12f00714769c641d1ddd535c796e74892b4184e081bef1b2ec7c576d0b2887942258494dac75cffebf16765867402f325b3c7cd943aef80d4a073c55c8dac8b08fa4aebe9ee367e9b75d584ffa02bef0;
        #1
        $finish();
    end
endmodule
