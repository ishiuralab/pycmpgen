module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [25:0] src27;
    reg [24:0] src28;
    reg [23:0] src29;
    reg [22:0] src30;
    reg [21:0] src31;
    reg [20:0] src32;
    reg [19:0] src33;
    reg [18:0] src34;
    reg [17:0] src35;
    reg [16:0] src36;
    reg [15:0] src37;
    reg [14:0] src38;
    reg [13:0] src39;
    reg [12:0] src40;
    reg [11:0] src41;
    reg [10:0] src42;
    reg [9:0] src43;
    reg [8:0] src44;
    reg [7:0] src45;
    reg [6:0] src46;
    reg [5:0] src47;
    reg [4:0] src48;
    reg [3:0] src49;
    reg [2:0] src50;
    reg [1:0] src51;
    reg [0:0] src52;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [53:0] srcsum;
    wire [53:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3])<<49) + ((src50[0] + src50[1] + src50[2])<<50) + ((src51[0] + src51[1])<<51) + ((src52[0])<<52);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16291d0fa3a763eab5be48b75270dee0c2ae2ed9752915304f75d61a22392c7981783f16d191fc65c5d57fa9313efea4860fd0da4306728455ecc3123c12139ee2a3ad0bb9241e8e472b3d8e65150b34bf051ff44e6c9915f5f154f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26eb13c1356d11abbe40a7a99cbd4c4a0cf23a6988c68053bc9553bab2f1f76f97fb112a551435ced2955f88e3d142622816977d170a8008c8b1dc1c2dd1b913e605a8364ad99b65980e89a760a56b45347f3e16bc0b9796a9c45c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46fc05ecdec3b46d3c55021cabe454a5b85d8e6a394cb3c3d57aa7e97a5e9b7db1c78c1ba8940c3cf8460503ac21a2bff8bec77282e6860b684bd66c35e9b923bb0b49bc42d6ccdd5eee85d3c26ef7e6a88ad5060e3b4f4c4aa16c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2ef5bf7c1db9a0bc98200809977038d7af4ba638d4d0bdc38097404489cc7c4b0a7db8c9da76b8ff63f4e8c19e1e2499bc2b7f432517d81708ec7ef473997d61aa2e0eeff1ad5ddc9e8943f0c372dd990300bc4932a5b0e72efa0e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38d7b06467d0dc3a919e497e8013b806cabd0935e1535e91fe21f9f7c32fc981590a486f19354f9243967a83305da880a0d5d0110c10602d9cade4eee9ec3d157393f41d77c5fbf8af158f8b697642e5715a6a653496c980810177;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae8ae5d48bf24250f74f702ca2e26ef911c648d9584e2862d708b4db7ebed3b1d901e29c653138c83010e372c0b20088c51faab9c252eb7e8f04b47ae3eff24c1cf36d83d014bfceb62ecd176ceed6d846d9f303f3d9235e009afb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15f0feb57540365bda40a2bf184b6ed525460ea9df2da1541ef7c41e8e66cbb6af175d6d6d8fad07e6f86fcfb85307c910d604cfdda29bd236fd1cd489f5731d48850f584f379a47d8edd9197c891a93c117fae8194413782e88435;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4db581496d9e2aab166e77bca5d769d690fcc044a77386808524da1470038dd6f92425aca76f8edfed8450b60f4afd7c6abbe5c6e5c1badb68a42541377105803f5a4945ebe257b4bc3bca0b249ba96e3f857b1bd5209da74b29c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h407ce967d0b163deab9ac00b103f43e5aa6be1f850dd80045c0deae35d3677bbf31f06af1ed4199546e8707aa0610ae04fffb39b2df4d58da8e6855cf371800954670a1c3f748f6c87032da31df63666b1c728ea308c46e7a491a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1297e6c78bec54ab6ddc2ff263ceee13c9f7291d880bb15580068374e49f4a3881bf8a0089aa4b50f5973bf197c4e0e133c6012e1ffd57cca554ceed5f14ac2326c4226792508d3808f70712522a5f3bd56684fcf37d5a0796a4749;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1940277d9f12a3f46f021eec9d80794dd6b56bf08d0095b44ab27587d114d775e569ea7179e445cf89b983a83098ecf218c10f85f247b7c5d9aa9f05ca4c24435209ef6790fab7c435954016dc4e1ce258326f2c4e5bdc6dd5ab500;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177265ce7f6d8b48f1ec06384002d460812936eafbd71898032002fe372ace86e917e45d4f098e01a7b21c1dca7660a5b92daa7e5a2df7f3651f38cdc8d468cd48d89711c69783734bf8f0ddf83b542fbc1cfb69f6b6de2ee779ddf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4101f3371177d6b0f421502f45af3635968410b7b75082cd8fd53f5a5b0550619e2be43e5e198db593d897243d2dd25444e8a91859431d00dcd88909320ce837ebeb1893255dcb56a0ef8f12d9e5829d18783150b4d2ad669ca6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13dd279a43c99697bcdbb7b4c934493a1acea62b3497dfa06d56d00dcd9247d2f28bf04da77fe303004db12fa0076637a06573436b3e0994e6fdd4ecdc5e5d400a6283062b43c8d45093d55836169de455e9cca502ff2f4dc9e1bcf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f522fdea4479602b26c4ac35ac32c820cace67d0c4b0fa07e5d8050c5ad68fcb7748d15519c683fe1d39d9673f043fc7543bdcffde69dcca7ac717cdabadfc7a1285fbb50c6d44bcf43010c475e8dc53b5ad743449a9c0de2c9f72;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf99a1abf3d21b6497f43f9e22119364fbc5e5aa7aa208074c57540fa2d2672aac78716ab3257bd8b19c69fab63495b8f74062fa2c5d3d8c052ade1aa76efdbe8d0615ddcf44c50d70d89991f9bc5a95844ada89f225a4d8f0cd6f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he40891b340e0182a36f53eef3a9e93fdfe315e7cb0c4b1349d4aa4e6dc3958433d0d1e56ab95dd6d102e17aaf6e2c6904376260582f02e582fce23c6e2784abc746932945b6a6ca9b1e7b139d17142733e04e9fd8d0982a0798c4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfbb497010a038439213425e16477e4a8bd9c6e3650fe0d52e25bdb33a0c66961316461f8056f68f4dfe9883cfbaeefe9dd17c5678e5d7d136d218ae09795b8b130ac6a4446538dca5d542d233a13cfa5969d05380f1a5bae5abdaf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h149a5bfb90955dc4415629f4cce11911fe524da316bacdfba916dffdc276ef3b06faf062fb18b1aa7d83339e961a6765cbd628c89fb2290807eebbe11d2bd9c6b511a95dc0f8d7b0be48d073a6c834a5b80f224e00d957548e7c239;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c21aa81e57f6d2a449d336b9afba4bec47de1103e3a7fd1f8e7220482932dec029ca1679a297c241987338db93d2aa6b6f6298fbd520e6bf2627ee9648419700dad0c3494557732677f9582cc0ddc5dcb0509df390ed7fc93f072a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29357d676bff757c3752ec64d6e85098a16d9a6e8773451663f3fa8712afed5ebd5b662898a7144217453dbbe7fbfad74ab9075ac8fc590b689cb601448ea0524a7d3bdd197635d15f14c8a889b15f877345b9e1f8b362bbcb80ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4548d4e0580bd66cb1f62910402db473a13ac1a7b366861096d7551f02f1798b98a0006b423c43410dd440c842d23840253c752d012ad1dee5ade7f36f78331daee563ed8aa97b517ce8915be59182f69e28889401b2d37983c877;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c64ae51d17be8a10ee876263ffe609b08c7a09bc1470afef2b4df964fe7586ef7c00c833a5a370322690914cee4b0ae085c8e4043531aec30edaadb9d1733d81720796b7e8c5feeaf99d283191eb8a5d733ede2e9fb6972176324;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5a3c149e9dade3ca942c3c935d933c1668845742ef0ddb7ad3db6ddfe0331e4e317d1788206c49bf2bc962198335a83d4eaa2bb9a6052c0105f8ad3fcf1d70db39b342b5eca4c31d27ee711f61f6bf197032bbc75550c693f977a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e04f8eafd99c4d6e8ddd7d03de78b90e12b0b1052ba5b9459f38db6c957ed5ac87a902909b52ca5a6094288dcf15478261c07ea8b626cfc1c78288b9cddcb14d987424745335b3afe7d4c72c52b29c2de119e9b365c21d95d724e8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4f5fd91e569f4ac97e42dccbc887fab184d9924d54fdf301474bf5f80532fd8b6a10964a2c8c294265a362fa0de7406a36774cb98bf87abb197c3afb872d62d50b4a99d90dd46793cb5b0e65d74340349dbf1663bb89a4b804ac9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9ecad7abc5fb01adeeed6ae483f9df4d6033f89f9426cdceb0930bda4ae865c806334e521b19fe9564a9b5bbd139ecd994a2b77d678e7e723c4bfe839fbc34fad920f0c4527a591d217e96af5591af691e7fd5fac0eb462f2353f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h181f6f84257b0d9a80209c500f425d5c853abea594994501ceedf086273f91f9024ee523c942b8c42e282c99e0d53d66028b29cbc58db350394031bf73cc8941b555e1193f6a7581aef7bd1c013238de1abfaffe1e8e3bbcd628b9b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c96898c11c3566234800a00837da8d7b182ad560b2c3c476f7b0b27548f8efe037dc1fca0a97c1b26c2fef6925ad5bb889b74f124d0243696270ab596db54b3a76955a5e8c3238242fda238142a8ea6164e214c72c8b6f598abe9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73fce1e0c860cda9cb21a10b94cdae8f1bb57d744208da2b11f75616716464f98e680ee36cad9e4e306bc2106113c98c6bdb86fef7faa0c8a4e4682ecb1ba11263c663f53f876d0c72aa6b4a9d9ffd1ad1251009c21e6f56014064;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb8d4e94689aad5ff2b4273213de4793e094fb3952a738c7a4866df382a41cb42025bdf1368d9d21bbf0535dabc364de06d2336df1c8a840625621901312635228fed9cda9b49ebd5c97a741b0ead7c54a1253426cd89317be7074;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1186cb38e8c70109f7a85ee81dfa775d833ae1c85e485d355ee92c1abf4746a64a0753b9226a749dfbe9d0d2f2abcb8533fe7f4cce5365f0c12ef3bad972f47a7fcba542658b0fb1c83ec6049b0360aed4b362dba7689dff8e7ab97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5a6340ffadceed7c5d65d17424b473732d35ffee0f7f32f813aa3206b3efce3fd189273359930e3c869c773f7ea0f1388d4b277b5bfc37f195871e3ac11921c58e181ee26c3bc7c5de44e3367b96895710c84ed2ba9e91968c8d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19634fc94d19adc7bb42518e9c0f87e642f836b78409eaba1da8cf216d26286b48868de7a316ab8f682e0161f5deb120033bf793305dfd254cc89c96fbe1a1eaaa28011549c652da715befbeda6e5aa06e37a595dc872c0e4e4afbb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec2635530d0d791494f463d3a7c2c152f53f17a06971f295670656e01a17c6bb20cfb8e1a66dade1ce88c8e0373fc880abdaf5b37ba5b6bcd09bb2e49672054e1bc4ce08453da5d5dabb7e1d00716da6876df70279ad42864e0788;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143e6a41d617c13afbf8b91a2be23d108f560ee92d50177fb474d7d499d5647006e3164755c195af63f5284627df267bc5c436d4e20ac688c7e85cbcb1392f2b1673c34ca4f2f815a4a7f703ea09e7324d8ed6997606674b00b4154;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1189094fb7d9ad432ab02f33d51d4b8ff687728286806c6aed4c5e9cd6a873a122adb38c023085325c64e8c483ac65413aff725815b9d6a5a078767fd6ce63743034e7edd211e208030378d09408d0159c6080eb20b873ded26cbd9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13e788c24eedfed14cd2e83ad9ee86bd2f08533c6147f5509e3df8b5a9a38bf79d35834e1f7ebb8ff8dca65c4d074653f8af9129ff97e5b0ccb4ffb7f37a275bab13450071202134fe88d049185aaec77230c305844f384e9de2aaf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1673bd9ca806b6094885738614fc5e9d25aa481cb1332e53d1883d45c735ca1d8b2c3b9a4fe8573b86796eae9325197c2b90923fe4a1af2a5700ed0f9473f25b534a048a9e357b0974fb9e5ec2e356170546b1ebfe431ed4d326564;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc7cac981dc2597d21cb44dd01dd756ec54c6190dc3b2eac25489f9f9b49f3e2f409efaef26a70f8cf2387cbee434bb2f7cf1310eee92ebdd3558fb014f830f871d53a2f98c0ea02747d69dd15fd9c7bb24c3ffaa6510c07d0e16f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68eec56f9c80e2be08b44def5ada43486c213a3d339c9a26aca5ba6ca3b686b63f784a14250ce762e2c7456c52536da1119d782c61d3df97afbe27269bc8c541f934ca70d1b0da70bb0ca6d8a5c92cd6cccc9d2664eb9df3433bb6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153f08a19a67289bd533d4a05f4c19f853ae0a4b003ff266d89f7a87c6fefa7281debcf92d49dbb9fa34b7023d585e7bdaf1a43088cb196664fa55d51c594f8a87a076a3039427c6c269756bd392a6ecfec87905f27e45ea5b0c4de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13cce14e8c9c2b366f53dac79749c571f24e8b11bf064af2cc29b68c581deb883d265404bea0952e98502a95c4bffd63ff9a95802ab71d8637d835d6f83025b933d7d923786150eb27bf15bbe9a4d2913438327bb4848b2e73323c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e508f0eb5a660de88c45bbe4edee9b1593b51b74ffbede001fae1b18b00fd6363d88049d77de7a8695a5b28d4d5d77d0cdbc2147378e68080f69245ab26127b639e28239b1661272214726941d1e3d401d918ccfefd4faea1f4512;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e5fdea173323cc02999a1ffaf2a2511cd4e900146b3b836b22a0cd6dc79255b87e5dde2861f129913bf59213a298d2fcf812bc9eaaa5df2de80bc3ab44796dd5d272a5f772e701084440e042574833637870845c2b02d52b5a710;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192eaf0c4a7c523f50e2decbbe51df96775d4895f58c7c65399ce35a6fdfe6add7a072c2a8fcdbe28d51be384f2f092f85079bd4bfe592b9b6269882decd44379ef1957ce9e3a86f04cd61aa727a2254e7b1bc87168c80ed12ec197;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1caaaa3b56e562c8f4d69593431b77209c076fe195eece6daf20b7a3bf4c47d71415ed8d98871f410fb628078c2d71f75981bd410a5ac6e94282c9a034fde5cc8465fe747be2ef7bea69f0ae3fd784fd1f2e69fbb66a06e734e5f32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41678e662b65045459c3018d25ce5743e35a8e61bcd92abd1ca0c28f9ad7ce18e7d03ac573ff49fa03e54752babba46afc5d8f613e67b4a47e8552214bea5208f584465a72bd0bc768c8dd9f3b84c96b42c19b5591073388e5c2c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa18b850295253a39ac52d75b76bf682171f8fb7e2c5faabdd60c79ea159cb36ceb5555bf02c86b9d923361b48a8efbc07172a28e9aa92325b30ad8b754a81087f37966e8396b94063c244965bfb23abcd2966959f576417108ff7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19851b25459ee8c80eaa742be8b8dd780e38882cc4d7de260149ef5e91b1d7e60dd265830a3657d5a690efabe205befc0bc93326b79e4be1fec376acfb85bed64ba126ad7fcf2a32403efff931792c5c1eb781fdce83841eddc4cea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132079fb693d1bdadf05b60ca8445205ad25b704d0bb8b8f0f75bc4fcafde09f8d20b60f36c52b7f8de28bcb78255ce9259b3e81b1ec2180d040ec6fb1964ca9aef887797e4d223ae5966e457e5ea59ddb183541c7dabc30c8d530;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf8aec8cfdb2ad000d27afd03e6655613b011745cfcc80dcea8e1ded07e7220d974223a51b6a2d6c7d8cb1cd43e246b7cd0e5fc17e63575fa45c19c79d2ea8a29dcb60d529da7b0ae43b80911b04e6023eb696abb9054e319054f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19332e6464fb52319ecac6e7b584fd67682f15a3f918691dcc8e7012d5abdd46995f7633007dd4e0fc658f81bb47f65f67d7bee0084d97f12daa11ed9808bab7e387268620a13d004e1157d19803ca2ee911020296162188f647276;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173d32d8e1f93359071c30071c75c62a147f51c316bb5905224359ab77f0037b21bb0aeb395f89e8b41f8d26f229062c7132d05dea2d279af32c7fedd74cc3aa8b15bcdff9b633ee263d2d4590912bf6a0c7c85edd4ea70a75713b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h980624dc54f3de36b38b097867ebe9ec7bf6e29654eaaabbb3582198289194326e59f5dd9e90279103a2e0b487659b43f2e8fce1ed840815c211e688e9e0588948f9d2e68a07d1f10fad67ed3e4fc03185d36c3796c77412d741e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0663791abacc60b8c9276fe8b0338ba780a36b4cf287674cf437c0b47f5425e7598355c322bd878bd0411a7494d394aff51673e005d713fc68e9d28013ee3f01b5da597e0e1f3b3a73a97cb7765d115b4dace1904adb8abe06864;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97af8c5bb363bc1efd8f68bec32d405b63bda6f37450a2b01995f0b355b45c08f2d2c045b3d45d01c6b607c860b8eb85a0822d5ce4f1c94d2210019b9467f9bf76474e44ed3f99c0afb5e19e6fa83a26245a3d97b822c3c20f1934;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcec684e867951da45d55149d546cfd5ed60c27f67739cef33ce885e52b40154f97b81e06ac04d4f38bbac65e3972595c51944458b658280c0bde128fa4683e95c85979a464258a2df7e25deb514f576581fe2b908aa917b16bb219;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h933a4e0ce7e9f6d80a4aa2356136a91b33aabe680e7e1778a54d20a8b356ed2f585df4f1c8ea4fd095f26eadc5d0b7605b995ec03d2c66971a6b4921677c07e3355953deb64bde77e94370818bba47164ca631722d3fa8a861c887;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7c5f4e81fd19778cf7f2ac922cdd21c78d778d7bce5e7523709958f062480cf787edd07a3580114cfab56782a93408b4ae069fbbaa3df7f391264e1ffdf4e55124e4055d4030f352144a9e93c9f940c7f348239837827887e404d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h778f676bf3dca48b5ad42a4ffb76c8961ab9d4c285bc5e31299da93a328046887c66be61943821c2f0a389d1d42dfe15b2a2bf7c89e6bc5dcb8307c4ce412213396112073a510a2786632d64a7c2ab8b16a4ba9ac9f21a903ab5c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efbe473fecb1f4f0616543f430c495284974f301d416d915ef71cf1e4d596d41c441915fa6b93aca077f8fbe4f9f1ea6bcee278177487a9adcf03f313c7a8aa77ec53df710a50a865f470dd03ca5145c0a8588547967bf919daa6d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177d0ebe19c5dd3a1f485693ae07137a9e4f9901dd6a4632434793dd635e3079027e4528288c9fae4ceb7c1b6d775e6b48f7e163fb96b5ee5139f1534d42ece44e5f02af08077330378f8363952aea190ff903a35d0a93d0f90c1da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ed9d0b21054d0a42457c9ef6c28bd1f2ef834aba98134d1d166f4d767150ba854805f5775d1c1df09720e8650f64e60fe846f8b05cde60f822ed4caa4b73047e602e4399f7a8d2bd7482c8c3283bb79ac7516582c25e6bcc5083a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb0247ce2ad0a13e135ac42a27a1cff69f953446b6b783bcf85641fa441a0d0c9d7a6713101223f0b8b9d896cdb2a3d98b559c78f08cf3743706d96d3ef78ed1b396e21bf0a81fa5fc2d7f8b694c21afd1460703718f872235abe0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102d74433d88a438d0d98550402674114a400d89856fa13c09d1b956eba435c4b931a5eff9c477e69acd921201b6ea43b46229359566f4f969166e73d136b2270e13eb0724a43bab13818b7142227529d3d63c79fb32646b76ccfc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133d5e1ad39265339e9f25791c4aa748a2ea76565419c2553b7527860d70bdd30e6f33b30edf699154af3aa948fb6e476d8399ec6320c69311d90f30588f24f6db43b58fe0525c0056e4b626e418a6a7a24624c732e54ee413fd7af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1495e3cc71ba822959b1fb465de2461d4fd6b2a9a00a92acf223b7279936cb911bbb095ed2c37bd6d9abd4e3f7ce2f2985ad13d0492b24dcc5823b873064091c58cfcd1b07e978e4408cdc2cf9820d46fff8a7fbe3c13bbf93fabbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h674a28da3de2f113d3ab40fddb712d564719c86d8bdce06cdc683a6fb58035a8dbdffbbb20841b97290639ba4312f27f025179f5bdc829d7255173954861e1b94969f6b5cd28396751dd3adcabe757412b2c4dcfd252e818700aa0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171e11ffa8e51bee35c7d230e02c69cf78e7675fd827bec8e2962d315130352b37c6edf11333075739b4e6403b99df35fd7c8934e2ff5f26619e97263fc2e16e92afa1225a202462521d2999682454ef33e2833c4c09fbdaee24d3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he35e65ad0876794f9b9e2a5f5f9d07f424119842c95c179876ac4279b40fd25aa3278a2064c534132554c07eb7dff620720a5f7ca7e46e36e3b639ebd6ff153743d5aa2c2e16d6f7e8faadac0322a037cb2919e980d3b097a53b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha3bcefd695c74d5533e8f841d22cac609fa8bed3f57417140bf24c772abb4690194219f22157be49b81abe7a16dea5ee9368bbf18d2c1d2cdede0b93d88ac5c345f7fda8e95abefe0a9dba70f7ec363a14b1dbb2fa826efd17da24;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha31928a9e1ab34606105d54e97a659006aac7ce74909fbce30e8f726ccd7cc0cd815b17ac1019c78a1f86bcb98829c017b5e516a9589d395c2863e224b4622662a4343daa8258ecf2851743dee90d19b7230cf2762d341360f712f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4c054011f7c749db9310f508afe8ea65895550d76a4719153351a4c9f301491e486a3c9f0a01a4604c178833a320e8fde595d385f78c6a706f8219232418bd881a5d45f5eea1ff89b2e1636d7a9f7fa76396fd10f0d2216d5f82f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27fd814a5ccee6b77340f5b003aec17a994d733ea7124492ca68828770b39c15b3f1354aa22dc3687c2bec3255be641846b9386ede1bcd5144cffd7a8bdad4fb138b3071c63bcd579b3617f8a63eb9647a6934c809db1a064194c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h198be7179fc19c61ab99ecdde520de529df2b3a0ba4607b6d6ac136ca2f0ac26f0fd3157ef87282906664dbdf540edbcb123650bdb4c9c35b5a2252eea2a7da44bc3047f2f0e327013643539a736b7fff5c917b6aa6c141af027a36;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115b44cbace522140adc65618b3ad1e7bd7eb86f5f68ff511c2ab79b548a3d63744ac52ef3735ee2646708a2a0d360a5d290bff555ac32354546b1b2f6626cfcd9f25d3fdd2b30f1de32a8106b6d2eff96430d4d97c9daa1c733d44;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbaa147931924ba0a30b872817f408ec87c9a16bc60e3fd9adf977e0ccde0626a5bc7e175e22a6f4d067a764b847bb2760f93a41df6bc96085009fe989e53ca7f4876628a5300f69c73464d17d186bba15395e18f71fdc9e1add45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h364bcb495915567b6e9abd4aff5d1462f9b4d67336578780dec77105adcd7f65d850f16909e8331223d46b395468b473a49d800ca2c470b2ea08932e833767a810a607b97c505fbc110cbffb1510bdd17463ab3fc8412118d4e37d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4afc2e425a90bae8aa260d67e539b1a7dff845fee2a58a57ae26b78e46aa09347eca07b2ce6f9728576378cd1218f5ef94df500a01dfba10ec80f534e213c6fcefc1a53f0826adec56f9e0d22e9d38022d06c536d8ea784cf1f665;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d9eb484b1a3019a0b2204afa7b6c6290461894775ffa2a959fdb8b68fd1932ee0a37fe3231700e5c4683ac2bea00150937d2b2d6bd2fc3db857b27d960422ad373dd3c946832d26814ab2a2664e9959f84bc69d380da67f131c34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc25910684b247d0132bac4049ad568fe4142a7c8e162ce3c8a5059c64da7f53644e391b229284db65015233c60b4ae66a107b8ab0f85a58324686cd3a4b102904b9e862263aa28b0d3e315e3fc784d48857911815525783f3e3c62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ae018c43bc6a63fdc7e51dc958f51e18eaaa2c777b44251935143f511be87d97c43981f9b9d0c65587b8395330bd7b27275f8efd504186b37946d82f3e1012ce0d3e6751de4f4268330086395ed1aa1721d5025f92452bc8bc9707;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h730fd80b381ada1cc65354fd04b9dc6af16160aa3c809518e0a9f34b91befbf14166a05f30cb5b29b68f5c2868c5d3c5555ec9ca55eb6b37033473b13b636ba05d272407fcd4a37fb943c97f37500c58a1b5564c9dfcf9c4a6d631;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8d153d80d3ff9acf1773f2a6a4eb34343e23e834e5c51ea42675e5c892295c91f7952159881dd1f7ebd545d09fb5c4cafd2c9417a30d35afd13b4ed9dae284756f4e59465f15aaf789db63b283e6130993b0136cc018c1006280c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f8e4f367155c3aec567f22344d23031e7a90d1b7c863bd428d0e99ef9409bd0c54b0e087343d1ab9550be4ea2a27d9f7bb0ff6ac8b3b74612a3c47d3cd1bb45725d971db6246ca767bfe4c53562fad782224f25157332f87d0618;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'habb5794b2500f82e57ea261ea6257494e9c10ed0f17d5a101d0826f0af5f0ea63a0db4ee3287f141539a9dfe4e55f63b7f29c2e8bdce3ee7cca827429afa8d1aa69d44da45c5de9515e6a2722fba605f5ff05b02a67cdb1200ea7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1553ed11b9006f71457e52bebc36b72ef8feeed2b849ac78bb9edc5091b75f4e0f90d90ac6cd010e417761999647033aef226c9cc84afafef96800fda35f66c931be184c9912ba1009d65c5a41d66a06d8a3f799e5cfaecb60e9ede;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59980a958f1ee728feed6f4f31d57fce317e0ac34d87599ffc783359abee2396b8b7894af82c95d3c3d2c4c7499019879a225fbc01867642380a8a242cd3d92acb08d4219bce1a6ff5428244cbaf6ea71cca48a9e416373990ac5b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a93c034e201ad2bd88d2b0ae96cfe6f4b459085ff8887d0082bda65ca376d04cd48cb9e59a6207174c607016627ff3a5b6bf1d3542e2562c8ea301c6ae3c8c1b225d317b158705abda9a6449f94d45c70852ef13de4481a5205e46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c16f0c8140cfbd3df2f45f3ef47d5894772c5dac860b768b2c6419961ed3b98beeea439840c62da1d282100f8d5bada8f099476374f6ee2bbe3aab3790447a0319b66a601b2876844e41028a8620b940d355634875123758d2e76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122f08d3d61d6ce91b75dc05da6e22ee3636300dca0cfa46bc248105c9520ee80cc035b56eb6076a3ff8defa664fb731756c21c695474fee885b2d6208ff6853cfacc5ca54051c4122f8d114962e1202014a4b965ab392b1b6daca5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbc8cfdc7871aaaf75be428fb316fcfe7f48da118d8f727832ced8e35d6ccb7b92199d80bbf23e1d60e317ac95c38bf1f24ae573444a4de1bea86ecb646397267a5bab37577454c80a205d82d68ad48684082d6cbc1968f792047d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16727ee83538fb7807699271cae3bd00bc3808a424685e0f0a1de4d62f1de0014f56ca939988d4153ed3488ce7ca9f80ef1d4e08b53052ade0cb270bd086b81f6c6f3147df86cce863cca37bbeed9e875aa4402d0c6cc956a52649b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e0cfd29ea031557aea2a746d04a64c77a742a67aa11bd6a8a0c24f2dde549d6c7b28d213a3919a674377f8135c895a7bd01693d5d8d42094577bc9e69dc9de06b7e6f81c8450009f19dfcf70f645dba4931be40c79cae21c24182;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ee8e4df6c22ce4a60a4ff6a7da842029af359077c5cd7cc423c9b72056044448b02e0b35a7ff659c9c88304c7596debbd10a44eac6c4df83d2fb5013fbba6ba8bee662e3f4326643088c5821f1353079851f1cfc2777ff224880a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58a6a148a6875c96f023230b893afde60e8ef68f093513b8fdc3653b09dc7a8f2fe08f56306a8608144c7141615bf075daedef5e3749d6b4272aa922a69af11dad129e00a30bfe51620d418ab187519e5d76f6b322731fa9ead77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha10ac7f58295d3cc0815323059ebee1657088cb1082e570dfaa88fff6e4eec562f90a2fb095719d575c3e2ed99b2f1e566aa5ea37f2d2a075b90c4ed3309c57c42e5a3b342f69f66150a2918ea15425497b62831921ff86fab79a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10bcaf7a5c53738bbc003742868ceb3c4598fe487302aefeed5788e532a7fc2ab2a8c3e2d640a4ec313beaca870432c5d5082d9c0a9b9341661f082a9d31679d6a731a3bad29c1c88013b4f8795ba18bd016dc5bb84d7c5db266e66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6ac082848c0839e0a73d77f2676da6f69b39c6bc9500785bf59a55b9b2a5ec9b65c8d1e87d26085e3e043f00f11a1a768afadfafbd01fd29b90d11da53ad267c4b9dcb3ba8bf43435c5f1f1c770bb25174d79ac557d4c9713ce91;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6a3ff2cfaec2592d3103d0459fd18dcb7b46c0587613656d08eae1af20dd521df5da5e6ee09fb83d5b433434453a27a1ccd95065c715bf1b53f6422e7fade835e34bfcbb9579656ebc9a796c59d52445843226d3511170f03861d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c686e19e5ba9e20533b265982ab21fe91bd21139e4b6384a2274dd216b347bfe8c650312efc7c073d748b9570cb1c7fc8e44292c4e2a5d71705e82a4ad9e33085bf845cfddee43a03fa8201392a860548675b0c497be78fbc815f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22d23c3b05e6000e2968c26fcbd5c4e188476f96201ddcbb72e9adf106f2d7d49b21ffc964468e2111e8ba17d9b75df33d7cf92f1bd503421206a66f6365afc4e462f3d7e88594921ad5e00e712789a8b86ea92667cbe418ca8da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104c9f1897aa8d754d57b3032b709fa1ca46ecaaf0f6f374313b86a50fba157c2dc8505bcf7318981983a74a7dd563799ba18184dfda105271f739477c898c45b0b06fee82957978373ee50edd1516bace0d45a7162cd5c82b24e99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha0b7c6d5ebbd91e0769928cc92599f9fcbb55a802d78270e032ed7f8b9593fc921c0241b6626c23980578ffe934ea90844b7fa9d57fe4feb4b224d17ba6f77685e6aa416d256c743e3982d612f098bb73964ea71d409a832504cbe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb874b868dbf47a1d5397da9af5503ea08fa293efa4705552875f96f7de0a0884bbc31f5001d6266f1c17634c5ab40f66730ee70f8d00ac38bc03446f41a46ab6a39317536acb5acdc9caefa75c8bfbf9f8206cb695294b17e67b4c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1855aa073409303a316988855789db2d00e2097dfbb24b321b9f5562f2f6792ba5a133d23b848ef578a5f9ed8ad9100634f359fe7c4b7351f8425ed7ae9d6b7b3edc4d5d86f9d6789601e73d330dde8ddaccb74ff2c6c1396c27aaf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h722705a72ac5f2bddfd8c71d06bb6f91742cc0d2f17310876c8db9c04311929b88ebbaaafb01ea988f1104177c923d702ee62b551c6f33aee43819f4525e7c8f0b4fc0f5cc87ab0f1283c4e36d69e25d97199047f06ad8b218fb7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80a71c974ea18bc35cd18c239e0a628bb1ef6015731132129d2dd89906fb7b1efdb0730cef12bba67f391343e1e3390a0a2d22881a68e98e8e584835804a4b00edaae52f32483c98d67b81d784d313ce7b0482dc2a1e9db87dbe17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9cb23a5904e9cdc1c1b0d0a0bbb88a63d4e9aef4baa6b5c349fce6df2694b4e5dd039a0155292f3ebc3b80fe45d9e2055bf9b8600238551ad3ed6cf7912c766fec5fbecd219a96c71f0945eaaaf9494d97d7c1e94b608d36def6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e2307da54a923bbe89c7abb0a7cd487b50843bcad403a332f279a65b38bd8c85b46697e35e574219d352006beb36b41589f396d2a4e0b6b032171ecd95a5814631a54ae3d9c98265c98487887f2ecaf409acc450a0007377582a1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147c05559b59d7f11cc4d430a23083b70909d77720ce8edb9aa3b4cfca698e50e55786f731765d0b9fb612c09acfaf4d4b84c75d0b9f4c51b64064d2591352120f3e4b9a42db161abdf25e1fbbdf7dbb29edff2403b1be61adfa9a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19725630da787ca8b64918c7571dc73e1fcccb12430e0d2958a820c84fb6d5130e725580f43b19d48bd10f44bbac6b52a76e20b06272c50d762bba26452ba1aad9c5a6594edccdadfb29dcc4ccfb4b2944d5690a75486425ed0cc0f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72d51545e8ad33ee27b6d9860b80e582f6fb8976a6537a22e4ac4779752fc883d03e50eb109a5fa5f57947158625618a04cd740e82318452a6c7b4f6ecf5c2625ed307536062ec56b6ea5717a8a1670c83e7650f6e6b2dc46cd78d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f79045aa0db7e471f9e5b072b96b7d10b9a39d26e402e6d7e95d69bd0d58f838f7520d0da9f8df10986227be17cc98f2ef2db285527405628556708b9c96b768abef2e42b068eb8a6a25b50692432622d58fa5088891d1f80a9ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1665a5c794986fd1077e17d618618548afbd5c17d755e78c7c1455c400ff64f0643433579322b66bc17c65e4cc3b89dc0e51ee04860576634a1fa72a24d287ae903bd134f3e7c1bbbb6d94d813281d05e242e8b91eac89803e682d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122ec8a2f458664cc6751da674493f7ea9d8b04773112e247b72fdb922650acaf78f50fae52b6a103587910f4abb2de200d8283d1f8fc8ef6b57a08142b597eb30472e6f34ea728247c146fd0469f60d8cc4dc9ecaeed2edd0555ed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d91262be382003156e8449e67824906c4a8ee43002de3549a6c93513a2adfc9289b6b1098bd43a44a2c7288e26286280fd7a58264c6827565cd1433e2e54a9d711c36d2ebcee62de78a8c4d8b9862b5c31cf20814a29f4cdb27750;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7f86079018c8c17c6d23648fecfbca3dff33e5934e039e954bc02a2a07c92f8f9cf73a8cc5b12513a51b27db38008f3b30f54d3adc8798735aca305a091e37e28fb7a16afa7d30164a783c10e3e263527b962da82d69da100cdbd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbeadd944a860c117f54af3b1f231ddde73d376a4b7a4e6318c52c03592e5b27d5a7d0d8cea512e6b4ff332bf866c53aab7ddad922206674d6fd9ab3202252229c3891031a6e8836d4dc3592e084ee1cb573d021ba27ff1a85812d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aab3857a0ddf7b8bf94f4352b0d5ac32c3546a282344a6145873d2b724c3471d3479336e7b4fc533510cb108f74ce25dedcb91660d9ec80e845dded8630f8f4aea9f0e330f57ee703f90c492edfa5f16731c7c0be2d85f256d008;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b7e8ac8b34f0f1c8779018ddb228c5929ca6a79af5e3daf3d13c48f0e13a1495f1fac41c898487bf64f2bf30db6badee4020690be2564fd993f93e53a8ad6d11e26d8ee07b0923b0cafe9527e7979e7c2a7edc5667cd9d8db0fde;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e02017bd1170c9ca9ef3866f171b004f72e2524049eb7f9b9ffab1664aebb6c656f2849a1ace90a3ffaf1378368e66320f9f51aa8cd99e7fd9d90809d7bb4e113e589f5c23cf9002cda63989038eb71414348d0e62929301722f6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155bc5864cfa5516b237f8b61546e23055c659d498587f68c2b03ca0d5a5a35e0b79e456ec0596f2a9901531d193069747030551447e2cb8b159897a5a72b58d5a36b0b66acc4bef60c6a305e61cdfd41c796c749c30da4e3fa3cda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ef2925b4b52cc505b715038569e28df9dbfbeaa088c8dc60b4634bf6eb5a451ffbc02a42086bfb576e82c16af305ee74c66b1723e5d064346ee712606d700081481beaba1079a9e24af6b50cce414b9dd6768b011f7fa21150c34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa86c12324466d93671f211a2206b5e45d474d5c34838fa448305709b0a0f9d70ad50fc0ce185c6a995649697e3c6c5f70d144aa1ee38a19396445929313b94a7883eb52ad204da2b8a7a22373f9146ef44ca1c5f7becf59f71f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6af2340fb3cc2329e3ac3f4fd3967b8bd208b5cceb3096fbdc0dc1197a1b16b207b4f4437c49b60204cba2d8a3d440e4b0c9fbc4486ee1e054aa58ed29b92c50de741133b3a53e6feaf25e6ee75a60c9829f15f4869fb02314f21;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b881cb08c3ac1320b775d885f389916355037fab7b5323b6137a49f623e303c7361dcdb31613e1729736cc87ce6eb6945a9fa52a0560a57a0fd824c632c7a3060777c8ca1a31f8016b576ecd375efc115c9c0e0145bc54d730491;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1212b3e0645e1b6b99e25d4aa0fc9d15928a7bc582e14d87431e300c4442e802c5c64c454a85c836d004b453094f4aff089a69e2320814631f7d380063033aa5d112375a679ae658a02b30aa2941110d082b9867174264b568832c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51171624984bcb2f29aa30c08ba35ee5e37e31af9291f3f43dc0dd2bbd0e5c06e362316835314b2693e33824c93441065cd83a8753d8fb5165c20c2cbc231067f7eaa0b82b1f3c1e0e72c368d1f94991b1fe52f7e8f0335c955c2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he98cf84d6cdc568ce8ebe9b74f78fad2cf198e514a327554213ae4b90a3dce53b239263ce6fa4e069b34f01b3980dca9a6fccccb91b45e6bb00f96f4b1cb889397f15fb6f1a2c3f6a17d422cfe445568ab13917ae2cfd790c15a1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac34a91cc7210a015aabe4dace0df0789bcb76f8aba76d2b0bf0a6102ad47f117752b4772fcfab0c3357cdd3af8a62db009e96dd3d207083a5d872832d9f0096dc490a53c17a108279d8f1fc85573c6b5b3faac76cc9a51b7ec39e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1222e5171af5728d51566324e7d38a563006768204b7ccd60954e7a0efac4d3e0e21c70a3a42ce5a12feea98a101cae66e6a0c560de0dab16207ad8676d4c80625c61bdecf8a1eefc905deaa1677a315478d5a8ffb68d53d5d17fb0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdf68b80edfb8b0bb4205b38bbe01d1df81d7810860ddf6fccc0f873b8eff79ffeb9ab36d50059ebbcd6f0ce83e0e27cfea6ec6508008cfcae6a73530441d94a02c067f4be3a4a17461f9c948726fad58bd67c95347e45aca7c191;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8efa0fc11575bfc09d02b42fb71aba4c3c8df8fe34e70f7c06d11bca2a6d7682c86da5a5d9cc7654e62ff8046cc4c98470d990711518619009a3a47310f25c4a7445640611b907e1c44aea35ed5280b87d78532fd0d94356d9460;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2c38a6e0288b8db3251c92cd0e9835778140cc380379872f97df05a10864169076744276bbd9a62814bc6f0d63ba4465720c10c06f48018408262d8eb18c36fd95f1f625db3656aa8783abb8e9adc821f982e7879dae608d4f6b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4254d94e0c180fcbb8f54a99c62417efef6181d08d32c7281c1cc105f28bb40867ff95271551ab52015f1aaa7191e1d10c496a3a533611955e5e10592d2285174750097ccf2efdbf1cdf2c61bdcc8ba3ec473532ff0b75972f0726;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h938a85b236453d36933781fda5aa1a0153cd91c18bb1f520311a23a4ac973d1fc4c6e0f0181d3f637911e397486bd0f0f774cc850cf1d99aa64152c816843dd7d7beae8a5d94548a8073c6d2c61a5ba0d4953ffd4af61e4e26a24b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa5900dca21dec6a773156b8993827213e541d17df86f66d31a8747a765e637d4c8d0d5050a3a5d9a38108750ff264259f87c325644da40d74bf5152b9d75d91d70c67a69b57403ca2f3f415aa18229bf31ae926504d0b6831ffd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16778fb80557113bd5a35db1eca00b3a78776614620946fa0dd04fcc973d8cf6bc332b29bf2d11d7f02f3cbdad4317cd38646b5b780ad7c8f8381f16c0984e63849c3cee82e8a58648aaf481cb1e2b802401557cf74da4abb786f34;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b43f6836f1364f9f3279dad08340bf1d9a6d795a75cdb22883d61fc3346e563c6a023ba7c83c99cce26e66fe18460440796188b521e6fce3698b66fef1e82ddb4e855202a1b52fd7a720435a340065967b46b2154e11b77a7b746;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h45274c2e1049ca3908392b4ef1f38a544bb95990311bd8f7e7e32faaaa7d9e4fa2a4004007939376728fc23a43361d86490b7a45c75136960b56102bccae382535bae11daacee31f2576be88bc393d1001d6538ca07e381ee39d74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168b4df21bc13ca54e7cfe605088422ba04d976332750dd46634fac2646efb27d31ae34b77dbb2dfc077da46649db942daa0deec309ad842c6b694a8560b0a69a0dcef634a254af2c855719ff77191c6ad98eecd3eaad4d4dbb05b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h636d1aeabd25ac200391c8ce7a87a19ce5a97098bbbf5243667a92d74fadb184caeb075e799be2ad4b65236a5b084f273a3e0d0f8060b0da410be8bab1211ac37e89fa54e09d87a4516985478d45b01f58437881dafa5afc95d5a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1093708dc731c86dfc8b3caa9aa38399c7e98ef6af1bdbe87e9409e5a114e7f67a05324ad25c00b5c399f8fa1c03aa685668085f7c4d6e1cb4c660eca1e2fe5bd27e269b42ef02f502d96bba8d9f69dac152dc1d4d446a9ebe25b55;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9a80f2a43baf884d6cd1ad2d40c19bb93a2e9311a6be1a4aced84b3897433693ceefbb93d173e89d0554940d50931b8e00467d494a2eaa9d25123993d4fdacb7d9efc98203fa958421ffdf4b8efe3978818d5f1bb20f30535d6bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa2b46e66deb5646b5425c5e7335a51776bd891f831fda05f3c6a8b09c7e95ae927514c525e9424d26ba0610179b84036d2a9770ac6eb0aec267a30c25b8eb6c95a8195bf7750d15e92a5c4f8d6ef7c19ec067ca920b679ece6a72;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bbf5f4b8bfc19cd426b4619fbad7ae32499bf2c3da6a52b78b7f668815a93bb33f76048a22d754f540e434ae5ecf67c6cb9b7291dbbdb8a5ecfde1f2aece4119dd5ed668d1b4c552cbf6d291312e9f370976fe644635e91965ca1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc0212659aa155ba537941527625259f7246dca7a33dea59e6e75966bd7ee0494ef7797b1b6b085a29acf3babe3f44e77ec35e8a5f5b5b5f83d881caa5f8032c2bf78474edf159a7919c263859c688479fe06d342a5dced379b31fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c4d6524bc7b68e91d88ec01b544a437060e098fc198aab175f19096b5ac4e51dd67815bfb4227aa124f6067e143ccf72e3a80700b0e036cdb75d30571363e812afd8c191ccc2d02e0105f362c9e2263d56427ef285c820ddffdd69;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f7ae224432155158ee7fc4381c1f6c13cfeac07c149bef92da37969767485dd6211c5fefac8fd411f6831fa70ccf1915448e3d91cfcbb8bc922127ffb8eaf7bc0b034ef3c4c2df6649349540130756171b06cfeaea5231ce2099a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e119756b6d29b78b1e9c7c65fee5a6419023086e1a3beadc31a8efce5ff5d3d24d6413840738afee56a0d0720d52c593f7f1412d9967105fedf523b22f52abed76532f97491415db04a32888ec2a440d822636ecd3446ec45e438;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14d1142e1ab629923fcf29cfec394af0f168edb051884cb02cead37c8a844e6316b582622da1e179968b2b767819341818d158f9e06eca9c61f9f43005fe25aa02175a401439d07f64977c889281eab91659303796e5745275116bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b4bf1b6466ab54c345e32a32b8793616377eea28944fcc03af2209db9755422444270bad14083eaad584544b23211355337517885c82b8dcc859f42cc22b6fb7c3d70212966201f5dbb85b2f5728994b06438b3a93cceca9a32d97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91e85e6b3ca8959aaa1ba408126018d6649e44f410f128378ab7c91d208bc8e052045f80d5a1ed56dbb3b876f4f33e64c21ca74c155aa66e005d55643b5c7c82f0d0941538f753bde851f65f767476aab9e52225577d2a7104e783;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb71fd451e8e12098704b17f3726f55baa3f78f807f8b1ea14af53d936eaea9a74c0c2a0fff020ecf72533a5ac01b14d0b39b69db2475e9bb784f0a1eb53ae79576738a21ef8457fd5b5570a65d68f53b607a26a22df3a5a580344;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1128d68f8224244be16fe37fc57413f1225648cd6e3dd447701db8442a26761ce347d5bb33089c545657ec793c5d32366ac10067c878014cd6e000f2e8c1c7ba8ddc065ad9d207b9c1ba1e07dfe20ab87b0cddcdefb6ba3ace65d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a2364e23f64801a7a4122cbf8e5c50364b83407f04f6d86e3800fef915c147d2ad167e2f070d60839acff13627f197c477100088554bd1ad96f5246570652512ad9558997093388aa8153017e4dcb9f23a0272bd3b19fe0c260fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h145cbfd7e0191e12a8faaee9d414696f2f1b4b4dfaf9ecfca7ef2d1b4c3b12ba7e0b3ab8f3b2b2029c5793c68faaf53c1d693e96110c0f6a3eb2620a668d2e7f836aa4886ac7ecfa9aabec5842f19957ddb551b4c4ebb7faeaea0f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa165e379576ca4d15c2f68ea8286f1711f10621ea63cbfc3b84252722c0a2d3e2a4967c754749e98e1362ca7fcee76f465eecb2c9167f62ff1bfd8ea69884db380b4a68fac0054770195369b23d46755e8ea7276eaf345ccfd66f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h91ec7c26575cbb35f7fdf23a24b58d72280b16e53464b33028d18ebf1010737c122cf377424291a5a8b38b946ac5fbf330f94e7d4f90a72dc44d059d4ae5a4356870e74f39dd88f485f4de240a8e0ec5b1b0a6f9eeb7917b73d506;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d15de1976006a3bd61f14f3da5da073f68dd3ec54969eaf2a4370c0d296f18a060969c7666774529fa7fd2ac177d0d103c5906216ff0da553feb76e3d1aed547faaff2f98d6104f97969852b97f63ab0498d0d127322d962e4f7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1972b1aa9ab1b2d8c6c40b8a5cc4da689a968f12a4ee1b672e24e5583a2f2eb3ab2fe3f9a659c8099b63bcb6926bce3bae2b57f45c056dfc17316915360e27e54e7ca7fe06c01a092a12a767d73eee4c7ff17cba440c03394ce45c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4e0e41c46c343f77a26dd01aab4227261fb4507271ea923bbe1538d6e36f6cacb3df4424969086405dc9d6b195c541800f693224131b519e0ac8f7eb15b95a6fd0c95080e37ff8efaf2e3231566c7ca26750c10e5d53f821427d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc13b8b617c9b0d66ae7b4b3ee0213f77ed8e796698e37eea46155c2d17c39f7e88f067f4108395ce4e51024d53290778e8862062ad94e86bcc11224dd71ec59d7dc2d45fa4f606cf046b5ff2bb7eb96983021909c1431201b9e11;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef24c05dfb1219bcf50e99f985f118f3b2d9ac14391838793fc6a572aadf4de3d76701eebb3111fc8b044c7a501b7256004e3bd1bd0b930ee817f58ede8b082168e5d84099b3e73df9995444dd150d407594012bf1059f7709718e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf53f23636e496ecea5b26b8fcd0eb4f1d78d9655b95604a7e8a94ec203c0413f06a02ff7079a9299256121c5290adb0f8b7cf519e625ba36a3934c6438082cd004594a87d55465011c313697f44a0eb3b3737daaba33c3d0a47f7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha766e58cc2428a9b37d0fe2a5ce5aa1e3e2c90ae23e77571420ed694e594c4d5863438ea9b555ccaa0e99d208afa64c5a8ead9961c723f8206b1002402ca823d36c8f45fe1403ac6bb9954021493a71f2a6c93d3f6526055051a7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb84fa6b7b53978a4784a1dfb092a303134d3b0a5699256ca06c7005e8f3d57d263b5c629787658068a3bd084a7e5f5df57eced8020e499b9e94fd02975479ca9cdededcce0411083b8c8d14162b670958e5d27389ab38d7953cea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b4db170218c4b292132b4bcd90bc52f33e489ae22b8f672da95201ab5ff6bf589aed33e9ff7a043907b7975da7e1bd74a1e6a61463e9cdde72220f450eb07da9221c034382383b74b28434a22241a03c9dd5aab6fb2f7b727645e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147e88245385c1263bd018c6698921d7c9c4e2d9df022f485b530231d793976544960a02f7e3ad6bfdd2b31549dfbfbfae8e0e5dfd7d4aa0d7d17248abcbae0e8b3bfbef383cb9d3d63f8452803fd4cdf7c1bf57a1a84fae1475c44;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1392df15f98de34d6933f73f08fccfa4a4414f74e66855fa252624ff30cf642f7a9a7b39adc95462176b133f4d2e9b1c40237479072c1b142fafda35e804d950db73d54a5a5f1e58e7b7c42d1e23a3559db375b13b6153962657cb9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b635660fa961934b427e6f96f7adc2eb46ad2dd62047a3ded4a71fad6bbb6dcfff60d0742d4b4d3947cb51a311d0b74c7715bfac8d4813cb3b1dba335442ee7ece0ec8b38e60ff5b5567b47b0681610c06f548218c29aff79e7554;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c94def09eac3d41bc7f626eda7657f29dadb5d2c9c7e5ee9bac5f1d1bc4b208d4cceeddf2cf46b25a63632c2936dad78f674b317189d07965ceb28fa5a50bd8bb4fb11b49d1a5b16724873581f5709225664291bba2f7478386774;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe1800e7ca7bad7ab9f2ea0c0764a278275c9779c580402e7cc41f5228cf296ab99f5fe58f9554be3ec6af3aee14ba8a1ef8fdabb572d0721681c7bc98d293b655a2bcfcd929cb6fa3e68b83094c6c0e63b0c16c1b4adb4e8230bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1795550075eda26980285666d7ce83427edd05723c0a5218a6eb63ca653290f2c3ccc9d581b884f794bde537d3fd874d397fa0a646e08d8138f214a642835c214388e2738dd0f7ae5ad285d8eb4001f89cac17cf5e621132eaaa607;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f16762252a587b19cd91e2d311980f83b058ce4cd6a1648aafa30bde6ff8ca5d1d84cc3e8022eae4c657c6391ed5e72560bb8f84f457265ea191823151787ff1e2ffbb7b1c62c7cff652236eabb8541338cfe1b67312cbce3b89f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h526d13d2f064d1b85e201a894a4115dbc85ee53149063c6285a72f7504025db32c1372d8ba7d8e885f5eb7674b7654849664abafe880c9d6878b35e3931cd3c4a0344d8bd11e57e2c309dddd9076b6908f8916428ee5b66d677e41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c2d6e3d1b2607637915c3d39191a189b9aa78897b22db01517ac6ac972bc3dc4136a2a1ee6bb593e3640f901b33e2e46aa2adace33828850c89e3d193d50477e0f52db91902ca47ad7b55fedf7903c032db4684a65652a25ca6c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53d3ef8536aec89b95655bfcea04360e337c99cc4d4c03ea785aac4b5b5aa1468b711f4dd18457012bc44bc7124c9cfe04c6da3cd9717ae1a6539b955d0689020e4376d475c9e09d5fb0c200002e9d483f996e09b3ed36619f34e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h516ac843aeb1708341e895c8f1aff034fcef0527d6a763b502bcdf5258231d7515216562507ae5dfd0f014bb932fce07943d76cc6870498a4801b3175d237f3f0e7419f157abe4b9de333461a156f34925105a90a06f052f544cde;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e79655c6e7b40f36d30cf5ffdf56e357a18bfc4d4ca14a91b3548532b5ab2d7213c7d240192252feca7436dc360174f915349fae74e909da6527651023753da30215a142ed3ecdfc026ab4f390ea407dd17f8cd1635dba1b7840b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1476b862078ed0cfde589ca5f487887a6b0d26453a8e9afd8c90dcf71896faf5449fc4eb62baf114ef1b7aeda94b649c898ba801a2fa0af069c6cde2dbcd3af6ad08fd50ceb344de71e754b2e501eef4b139e4c6d0e1924c1413eef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6df8edb7889a5e28f98c76e67ba466178ada5d8640cdf777f9f3c7b04d23263a36b1595ad517f40fbc918d825fbfe8702c9699bf0a10ea16a3828af9bce1b1767d957fadb3d03a369385ded7aa94fd3eefeac96db298bcf532d945;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h718b5089864bbdf968a0640927865f5ce95841b71c4f01a2b557b5dd192e442f71f61a27c339f2d3b99cb42bc2a633edef320ca9272a5c8be6f14b1a541b6133c466d2c59b660abb83ab9107d4a1db0ff6f14c489fa1b7ae2cda8e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9dae747d0e5b819f7d51eb3cde8835172878355b4184fa805d721b860183ed04bb4375a22a80f316d28f169d0cb765e49272d0ab04651b77df2b217851d9fc54e1e93bcfc58f11efb4506e9321b554546ce764a81da8a6d40d9307;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbfba6ab7a6c237f8377041ee97985ab048cf6239b21e25eede26665470e9e41d7ed01efc7ccc431281a1f2595c901587fbbc755db100eebff4ff8e275177d01c21073eacc567026adc5e7f88b3993591ee47639433f6ce31a8153;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b39939d5acecb2412ac06d6e84cfd2c88e0f0b9f6704a4d53d09f08a4bf505cb1462e772575f346fd9d4f7243a042575d16a276ed8ed046828570d90e3d3c3b7547fe06b26e42ae08adc2e82e51ba80922dee74909847425ce45f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57826783a9bbba5e17078b593131b3c5614a28a89ba7be16671d2219b66285a496267a208883b839b414509c4ed66b8372603bfee203d602db8a977df5e42850b6a24d29befb0762170b0bf8ec1016045723716f430966e6e808d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f38688c1db9ba3f8ad24427f912b460d352a5d9480f987ce9ecd9445813a6ba117cc00476dfbeeb73ed3a116b887e8318cb2de29edbe622bab2634f137a4329329654490a33c268fa51200c3b0b16f4633d61036e3f24c935cd46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188ab700e25441e9c3e8a582f4dd6010bcdc28012049abbe9d90c41a3e0a49d95dcc3619e1414f7e29349e9dd20aba45193fc7be44b3fcbd7cc77344cd70d972281c54aa9e74161f6eb1a0cd376a0d5391606f994eb8ead66efb399;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8e1533f5aa31b2601bd36b8832f3b4ff411fecd6c40ce1b90be4468f6da9408031d96bd9f64f4025a499d0f3d7e0a4e7a3eb1a19bfb87593762ba6bec18582194c669942c0f166aba1931af2173021dac31e4abb73821061e94b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e266ee14107600f4ced386fad5f5e1c66eb6b245c35481e5564529051404bb958fb8992415930d12ffe509d562095cee5c4219f847133cd4789b02a33b26aad4673486bbb81a54bdc4d797a3480882c928d3cd620cc87206104228;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4213ab123b1697224e3468c1867d70578d44642fa3fdc1dde91faecd827a08cc856c4169fe04fd821ac6653df64be48831e76a6e97e43db35220eeb21dca94e5100bf9475fa23a124407460c19d1c42f826d50db5938c3640a4580;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff7a3aa1ef655a8626e3da509c4d038e3539f6729bc0000d10e80a9d5d7d10e57eb1dac9f8e4f62eae23a6511ebccb6c532ee7b331427dab0475eee1527ff2d0472d7d3b1b4e2ba536c94f2c09498c42eafee0f02f0e8867ff7754;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf94491bd83c2c6f88ca22cbdb4970d00a1afdfc9b7dbfe8f0bc5ac43bf0993fae42967e62786bba2bd85b0c6c571e6affba9ecc520f1e3e030d8680c04d4bb9c901a5f3f2063481a2d3b2673f7984e91d75c6d0dd353432f8e758;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8382146eda048ba2915706c59382975dcd689dacb8a25e07e38e913c563a1157d2511f7e63c929792f67683859224e774f16be35666e7d7b3e10c6fb03740744d0c6b561792afc1ce5a092855180521ee8ac0e014006950144cbcb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1faa223f3a024da067b8e5b44fa0d963475d2ba554a1406017dc27672b0a5b05cf62ba3e7d6a950094bbd00c12280e1b50eb4941d7f800bb4c4f14b3d3df5beb7c49cb5c2116bb127308f98f1947b7fbec423012030ee9938c1d04c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fa5125387d34720e36e21c801b30c9145a2fbca2db31cf763d7c837ad3cd517e3171f7af5f8229505b836682f192946d8e9f48ae3027a9ab04141a2bddb69e2a2181425203406f7e8858a2c85feb85c20607ffeee6908617b7909;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144353b6c17ee4be623ef3d50c837f10a0292aaea400dd29ed9b46ae6d978eb38ac2c03020ca4fb89d08f7cadd2ff6807a18cabb9141baf1d221f7820c19d2fabc27711f2cde84fd52e2cd37c591b72aa1a231747d778733a3d6487;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f00f8d408fba8a10f56bffcb8ad0f84553dbe0ce8e958ffedceb8ef0b1204d6f74650b293d9cebdd4dc7d14a85f017306d5e0d7c74a6fd421b80a80f4048b75f2a1d6d1e990de94d69e925f9ffcede8108b58577f1937c202cd5b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1754add397213945f3a111a1f0d345ced3af6f272c201dead080009ee2700bfed5ec7af591c0cfcb88a989f8ec4ac8367b8f77f0eec76157cedf487ce3426caca54612a70f6a80d0e6f19466113a5f300b0d5b97b17012d5e33648c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ad5e299fd39617c580c4c6c92a926d780d223ebdb7ea64143f62fec6a3e0757bb3f2904b3c43ca45325795e5587ae06b7bfb6056b0f1279eab3453d3d128f134987b15131881df45c3bfd9e16d57c855dffa7aa73c4b88e231aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f4beb785a000562ff9fdc29013360f74a28c877e5b1dad3cf2ffecd4493ae307c0a958b01370793727b0917438bd65ce1799983f7991ccab4873ff6b3608e86bb62e0c12b2e7c2c87788c09e94bca2afb212d2c5b5368122f9ced;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2c806f8a5f646bfab4b304ac5ce9968c6ba649245ca6acd07f69595d939594eed4f7d06f1d10271ef88c24222fe280c6ee6e1b8195f0a1f2f545bcd795cc345d82263a64f6b5387628595afa264a6980fe498f0df254c84e00923;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63410a7358abc7ccbba813ee013d4a73dd35824b1bff1af5f7d7dd3848d5324b82fc491d50bcc42479673a96e229812bfc98875fdac2228d8b60ffe05de75118a06ee10564b542dcea8daab54af8794f2e1673ec08891c58e4869e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2b63369f288345f652f9f52026b6dd8ad0c862f991c7eb94a9d9330a6ba8d809d988208c4a2596ce109a85432226801ede72aa21f0b2f6fa17555d7e1a323a573742cc517cef880a67971b4e5200e2ffed5570c8978d6a2e2399c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a2ef9b2621102d8da2ae436c55c8e7ccbb2e031012088a20e115ae7e2d50cbf60fc2cd2c4e193c4af1649ebbe0f8f5d24058570b81e687c48760fdfd221eabc8606a7d34d9aa876291247b318fff366f40ab9e38eab0469f039d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca4905623b52ecc07c08aaa30196af5193541bccac5c516044b1c6e98d12a4eb45710dff562fdeafd8bdc1102924814f06ebc0ab842c17b7f9407e656eca50cb23d14f3c7286ebd6f67773a7643dd781f4b54ef9692674b020ff31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194dbcf195165ae72a5a9fa78144544b4aa71acb2bd322d97c052d1bc34baf068b8f514efe43b482a9750856c345bc328c99bbc66dd70876c2f3041e939861bfddedfabfc1f965eea6bbd6ae60239716ba38b35078868c25e7d5fcf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1534e1f2d2138d0d21e4ff5b75bda916c9039d886e1b16a5a6201041e27a43a897d82f759ff16de19c370ada18dfa93a559937268ec92b6133aa4ecafea86bed34c8cac239df22f74e7b91d82c5462ff4560731b8e5da7ac6846f5e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14dc3875715124a6d19787e95522cc949833cc6450cfceb4654776cdf874370935b25cad0813da65a041644d6f83a277f446ae849fcafa0bc616ecca48e190c3f3644a9f31b1c000ddd006d80e47d43fd84a09179307e5f346e2b90;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b686a3c285190c6718ae091d7400b05d791b60713e928afe4b5e5fa8835d44fb42896bb6dc8df2c87163194bfaa89b59bac7f27da4006410c0fd610e114f62b7c83eb2ee0173591dabcf420f5ed259f3ac434a84854e7c015e79b8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e4c4b806d11c0456ff829d49e6059e2ae2008093f0895e5557adc8ef5b17e9bf4d66438a8df5050a8493b98e0cad85b634e9201d4cc761fa6bf03be451864213a6195b3646a638ffb7d1de4faba4d87f2998fabfb2591857d614d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6aa73460cae909692bf4ebfafb3ba74111299ced43d1aff92052681251f35cb2bff6d860d69241bbf2e2ca0273e36f1fe924efae4d2054cfb6710942889c62e8191f78b36890b727607fbf9764fce78aee7992439c4b366a42d6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc51437a8e55e9094f96c780bb67d7be6e5f59bcf54e786ffeae3a201b44fb0aab20b9d40450c852c358447055219c75ff452f50fa7e2da9072a977aae49a7639a8b019651ea87bbc9b2d550770c51b8310b745320152e339f875a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbeaaa9b5e1d890e0147209b81c68e512f2615a1cfb6b99e750ae6f2dc4663f905f1444e285f0ea10ab4479d5ea10bdc1a74c0dce685e4b9222182ac6fee93632a2d60b46539b223d073bbb598778d225fa50aa6d9160052626ed62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9f9d88e3501813d36eef2a83114d0ef0a1b720fe72af6d467cb45b5966bc1c0ff77487f8fc0dc89e32643506ed9578572c71658765ff4fda76224baea4972b06cb9c8e0639c20d69bceed333a5a3215fe230caab9d4c8242d04f8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cafa8bf36789fdf8b273cfa676c463d74bd43c6e639c2baafc7db667703eb4c8c9a66bf6ab2d953de31de518f00c6f67369d92673de6560ab57c167a920930231eac9516f769e6886b43869e56504c7850dcc52fd7d7d2b9ce984;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1477b754b07f834777b48dad6e0547acf615898cc0b46ce9a63641b6de68d7d0520515dcb933e40881702e614ed6b12962b722733a3d964c2bbecdd1050f6a59cf7fb1317c1aa366ae47e901108a33e2aa3518d11a580984220312;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18984a6c57af3541be3248a043d1ee12384fc22bc2635ef480e51463b8143c3db6a3ca6b0242b3710ed3535a277f37c3cc4c4f386f468ab18a293ecf25959c939fa7348e94ed83f7170e28cd8556921d3f86edd315326df16dfc400;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6af0a2fc5d195fc968679f28dd8d4f28441b9887032d70b2cc47c7b9ca42defa23dd41d74cbf2633a2b4a531fd2577b45699fe8565919a56cd79e6f2957e642778f18d068582b82ad2304ec0d18e24546fa930b1356a1fb39cbec4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h781147ae38e69b226a9351e703f2df1ba5f3d21296fa15f3aaeeccd900758885466c95a57b84601f92b0b35ac3d35a766a39c5785b28ccb68c688297e8056219aac22800d9acff77746b63874881372266abbece0b1021922c4e86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194a06f921fc0dcb82f95664dbda9f0c93737dc54e7ad0a9e48b6a12cadbd80e90e3f90740428ed8c4a4e5f740289ed76074c4b93b4c6a5b793d254da5da640b1c7e6676d461f5fa5ae34fc7595cc062308061db4bf537a923fb86b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1792e2aa5eccbbd9c0ed5d3ea337c68f845af6ff03c83c59a8209e72d2f626d7b0445fe9636e3986d563ba6355a526a1d31634bd684491054135a20a22e12082add83871ba927056a2a1ec11e78c1f7e6020172d3c111b0c8885bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h530da204d2543a723951d09f0c2f707ed0a6d0d86c97320be4cf81c50f142904a5d306a4b8469f579479dc4fd4b77009035d7ac7795a77734bbbd001520174c43e406ff7a4416ad33f690756a51dfe3bb22401465abbaed02b96f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h370308dbcee3b4ad84dd18716518af08ad15c2d26db01209ba7016e7fc19c80ceff180b9cfbd398f378ca35996ed9e41e2db15dc7f278006286f8e3dd540143e0ccbb997c40962b5945b9508e661d883e990e4b8b9396766f405b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb0ef9033b6760e84bde282a142ed79c60b2ee3ee28fe94f384d1d9e87343c920a24b435badaca5afa4bb53561a903110af678e0f2f8512db60cb11039c6942b02e34d28a0dc3733de72b1a4f0e6970dd518ec274aaa2d202fbec4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f49e55eeb36466d439146ac36dd741563dec5714cf92108c7241463a85cfa7cdcc870bd6477c8efe63c0f5ff51e198bf72e617190aa2e6503f64813bbc256de054b97e7a0566d979708b74ca1bddfafda4e2608d0cd3d9024a8720;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc26ddc25d68d486487920235dd5930dae5a58a04321312700e4d8090e92db42abfc8edcc9599e58f99a4328927f3b9d39ddbd63445f3817ded3e865ab54f9f7c2dbc43e677973dd888c5e8c75097222f692f35acc038770740f8bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6e242aae3b99622ee9645aa7f5e3a7aac52df67a9e77ac112a25f4199440d4035ce0aca52703b55a978b2648faed1e53c8eb7481e5861d73a765f39b99e591b60abada903f92dfa4f8770268a072c072844664afb06ad3cede511;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc849edffb359a5f6d005af081498d331e474095db007a5e0a5a4ef732d127039e4da298f0a491626f3511863936e6688f02caf262e10b823b42c17a8b91ab558642a0f06db8601f0a8a8bf826adcace4daa1e3d2f21f0c7e15aca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8da8eb193d3881da7e98cb6022583d66b46604964d809d33e6f2c621df2be2d478134c1b24187528d8ae9cd88492e8ac5bb40cf396773d46c5f51d627bd82e24d01ac896cc630fdd4c7dfce9b0d0a7f04fa3a9c667e57285c9a42;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa3b53d33a1c8820bb23355bb29e2ee6851718bd4ecf7daa7a7035e25e23d02060a69cbb21669e1c1f8b5bc90c441b8e935c2133c4760ba0d43044062063078ad96245c84697078ec11d6866e30039728c204b5951254e47a6982f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170886037c31a0a78aed487382f1276126fcd179d592a0870892c3892d94fc247bdd59594c19dcfc89b08b292954f3ac02799d520d985b7b7050445a32850a2b4ed7111f91d72241cbf2a403b1d82d16a8a846fb59440dc8f725f70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57ba801c6f6698b18ca7d79e875203325950cc33e695d57477d705d2fefdfa0f2025ff69560bbf4a4fbf3ad747b4533538b8f717b19592e785fa7dfad2daab3258928aa3f5de3a0143b260e1d2b5ecafcc9a7385d63f85bad71df3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h281049f6073507f634905f911ae7b6905a764f214e164ff9a379722e1a4581f8ee1cd41e152fe23c46b237277873c04194f1f37c38dedde2cb5c3cf7f18c9979f0652d8671318a7ef694c13d73dbe9358c3cf16b7bc406ba75cec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a080f04540b8b01a3080113663ef0e48891528398456978267419c564193c33b0694631a56e648869192157e16cb778fc3867f2b00a9084d485d3b9d35e139c8dae7e31a375e1409624264cae599cf6b7d2e76c6c62f0700be9ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13540277a2ef0410de58f0dade15650ad2985540c8e9cd580c6658664d0ff96584a3d4968ba9000b9df33fb2736b24e2a3254672b78c15189abd8712a2cf1869444637865100e75805a78ef6487e0b31a9b057c652d1a0d022f0546;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153cc67c45be3547504b259ef27f7f5027b0de44c1805c63f8ea7f5f81d5cd267a1a2b8dbf09823129bd65eb22ddac999b18d711668837fc07e28dacb175fc954bdbde4ed889feae62653c0c1025e1e287fa08e7d17da0739cca9bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b3ae523574a723d95d69065dd42ac00f276a4d2ddeaa6aa22ebd090299aac6ccfe773a984ed858cdad0e0596ce5341135dbdbb23e23edbb53d1ca7f0bf291caa832a821c50adf84b1fe4d7d5a38f2a71e702b0b73a1dde7b1389b1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c9a01a451c21e4d8ddbd09c608779e5550fc29a7efaf2543dc03fee5056385150aeaa62559919b2570d5f2c77b25d60c8625cffba4cd48e927f8a029cfb9f807a676ad2445ce1a6b42f962b6022bfc135b8d867ab12ac9b195d5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa52e05182348f1a1df34e2f964a2a0ce56c4f176bae94cc7aae973bac2c1d72f844b5090d60b81f1385d4c01dc3fea5c46a75bcad0e8e12e73d7303a8a039bac6244db93de6e17ef054abe7ffd425652a269d806941dd99de2b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d6722eb78ac3db439ee757c728559c08adc2e3a701ffd8f607d24254a49a97ce6003406967be41af458e8ddcd38a70ec024be01f2533c346f6809d7a63e4f2c2e0f27db92926b975d905e60369571cf63eb4cffef5f10d5896377;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h47126517cbc8a8d71c2b4350390d94297e40b7eead7548470c152200f7df7a998898827053b7dc76449f1a5f16855fa924a7c10f750dc0268e0d91ae4bc0c68c4cbc722775420a29803f9b9678a7a66e743ae0d16f40d24e6f39ac;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b33bb8553d1cc63f0281e4b8a2110b226d1a73baff41f73dbc493154442466b62cae654548921d563274afde3b97d274fbc934cc617e99fed3536f917258e286a92dda149ac01d4419dcf8c14a22bdb7a56ea4453d78a54dca85c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h150963ed2f96f3faca29a885eecc327ec0721cb027927e1c453edc993a5cce7dace6b99d7f3938907e28f41c470c62be8b92e7bdd4f6ce753e6b448e0b4aa20e97f84aa356cf0d0dede5061ae9357a409842fb59103e6fd09b1664a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd01abdbba070eb623dcf3f14dd845ee5ff85934e5960d9e72cce4894b38ee4fa2cc1ea3c29098efb2212199dbfb7980e16d7a72da08d66290cc8a3868aa5311e85427f4941575f40b166923f94064558e2875151edd1f1e800fe6e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c2e988dbe17d374d8aa0ad04e0643e41abc8fb8ca3e9c0f5c17c6fb5b7e27ea115141ff0ff9fbf0cc55368c85d70777c4deb589636c7c48a55a12223f40ae7da088a27f31e3b92fe6e6685b7bc684ffc04af8658f5344400b5660;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1921656c2d5b6688744307ba16314ae95d25cba7c25deb03caa01e8021a3ea3b848addb08eb8d9bb41298baa877c76ba31693e2ac294f83f4ab20e589260c3c93b24e105c4e9c0d87c764244347a69b495376860a272a5ea7ac736a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95245787b46e42ad8b5074309218d3e09e327ac14f788bae3f346facd61dd2562c336625893da94b02223641f07d03eea5271b4500bd633fd32368ee448202ab659178b1744c65a9aa6d5f930f6cd074ed5d2824473772063555a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8acb045cf4b2d140164f372f547ca5951b599e1b002457ecf872f94814fa98b8d9d4b528a3c408496acb8396d9f7bd6c5f53f2a965000697818eba92e4c682721bfe389e263352be417f461390b5f8f759f948aa5f9b18a51c2c13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5fb1247ba1a75102c6e4faa69cd05e3cde1ea35ebbe7e73ad8d6d62a7d87c4f30258a07da0674cf2d46d3e6fdf1e76bb04e372e7ef7c2632e0c0b31f738d7628540e9c770df88b47e932f19ea8595cb574b464d986fdf73c097951;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83361393d10a2ad386280fea2b7909b72cef18275c8f4a435fff2a53134ec0b7d3eddbe03f8b0cc345d2d943246fbb44003592fa8c2b988c6f2cf88c2dafbd3785cd2f878d0a90971e0708a9f3db75fff3492be9efb5b43edab7ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4699a00e151aa2ee1939d8bf44d609ba68d07a7b5aac0fcbda4c49ada69e407b26d205913118abe33cb0ee47109ef64b246145322a5cde681e531a2591de9d00477aae5ece835da72fd63aa29f51e5e623435d3eb00e28f0946c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0154da9603f5cca36177fabe7e417a0833701315a6282f2f470f229edba29236018f4de4963529c428efcb50b3c3fd0adbed1b43b98507be8b0881230e1070e76bcd4ce9c071657718b350add07546e68d296d017999c15753314;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb864118d6bc94c059590365ac97a3d0d40f9e7c784887a37ca03d3915c16cc5b442dc429162c6c9abe8bf83a14b362463d1a97deb6ad296fcdd6cd1ea1aa91ab7fc1b8dee923bcbdb5d15dfc5b0ef0d876620f45c21dbaabcd55cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16897fe58200da51fd88b51bca93d383a4f45317ee6ccb6502a1ce7fd82e423a2403f71397d2d303f5a6640698001ab8d902a334ca15700a2f2faf64977bd4ef486ca19c00674c5a57671dc5e9c3b41e29384787b41ac37ee0b1181;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7620e1df771a3427072a633f96024e11479d04acdb6f4fd4f17e382bf8565ae8d46616a37809c847aaab05341c2373c676fd7d569617a886c8a2957a40ff94893026fcb290eccc5be304dfc412eda82e8fcb8c1fc536f208df8287;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8f8cc696cf88cbc8ca48f7f22662f23fd6bdd39078d1e02417f29b0cf48a1ed7985df8a8c79be134fa58be6fac86d29f063f3d3208726ec463c53ae7b0181aee5206b0f2bd87253b39033bc7a4ffecf1fa4b3a5e53c154f93d6ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heeb0ea6813607c2950ed428d54b7b046f620439836588db1271cc5eb01c420602060ba3212d9085020580058aaa6dcb97e036009c3604e3146bcf993be0c0e0fa20ef7a208d5ea6bc00d1edbdd0f8748a16ddd734b0b1de497ed7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cdd59b552dac2c84e8027bf312ee99e132ad64a3ca88971d69eb19539c06152f028b705f72222c6b88d38dabd002f680721019523fa9106edf1034c66bf75f3340ec89036bc1ec0d83362f1fc86f2244fb8f2408342237858ee42;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133a226e0527a5cb8d086e630f0c6d52e935f134890fba11005304eaa71382deded5f6031d700a870ade8ed948bf6b8e926f7a806ba1dc4e2175e32a15c1478577b9862634faa8a7e8a511ce9ee7f82b5ad210f13226d18e8b5dbb6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10656abf087e1aa4dfa18c39dea055309215b91f5d879f0948702ba08137b0a9956df60fa216245a8b389d85909688644fda3a5f056be665e81ee99cbc05cb4ce3ac0c608fb83e2ed532fc5833c2434804fbadb30e9c5e5de5b29ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h259b3f2a519a766127c1bf9ac73a0df07e30520059fc4a41fbf93b904fda7dc8ceb169f4ed5a78a94b038645ca7c5cfd81152d16a545006b8b82bdadac6a0eb8cfa869c03624a7d0624124987a7cc7706cc130e65ec35ce5c873d8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8537d7009b8f6a28c9bc41dbab70c145c0db1cfa638e918052b55f82e443938b98547903e749cdd783d4c2e94b6cf5d961f3f07f74f4f357143dc6cea26e6d4c6dacdea4a3372ea991e93763026507fb34a012f9e5a518b217aa2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3f65db58b30ecb7a73318a165f5c18435cce6cf510022f320d11c5a7f27dafda05e57b7136a668c3c1833be98bc3dda370946b2858cefd8cd5196472f9fb2a6e3a52b4f5bd42e4ecdf11f52d2a586f60c1f6c660344f49ef277e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4dd9edd89ddcada7ccf66966c057b14bffd1c3f926bf7e05da885f354101055a0144bf1ccecbb51558b2cfc6b68ae918f2695587a5fd45a40fff3bff46acd19cafbc3dc7b508129d1c409ca0911bd193f3ba223eb7080c85e057bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf7c4e2b3f738f8100c368377aa8c42c65be72097233f3ec69c69a88c1e6210b58f463ac19f4bcac7ab722e06cb69c107719b1eda7d175fd784272a9953d7ed3d5dbf139954ee335bdf921d115fffe12fa2dc9547f482e3f0c5210;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c3c5aa61011edf165082c3600600bbe2930aff4f72f6067ccef853a2dcd3263f5a4c45d00106c7b1b9e3560a66e33d0bb235a88f3b3cd571791ac3e9fab25d7ec60bc8818d4479ec76c732328bc4790590eaec8628945f936f7b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab954cceef6c883e934f663f33d42b20964d38d6b4117c2eb7d2144376ffe2e21c5a763e44f1ce28db4bb8ee539a0fe244da2889b10324a51f22476ad00d4f8d36ee75fb49c4c44e0966fe17a1789a54bf79ec15489c9df3e99a23;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b877b14af23e5a2fe0fdcd29750a811ab16c57dd72266e31edbd4454faf76e6df9c44912253fb6acc0c19b310ee35b647cd543ce2da0830e013794f82b4a8d28d66ccd335f75fb7ed4a5106c4b7ee4fcc6d80717ce85fa0e8bffb4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d2421c5e7f7a6e2afdac95b5eb591a537a285577d1f37f30a47b3f45b4c8135547d5ec76344cd5d20bd4209680ffb42940b56c1cf37dcb5599050d6efb3f660fca41223fd45f9b58fe0acffd3651542e9dcacc7ab01512c48865e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1736505059e03a40d21991e6c4976f66cc9bb566bf427e284883c1728caf82995e4690d10ea81ddb12ddf93abb5918c347987c1dcf7dadbb37eed255a9b2f8a67de6c6faa67f001a3996feff59b6a863c6740cd38de8fccaf569a9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175531822a7828152b27a70010189fd706ff4e90773c09ed133c87c1e9152dd759c0d90dec0f24fe2b6730ef48ed6168f23b86dd06e94dcb32fbef512166df894007e3d07f102dec71176ea174a9d490d6814262c71966a12472788;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158bda157fbb6486be728e1be3df742bbc51c92564f35e965f321ab86de90f15e155552a561896bb23b83d683d279a13f4262968a0265557d666627f8f920b7faea4ac5007d1214cb2332bc984ffa2c2d5e21c05ef351691a658d8c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec3062ec9f3000bb07cb64ff3651ab10298ed6c48344c18cc4592b5a24eb2c8ae642f3135f00372442b806ad0e28c81d6d5e89dd0fcef9e7f7935a736480a99fbb1a5d77ed68a7e3bfb94e43b1f91721a1ffc11a0ccc4ebf839390;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7ba69a04c20bbce4a9a9b162870b39b286b5c7b8b073850d7e7f4e5cdeeca1c2ac5b57924fa6397a97ad20f920d9cabb1201cca68ac0cf69fd7248a164a3b5666a1f140374db322e3a490f5defb2a2f2b7061d03e88d7b38540b7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79cfb4214f1c8587956e7db2a1e7e4ed397a2cdae928aec1893cb13ed986fd2af81e190284e26462ecd9ee416ae57f5da71458aa7582ecb308f13ca035f24c9bc4bf71383ad954aa114ecd6469fd39c77e3efecfdcacb2bf2f198b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2106de6fa3fcccf05aaa8b2e7fe3b291a0bbb2d3a3765cc1a6a35a41b5fae8ab9918db0b5cbfd75941cf221de26649c5e8e987e3431605591ee8e385c24e15d919e0b24a1964cced5aeb450057c94f6f11c0a11cd65e776fefa86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb411a5cd9e4ce6cc5c95e7c0f85365d16fcdb04acd2e44d60c10d25a4272f705d7754705d0128fb4bb939d577078ec322aca0cd29495eb19e988ee023b51b572441482f37f6237e9a8051a9aaeebfb33270789d98304fd6f3b9cf4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb876b574f2adb9a2dbd847cf20df51a962816d628d64e3c10fac7085daaef8fd085f199425d59a5692ac57a39363ee154ee51d0995f9847576a5276aa45517e46f7c05bed716ffa7f6b38619be15f8d7fcb9b27bbba22b9193a94;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h225cc3c14dc18acd7116137620f9d1baa2e69155c5d6880dbe91ba60296fd1fda342fb89c67b82b434644e5708ef6d9682f602f406b985c7455458810a0fac597354c6f478d4e8e805f0fa5deaaaf38c9cb58ce9dc3011def6bac2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30425b3b1e58ab854e60f20feadd9d819aec15375e06bb14a3416698ee95462d8ceb2dba8b347ede9a857b51bd21ac1a743a5bcab3ab97d1cf022058994e895b82b786d57ce0cdbeb61283985dd3a31ce4b5266ecdf363413ce4f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he61d5a5bc25f64d3684507ef12be212163a40208faca087da2a7833e7beb70ff1a4276e9f16861a2b1bf67376eab16ddf19bbff5fa75ad91bcaf9149af7c3783fd95367e28d91f8ca5326e722a4ae3f424ce9b30ef032a9146b871;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1528aaefd3c39edcaa05a8ebfc020fadf146bc8b24a489cb5fe305d9f4e8dab27470268df3d02f650b13d05b003cc8e0c4d9f1f16e9e1c90b01ce54df41b9035cb67c0187f40be0586f25ddc2ee1b455d5b688f78d185ec6aa6bbfb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbeda87b3a1822ef75a5436ef2b5ce5b4468216062ab552c10010855a2e4114a4d719bdd868c326dee37f3b541940bbe8dcba994afd4d2ebebb05552f925b99f1a2e162104c6f696a99eda44776dd137ea7dc82d24f8d1f9863de2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee2f9fdac9d0e551952d3f4c78108ba6f6b82c9158c03cd600e8b04ae6470e36d737ff1ee28b5939baa7abdf33ce703f91e86bcddc2adb7624c21a4cef3adf5ac3a409cb2d41e7d4dc781a79c42187f4dea6480f234f27befb1e86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16df320454e335a164c291d2bdb6543329ce679935cfd61028f5c550247b762a99c745b5fe637efe27298a53babec1c1f5b6732fdbf9bced83690fcf22536b7e351fa1362a2e3579a504b1f5ce898b85f1e683a36c4e05dfc399806;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbf808f91a2d6cd13f30984a66c2fd8a79eacab6e7ea2dc91423f07ab56ce4819e2bdca9d9f9a6ea6e40603eeae27430fe895f97a83e911fa4fa16b5f6c438b0592002b85c36ea78ca8248a1f1cb89d280ca279d33da469cc226e2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5368028b937fb0f1cf07783fcf2281cf7094988e132c98690729b6530d53450a9c9f6f7b696d40babde95848161a11c32466eec81718b660946c6fa18ad680b651d276be84bd52015dcc0a6bf77cda43f64ba402341098a6785ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ccf2a2ac8fe84ecf6269bca032898bb43e6a4f1415b0c11681fb8384aa5c2f8f1779a7af1ec275c00db4d7432c4c5da778ca583b1d021b6bf4718087e3f572edc54e521f90211005e9b38fcc6e4194b5bafefc966b4796b668dafb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b88d32c56368d1d43df144e681ec637c569afb0848ade3ff222dff488c75193903806c5fb0eda90630d26395f79c89bd484325adcbe3c8a84be5630dd123b752e6ab792255182d19732f902b7268b6459a175074124a5743a92995;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17058dbd7f4285662640fcc2cf4979d0e123ccb6b3e3291c2da79e004386e9c5a730de60baf349a83c593cd28231236ee64c83829f192c4393c544c8e9a5921cd07bc5ea6af50210bb87eb57b677bc578f2f6c9cf97d1f31152747;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12633639ce9da016dc61cb3b1ca5fdad924395398df8c6910d919035eba1beda6ff85dd1051c52c29b89c9a376c23fe670239f298cd73dfe6ba21365cbd4ab38dfe98d975b00cf809f8a37f188dffea2fd60c7dfcdc18d81261246f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1099be9c019d0233bd563c31bc6948fc1f067a60f41e09602270a6425a958a9839b5385e1803b50a4fe1671c71a4d5428ffabc745bd6949e32fba4623daa977c79578c611b949c618f3dcd4f5330215a2423f7a4660fedd01b4254f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25b63788b81ac29a2981fd52d3c4d8d8595abae6dd804f3420ee29dae1997f38bc3237b5fecf706b8d49ed4315ffedbe24ab4f7ad54d539d774accdb7cc03ac219136d903ac4c82b97dd94179d999d40b3e2db1b5a700e6ef82ede;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e90c35e4b7bc49372d21a02414a69d5e389ed05cc89b3f36661de5edc292a316121d08c6cfeaa017574212f64aed2918c0393bd11a534a4b95c45c4a4d9c1d27259e6489c9da821577e2ddcd9834223418649e235c18706c79d78;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1634eb3610a6c4d14d8a8b0fcca22889318d9279eb0e856ad499024ca824e4101f1c84e03ca48ed68db57dd472faf642d374c514571b966b5686ccc1521f8ab52c32db461e2cec718d3ddc3e7f3a57933d5129552330c91823e3679;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5298ddff66e0e3bc04805b7c615b5e4270c3ad7ec7e9d2ce4df4f1865e6a9488d50302cf3c890bb2bcd27c940e903b9fba2ae2b4b33ae89be604434fe7f1bb3aefbeefe6584e4470d9c54b5e523e996cd194a2c4349bd43b560221;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac0e4fe16a96b1330988c003ec9549abbb38db94e3c8ba6d4650116a118873657429a6128deba4d54adcf506db1ba9a490db4f479e890f9734c7e9395775c06e1027afe7a8824bce076301c54c8fa385bdc33b199cea2f8e79a107;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c0f4de25a4d81e57ec19b0b2c0261539ee10cf6c0dd8b6e01af4322e22affd64d7f0d69cbdab76c971c1b27dff697e705ef61a2683fb02397c31a49e9fa87c188f49f340ad0235a8fabbedb455c366cd642ea8088232c70d9b30;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf916f249fe3fd35ccebb2bbbf99fa266d99c2bcec2e12b987f20faabe39b7bf4f1c2f17fbad02b29f6a82e3f45da7786de2719d0cc2c3076595990fe21dcc893ecbc6e5d96aa0fb129df32ea91898064692eda9ea243f73382ddda;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a3f094b783f0250fb83656bc5cb07a0194d9a1329636151cf1b278a854b2ea80b56fe99fdff3d2a4216ec31b4c56a6abda96f80d4c0adbe1ea6b59508653bccc80ac06783ccdaf264c545184732b126bd0bbce5c82c40c319db42;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185b12dc8b5719d2d78147b3500e763b621bc649ad17ef09cff0ed590592a99dc43d9fe47eec44e0c4834246631d08e0afacb151c1a606e4fa20e61b32b098b43f2f10adf8fe90ea39522645ba008c2b64e5d66f30b2ed7365c3db3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1308682b38ed9878c34576eb4f32c116c75112d4f36b6e26b57938843cecfb1a9025c3357ec9098ad66d20e4ee73bc2b4e2c06575d0407349508554e096e3ac8267a7ff1d26f5d2035cab5bcd06d30c280f7d99d047bd60da27d281;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f758464b4deb37f64e0124328b4503268e91dbd786870284797a1d783075ec22bd461e1074a44611548a3b133be7c33366cb92dc3b1567d460ce1d94e26fd0395aa67e44ff8af6ce0c2bd28e8880f75462f64b07aac5a5548abcf6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4987a24001cadc0e6b3b61f15f616f2df362069e6829afec0175477a035992d030df03f82ea2e17cecd4fdb21ce2a0e98f0ca65f41c5cbfa300d2b14f7e89abf51f829c92ec2307125dd6383c0200ecd07ee730b4f8b40d29c8e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a6c48cff81abbaf650e374d34e92b3ec4ac15022f663dade1d16259dd6e494c2287b58f318d17f62eefaa2583f455570f865cad850ffcdfdf63312493816ceb7f066efec85888000feb03eb047d01f83a73ed2bbb818524607f2f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2701dbb12d37d167db62fa6855a954f83d1518faf9e6c05e659adc73e871e86690c830e70db07892327099e4164939d0641c3b612895c52201c223ebd16b760032033aee35381b9fb4f990cb9108515f6198a7c664b917c9c7092d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c6aed9eb45adef7f44f23be4a3d1556697af428756470fee61d199e550f3db706fa99049dba3f06ab6459043b7b0c086790468c36962ec30072865d78294d9978092c8d86a612b738354bb690c38ed5c719ce48ebb095c3281715;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef1aab078f46bcf90999df27e8482ca4ae78ccc74d4d69ab9f330f38e8754df5fdfb799a4d425f046a05647dafb1f5844023366ebf3d09a75a89f08871bd09f5b3ee04627b96dee575f8d4ef5258387dc03f4019d0797bc8996cf2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7decaa2a12df85604017f1cba26223227d093d57308736c32047eb449b3de786e7ea4b6b04074616807de8887211ec5d7acbdb89ed9cb9a33292d6182af180e1a629f680aef677dd40b75fb05ee6400b128e2b387bd02640f8931c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a0780fb711bdac885dfc6d52db3cb8c764ef53710bf6e0f5ddbfb5599d82d6741b53775125c05dfe934dd3f015db796beabfe4740bd409bf7fe1fc33a89b5775a24cf11dda9d63664e964a53ce588a780697015ac15d51fbcb299;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12878eea8dd1672f996f6caa20eb30aab310aa7cf121b648907cb965323b4fed0a09b3b4fff91106a6bef128a78d53741b78923cfbe6273455a9146d2735d789c8b0d13dcea8f2dd76fb7d9d5031dcdcede2a8cd02ad1bfef2ed035;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196affb9f18e61937eeb1fcac10ff493b3949f3301fb9e1b00b2b3f0941cd96e7b8e1b88b4ace54ce1cd9765655ae838e3eb0892abaec6711c6e127564fc965875941fcf2f2c8f58b33dd8660f4b0e951439d59a9f144060853e2b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1023577e6ce9764a21062cb2a94426a77755e1797898b6238efc75f753c9b165897f5e7024cdb821d39115fb1c11e54d9c0ae18e4a04d068e03bf36effafab8326c4d4178e03f973c5d2a4a2b6aa6fed2327126b8977ad629f039e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42e7c3a2bf4072f0d973e6bf07387a7e9e1c98aa3e6593a2051be4a1432c4e39af46415ce8469788f170870ae986fc6b930d26002035248e11032bb1cf98a0000401ed8a8087f6bcf5f1fff42583cd811b42602f8d6788a29a401;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13805868996058da06f24086a38602134aeba4de49eae2c52a3af8f025f9aa36f25b1eedde615121ea5618019bab33005502f43171e2909179adac04b1b24aa29a952c09cb88933fcd1a0490d8e43978e2733932f3f57be3f62cfb1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h626cd632dc47f4874ea0761f2a58da97efb00e6faf9c38b34aee7ac42adccccceb5cbe03261c6246311652eb93a8ae5d33aed0ab75e796c0222ba6447db5249815dc04e6c12bc6a4ecc6aec98c725b2cf411bf45276981d881ff53;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c08d3d2b45563417a652f5299c8a4fb830b6900e79147c42bbd7e731040700d2574f8038819510c76bb1121f828875372ee274f4d9d18310741a0127226217da676ea352619c7ae645f4dde4b699b75d910c73b4d359868f425f20;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5089fdf0038c3eedd36c7ef5efab3b395f7d3f512776c0670e0f9160d5932747b5cd740df5ed8bdac8c2cb2bebcb33a51f8c451742b23ea3b0e53131632aef88b767cd7514f0f7c3fd713014676833bbae850dd187cd36d356d0b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b91b1c749bb8fa8e1eb9cc9b7f23862b90637148f6eb5d0016bf8d5bdfb21dd3ad6edcc96598a93cc1e89cec809072d718ac03c261f702d5ac116b918f7dbf8a78bc1473e208d506c5df18ee2031502fa512a8ea98d21306a6e9e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h56eb77719d6a92868e9b30b8b45a4d3e9576b68f4eea824587ddd9d13851778245c4e5e2befc8a48fc0a6369d0325780ebd36a6950d189fe3a5e06ac3aff25245f40832479be27b8e6c26113beed72dc7ff74b3e6b751abc1b39aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb22ccceb8ff973f8df170036c8665a00a5bae993785dc1fd5cea9ffbbcc83cf037d00c5cf6220cb990b3a3e52197c451deab9786182035b181e600702340158813a6c68fb56df1b6ec15040fb81cdf00dd82dc8dc9252ae5b58237;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h32943e38d093bdce73523d5659dcbbe1bcbc1a3143dfca35613b6d7c6cf6a61b526bcb359a635375719cff2da085b441e85a50447de6fefb7637b832fdd5c01372ceab29bd54dfab755fc96dbb11f64982253609f7c2d3c2b3d47a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1429197fb9ce415c39a525c6a78000485830a16f9ee55f1dc61a8bc2a56502de44df4d2a46c08da4f51827b21a0961d1ac314dcd3a7cb92b3276e9f3983f270557ed19f1c76e55757b210ddf9681f934a2142627d34e3baeddbbe7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'habea7f34be8d0e769f27d96537e06d919281c6bea88cb5d57d7e3cf65603663cee7f5fb7949ccf9cf435c8b608a0cbed9f76a181b69ce3f47df4b1122f093cdded1b1e730c6d496f6b1fe1c956c89a4e4ddc8fb73c480182cf9c1e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf67c504a56374c5dedea8e115e1457bdb55b873a6c984bec13c2571eb256a451348a5c5ab0a5a372e64156cd5a314bf7a0475e593b831502fa41841805b3cf9802fff68328f0221c6086803e10899cc1fd9c90fd4279e278d0d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cafa5934847a134fda018310c498a7af1a0d406c79a44cc62b95d138333165ccd5a279060695fb38558bae22164385b750195db8fb93841a8505a8f1321d3cb7a0962c53d37c7e1f508ac8e8274e5d610e51644d281cf31dfd3c40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12aaf195395e7054e385b76bdac20cbeb05a91f75c936240f343751b820872861ddfdd7158519858d00259c576306aae2f7aa44657c2a13926e8c06fe140663c7e0381574903581a0a276c01a912a4bdb69077ecc3ab1a171473c2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h920f38f293ea5b89ef39d70e3694ad1457a9d34d95dac7eb07c38bc3d2f5a2b41922a4b113ce7f37580e44eafa8d5cb6c6071824bb28ab012d01244ed2c4c92078cd3371d96a3953956af68ecd8d7cf7cc2dbbbd0521395b97e515;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8dd645215754687deb96ac168c2c86c0031dbd0fea0b7e05eb7fba5287c7be8d605fac29f55b0343d390c7c02fe7fbe3d15766a41549cfef594ee6aab7aea49333e5bb37e6f4c5c9d07c9ce47a3057be183cd6c9b14aa4b04e028;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha19a666da9f82888df6c5af7864790772b7bd1f54f88b4a4cf7f377ce4bd80edc0cf73c280e17aa17152049509f6c140eaf1b0824aa15f54ee67bcd8c23df60c5bf164543eedb841a2de72efa9846f1574e6419792db5da87b321e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8ea5f68d9241d2a8e1160c3c0da224c47bb7749898969b9f13adb695010c17d3bf8068944dbb52688d5414c58c2df97b658aa424822c660f6f70b53aa50cb397adae21ebc7eb934bd2021821458c1f77db7d3002a41034811371b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4afa13ef99027956c928ed6708d958b8b868f26278632f337a169d619a5bb0e36dd7e1e2ae0c56d4f2626e264e47d90eaa4f980b342037d6a672e6beeb4dd2da91adb5f6f442bd57ce79392ac5876999510fbba8cdc71db9df87ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1982950ba74f6c0a3236a6338a1360c4392a0c29f2e7f10655c4c9903537df9b74cb95e64a5ce4298a75a950b93a0c4a7a93804dc173af0ae8b92d9afa52f6aa393ad6acc3034e90e646aaf9a58b0a4cce1a44dd9ad8196e2fa8048;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80d3993defd3cfdfcd6a3d59149c3450cfd6500017c515c458e50e2d74b4f02e5dfce068fd16d20f9e87206932d66c5231ae334cce1f4058e702d9c92c907136aff01cc6ea026b889c22ef8ea0efc96b8ca335b3a2980c01270672;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17cdc7b093eaa5c11712efaa19f735c9e84e80e9c3ef38cb86e8f7d8420c85cb91e6d6187d5884482e1476fca9ce847f045661e78845e18f9a4f95e2a0aba5bfa937989b1795ddac5c42ae5d751b77392f19b946b9f9fd565c1ee31;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca3c668d9fba7bb068b081a89ffe0f23bf6159a468a05733bd35c6ae5d7913022170b093d008533e26d3ff40d768ea64d648ed2f915ebe6f59aa4e454cb4e3701c62ca16c3b02b19d9eef9010b0ee68a17c4d96c4ee5b8e8c79b6a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3845f5a32eb05d7bc7d36e23225b690f4a728f2af27e160cc41a2ecd139fab122e467bb66a8fd464c2f7cbed2f447d2687eab9e78b1d8a3f6d8b8dfdfd75f2f6f7417a77c97747e79d3380930c0fba315172b773d33711121a894f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he93c2a5d5da2e67cab1c81875f20d7687c926eeba718b41e396b5ac905807dafeeeda8b13e4a864df6347d568a8413f4fb6c61ac06b3d4729940dd4346eece40780889869d6fddd7a63fe36b4007bb83bf4b5b05e3149ac437c5bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h130079b5e0a0bfc5ff7582e6dfd27d6996aee47120496bb0612a3af9ec440d98081cd7c2cf7775687492edfbe0cc765186dcca848642873ddc04d27064d35f131b1d734df2468d8b513748522be6ee3f766c9de7ad6625ff2814e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b60640dd3d0cff922a3441a16e4d016191f774e74e83e93bc8c86c9d28b39402e69efd1b566204876b513aa461b97b3f3037ac9783ed9f05f1e1bed9adcd58f14133adf9618592c960dd31588a75408fd43532bbb46633dd9041f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c979f86aab0d15f8fdf9e949cec362c064915d8d4d54a2871cbf7cc7d4bc27f1c2863138ca5f54140f971853eff860365f866cd9831c2874fa685ebb1a8b8607f4f52dc10aacd69875b6ac94f3de967c83001260866747647e82f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4742ad5599aa22f19326b1c7d4544a48d81d4fd1d1c6a4e51748a269eac0b477e5a21c096655f36b979d4fd4002f3eb4ca6d914a930c2f0c21d33d9801850b9c0624df3a4a10c6cff065d38386708bfbc68ceac9ded05e375657c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3e3711ae6ee903d2821bb7106745429c9180b9d184247f019ed0788e60017954c53bf9b9e54986b35a25f06d0138190792b2530929075875b5b6ce5d8f70d3bb7f3e10bf2c3e1b12d6a5ba4d4d9e815da07ad3b2becd092a710d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79b176e3502ea6f458fb0a4e99e1351bc0e70aca441d6c8c5c9fe730b075e5d52224abdf610db699da978d3ada9dc4e43ab77e2c0ef306dc3a43ee1b2a6f3592079b20fb407c21a08cafc3dbe4044b87111bc003a64c8cf9819899;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19eb5db324a1339b8ce9ce295d6c97195fa86cf0f08a7daa4cade42de07fec288776619eb3839dbff5496730ab77d7875cf8413ff7deaeeb8f88bd692ae232bb8878af1ad68bf1ef0243ab9fc5a0877a31170d1d91b3014075b0d05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f82859e8bdda703332c4500ec4480f5f2e48628be1b3a3806f15a0d8d1a797542be13e54b52c1f638c138ef9ccc65fa7852006d9172cacd25c163a1b6d7104b66fe549985c8ce1c31f65f57cfe3c86461bbf5db4b61b9bd107f56;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146c0ba90cef1bfcd135cf85ff57e76d98fb657a6c84dbfe5c998d0d0b5e8011b16e774080966eb1ebd4e2dd6f7f239b0d7d08e4f3b3b5c47625368e8b464fedca04c39575e7dd4de27bcd9bdb4f57ee9d02ef5f0855ab49fc96356;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9781c8b18c7e7cefcbfde4501add9b2dc5af9fc37f9498639d7298a8af16ac170ef2783d7e437617c7c9644a59b922cef382d995aed150c3a8296dca8133215f9427f9a482d2b895370ba64b58003d17b8eb3ed569b8fa28ee8459;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95c05305f6d546a31633ddea3787da603da57d87519d8e224c1ff81f05e70022422f8bca40cc193fd9a608f875f97bb6a66087d39b9f2c723784b7aaca8afbc58429ca6f847097b00b1a490c9fae9b93d59f80949af0e548aac9d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h145350e2cbcb2a06a396cc3a3521f4f794884ad180b15d5abe46cabb0e5cd709bbd26cb7af9574761e2d00dd23580d99c3c5f6bd127ca06871df20a7ba21b1579148a3076901908daa6439b55776aceadc62b2d51f23cc95071a1b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fd12e7aa0cc3b39f4c6cde96ef1604d5df26a1c338a928d6da0c4b485eafff89ba8e133b2a2a409223cb6b940e0d7327c56df92932d8e40ac29deb2d99a9a557f3f06bb9ff6b0b24cee7f988465041e648611a34cfd21ce07feb1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h147a3e834d636d7ca958ccf4fa139347d2d0b9b449d7d974fc2844f4d4544de966201af69d580fb8caaced4c4201f4c6fce973b03775d111ad677bf2a86c3e8edab15ec5b35667bfc95f14e4d2132bb7df02fe3f95d5e33a793df43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ef5afeef2eeb70d3cfcba1fdd0bae67e013109df325b3d76536ca07d98d3e52d506558dce8bce7e2f32cb2a00c376a8b890a623d83b6788d8c1457b578f030acdba7bd9b11946f0abf85870a1bb680a167b971f40e7c40c0dc49b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185beb428b9f8260020780a199cd682568c20ab71b78edb71c627945466eb3efed5fdf37494df982b0f17da2f76760aa0eac6a0a03ee5fd761c7bc7b40c7a07352aa4576b2cb2448fd5fe716dc35a8f4f37a5bc253c1d5ddca97ba2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dda2115de6021caee0d85d05b1d48f90ff6fcd1ed6b3941100e408acd2e9805a50f19763de540d449dd34200ad27c1dafb398e318f1c83881149aac604b0810834b404649274dc2cbf96e04954d87a8e797774616f332c2d62a27a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62f486f2a819b04aca1928c50bd8fa777dd9abc7d2d90a311395e8ee48841f2950be4a4f276cdf4c316f5afcaf162816b7915c55e7802ed798d3f4c2861582f9dcba6609fb9ed75d13e15dd04ad367d4b7957795f10b0464247e40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b26fb809a1edaea209a13eeee0e130c31feea1d223d639d5841859a8b3d1cd6fa84afe337cc1c418154c4b8e7eec28b32c75e3995b09e85628ab7a55b6843ba733437d2bdb3e5830f98097cca058959365277ac4d79f71fce96ed5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d49e43c326d913ea8f9c11e39d407e4aa9276f030ab2e85fbb72d62b27a40d44d4555c5606bca7232d8c74dc8d55fc7b8d7fa704b77204ec420cac4d65a9253cee45462d71c7bc281d82e3387bc82344f51123c73c941dfb2da376;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da374e2cb179495bf9bf2cd3cb86b34181ebee4fc6284a7d5446c9bfeced730efa4825ce0238c244d48e706bb439fe702f4b0ac59bde4160506da4079643d43f51886a0b965d6f6c365c84dd785634a952b09fd9a5213777b66172;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbd5416e4d378a28869aff69fd30446ad5c707749da6f4276b92c301148f60a0f3f826419875659b57bc8dc0e1484df955d688453b3987647e22458b308d9be3560467c639f2c5a3d787b6f1adef595295141230ad7c68ef495873;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174c21327f4d342749f91999ee791c4b78b313210841efdbcb619c84158803524ac080d28c3267341969aeb5bc96eab9eb7c656e1c08d09e2e8a34879526495c27c149f77265e4026ecbcdcf3a7432e8335cf4101cfa1a0e1b33076;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d56faa37b04c425c6edc2eb9b9fda94d084f088c55dcea61c257ac5fcad099d15e706416d0c1f750ba27370eef07bea278e1d5cf5e6792e7c23ce09cadc668aaddcd260a7854f8432592f76f13fc30ac8d118f4111cd152e923647;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3433ce0658b242ce817248e51801a59bbb9da6f4efcd374e8eafb751759fc98f1825872ea928e4de220ffec44880fdb12cae68baf44c7409fcf278badcc85ad86a02e1fa40ff7fb509a8116e4a2e16d8638bf99c602308a3f9c3a7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c559bb280177c769308f88ce3bdc1a722161d7e21eeb7fcd71c3c409394d91e6f3a0906e90e63ed038860b71efd53d2f7efa2fa385b5e6815f2c077e7d2ea9001c70b825a2afa9241286978bbc0824ab1b965c123a29360c52473a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7a392e791f73afb636b0ab5582496d9473fb89ad395448d03aae6faad1bf5f01e2da46532fcc203ba33a0e42b3283b1e7ad76697f8435f2eff22142d7b1dc04e06bb4b0147bce3050be13c55c692c6c3eaa155e57ba110ea311e6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc96bae7e96df7471493066237785253fb865b083b90bbffb66da4e8d27358a57a4a8277473b6dc0dcd83b3e5a01fd7783d0bf2882dc52f61bc21eed435e4cd0f64037f6cf5804eabd90311e6328ffa15317e36ad3ba85771c4c2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78c3c08b7422e6d707916da788ac4a2a002b0a1a8a81cdb8f1eeba599e859989a5d0ad6b7b6b3ec1393cbdecb61a27b8bb363a9298173f3e5aa59ef49fbe909e5539bebe94b32b80f95388162adf29e72b73bd160a47ac3e753d09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b627ba7b4283c0c496b905c67ce863e08cc26d38ad963df69d8144464b7bfad045d20cf5dea86dcb0d3933174cabdf7dce6f53b8fd4afc28317ead66a6108d416b4c4e981d55bf1f3aa608e439df77a7bf45ab4c06a667eefbe0b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c6911172e02aa21d5bda5b1a3893a9d43a0c1e72ba7060ac4bc37e0ee8d6f9ecf6839b9853e05439316597861abee3be826b6c91b8f3bda00a45351e7078a51e2ca5160076dcfa8116958ac495b22135f00c54fbcf0472adcab6b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1407c729a3993ea02466eccf0de86648f913163518103e2f45dc8e10c1d2f8834a6c62aecafbbdf6d9802dae92d83837c4016cd9797e2d87b99d8bf8efcf33c4e90567126a33accef0f53167c668d9fbff978267d5481874ccb582a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6943ddce39e7b3c6d1415ef28db922738bbdee3b30f503dfe0c92e5f12ae8511a460f964c346ed7cc466830bfb97f05881353e5da65c8a0421f45ecdab3ea4e2d12eca5ff98719e5fe9c4962ce1791d7a9dcfeece293249fac5b2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b91ed25d31627f8b902b06a2e79b24b224a87cd21169dfb9f7a18b714b5c42b1ac88f922e1fbfb0851cca0ae1c7bc9c408945180377bc79eefc12f94ab73116a3c45c12a03249618198da9633779ca7e7d59a9d6215bab3a975511;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h311a73c9959c53f06c01ec1235a20ebe66b3255ef9f256d40bd1a7de5c9675fc4453d59ce847bcea96b7d256837937a1770f652de9df9852439bc51a9a51f784337111cb2925be2efcd5ad9ac2e6b4762f6fc379a9e55eb021ee4f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ac3af91ec6108d48c656c64b860c3a4aee24fcd6cb0025891c60cba9abbf925bedbdd53ca7856f0aa2c0afa3cc0d6f8786b46a8f309b6acdacb7edd10108c4072f06a7b442642ce1a514c55b0957399a34e3cdddf66aeb68dc6ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4986e2209270888cb8d25e8e6f5849d8d433665f09d2e302bcecee266ffda2d633cf875fb1f44f8f613ab119136f329f38d39aac8000bdfcc04d8f60cb51fa691c84493bb7a754f976bb684a569ddc28872a2b8a1dd37638ee190e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1019a4700d72051bcebc30601f6f862b128a1ded659815596132a44d9256ad278977316fd6371058f591950cfa3696de8070f74bcabf6fdb8a8cf079460d99371e51d9d904e206977d024db92d17c9d7c5d67a386860aa383f3b24c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e51ede7d1ff0915548d56a6b0d132a353d67332d291b488ca49f27f92acea15f21d9f0c3ebbb50a9f9969af40dc5b81779aa9878cb649809d19495b1d196056d52164a07a3a588a64aa49426119ce3f67995b2cb94e2f93a9d5d27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10361bfe6d0137827c993583078f637fc03004d58d8eb67ff6b7cca8c25cd87d7b4655501f68c4adba110634523a9e70bebd699988133e367732e3a1ed88566a5105541f0bc11ded0069775856d9fc0fb031927bbe6da7e00fe3c25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1625a27547a109e02c8a2ec4ac78107404dd74c595a33f1b039e400720666e6093d37572763f2c3e114ec1c974c35aa0e8a6bb4819d3c1fa4f991ff13ec3d96922cf18b6fdb72f14e3a67f0e87cc2223765c32155e05349bbf3c212;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8673fd903286a39f7b4800f28adfd99c80f63f4c63fb23415325c2e84e6632944de2f2ef64da6de808c29e46517f9acd97719d3ce6c79f45e9586f855a2279271b906501b092666d80bf157d9c028ba172696884780be95b6fda77;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2e0a9e431038e721e4dcdbda2a67fd08d086d35b4a71f21bcad7e92c636f41f65ed7e397b6c27ad1f66642b81af2973453c789e52f57fabd758861c5abb6817fc7c66cf3ba5656ebaf02215ef70ce566ece8d2fd00c62f8984038;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7f26113d72b742c7afd9277b07c242caccfcc6689dffbcb4c47199435daa4a16707e3a75839793cf7da47c37e37ec7697e6b699ff2ee9ed3ca1ea39bd8a3b8371591e990ab891d4ed0ffe7cc90e1d257e8c9c4d13cbbff7ee04ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h636981e00a658a8164c1d8458f5b655a7faa673c2bb5e15610ca54022a27570e2c6c164f16f4bb22b6d54761caff25036248571028b6276786f1fadfd703ee2b086b2fa1948d3ee5f89224a7f8878257480d6afe8879a2f3f78547;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6372435527e59882f07e35bb6b17174d7c312cb4fcce4311a92b9c94117f5e44c0732ac8c56ca9d2428470a6db6c2a93770298608bbe3e24fcffcf6afc4de60264fbaf04ecf7fcf03fab410070fa5c69fa04f9ab0ace4698895063;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49ec66db1f59e55de31d259cd21bc80afdcb2fd82cfda7f2bb0ca2be1a326ff886b5854890fcac60d35cd7ae7ad001a446b64fbe80f50224559c2843d9253dac5401c5de6528b28391854f882323e9ba3c5968afdfb1e71ae97de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e03f3a6e8d1c91e060190a0711cc5cfa66d22f96461b54281aadfa6d0752afe1b16ca0edf01d3c1fc000250ec44582a66205feb633d32cfb4b53dadc69994da62de5b0f12afb76bbeee4c5e83db2f925b5347431441f8dc95d9b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6da6cd26a05943cb0da6c18203a2c3cb00287e3ff5fa940968c8ab1057d053e39ea5f6907d58efcd07c868be63055e4cdbf94cfe2c4c716eaf4b7679c5469d108e541cec08ff2048e8dea38403c5fc08e6127b9b7152c04c1254b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h408561dd4436bd3c695834caa521acc93c0977d3b656f0c156e760e4f03cba4bc19620af5730985b14aa0138895a38bfcfe5ae013dff6975ace23931b63aa46d0bd55dfb73f58629068cd52060aef891c850f9ede29aabd4a81c70;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10908c3d61fd3a0cd47c01d08bd258524392fe8c193ddae80ac6a946932dd9bb480aa45e0de6baf8e362f1f45d6c849c234806448676991171b372b542989cb300a80c3ffc2b83601859dc596a7c951a19b703de65cf45469c6093e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c4525ead2af3555c41adc27800527b143f8c3a204f67ca72e9a28fcb9ea0a3f35f2ef15651651029df5db69d3e73f0b5975da75a942b12a7d55abff061268ccf75022de7b1970563a38febc0d3312a7ecb282968cedd5e981e701;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140caa705f14450fde03cb046584215d9728bc0094b09f56c03c19694ae53c882fe9a443c289bb66f9d97dff3ada233605c4a0447997aa1ff916041f6ae6dadce52551574b445b07a065ef901c448797172cce0f1df749635c2acde;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e5a5937741adab7163fb3114f694293d60f26cc525c7e07720ef66a6c368e0a662124f0b242bae46f1ec9797f4afb85067599445681c4c0e35194f20c53310eeb727578c1604bbb5fadd1f73c7b1466b5c9f746b60a1ba463d552;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e48b7644ce1b70bbf02c738e378ed82adf22703f15182066bbdd4e05c2f0c7ab047ac8b1c9f0f08273b4e3bc6208fb1d6a2d649a96c86467d1cb708ede95c1592fe9767867928fa74d820ca9a7ec8e9b4852715b3c1d232184acc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15132fc0e34b44a294a0de3de73c640105b0b85097d7b8ae0f4d6bd810f39af4d2c252d5874d5298bd94cdb750e586d153dcbb411964a9d83278958c212d1b61247a365fc49e8dff558cba04f7c7b54087f4b34354b5aa558b591ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb40303cd4f6bf9fb2e7c7dee678a575b6faf0090d3d9a89fc7ee03ee4344f0175374cd1642942a3f1ebac36b87edbc3cef22788e66bcb467d6fb85155b5f753bc37c69019691afad12eb91b4593e03315d9d4bcb2d86f2953d4b7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1da53f2d06ff0255ad0788c46f5c55e6ae2919ac72406520f942eb576845e857ec64f974899e0c7582f95ae17d9c1ba9d203a7cae5da362fce7282c3ab60ec025f3f159304a957a16a1ee775cfcb42ef98ae9b184105d6b372f60b9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab2ec4d50941958adcb4b675a67805ca8325bfb75d39845cb0afbc0f037e067005a7b6d00dfa527b22805d37c46e2e5eb83ebeb3c6224bf591b6d932bd832aed05c66c3703a270ef7d474d2b034c8856ee13fc3feb5a9edce0549a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd22b90b203b9f206af3571f0670af34d494714bbb8113d8f9a2ea9cb6ab0356b30ad48843c4d2bcc1a67b7e142aaca0e5b455b551338d685ce1cd1a56024368848782ccef2b8fe0bd2cbcde7daf84964cd21382524343858ac2637;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8fa00a077c1df28201cc9b9f7e7ed9c8935eda2b908c52dbd94b5b53d404a1ecb995a4da4b5c2ede6dd50a1c42dea0c4003f12ae5689763caf687d53b96ed643b0a01aee3289f96bbb8e56d0b4c2fbe6813d17b07dfb79d3b899a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d3981926e4dd25ad94f1000dcf1c59261fb4e6e60330e164b76b63d9caa7a7fb53e03db941ddee3ce5e50077cf4e660b4ba01af1816ae2764a4239509cb52a8c7a3e93d3c52646fbbee9608a7d90c98f8da42bd2bab4cf9b54afc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2a78c02030bf677316ee29c6e7a3cb24bb7d6773a749b8ea0432a335a73101b07c955d96589659e60ebf53b3aadd96d5a6004eaf0dc56345cb2dc7fa527c3d898a9d5c90ed55490a6971211dd9f71c82ccb92ed78be9c184bc9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cd45f5e1e1cbfae2cd45fe5182316d775f5d303554fdab6044011db198169af9692fadccd7c6c45adba4b1d2c4f674fe79e033b9c87dc17c6de4a7682d18a2e8c796ad2568171ff61da1fc0639bb0174caae84554348b655cf338b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2fb52d3fa1cc6259d47d4adc1b263c4d2b56343027cbdddc7f3718b07950f7de6e3b63d121c42c0909438ded33831cbf59a9ce449ed686134d038e446eac45bbb2fed69156ccbf202d56ab057445e29ab23f10a46711b11c7a0081;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93bbf510680a1b8e56aadb5965a07be2eae1f7a828f9ec6f144ab3e90417f620eb6ccb3caf3b459abb5aceac40a36dcbed82826a14deff138f24cc5eadfdaf63a8bd8d2a693f4c1464df57d294a17cb964daf32fe8bda7312196fb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13950239bee10521c1d91e3081637ccfbd5b4bdceb35cb7a81c7f1cb8a2b686a5d078dcac61e603e78cd450a3ebd861818ea14819b7fbe5c5206e7596b62f461c292304f1be4182b639f5b853c4d5084c8d2176007b2c02749b19b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h982123fb2ede86a2a1aae00600b511a1a089ea17767fca446da15463ff753ee01f0fc4308384680afeaa6b6b3aff43bff8371e09484d72067a12ee654e4738ce8f32f76694905bbe3d84c1089237cc4804767d53ded9c725d10d98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4636f735550c78525eaede4c01fa6e4e8cc7f94f6ed468b005d28bf71af57be49f0711df8fc0e40bcaaa23565a60e42fb97b96c32ff170a58f531147f6955af149be07b2730cc9d4c9702ae181eaa2fb4586e1bbef5e51228b394;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4569662770f191d8efdb74c9edde5e308062e5068afef79d74c56e8dc0309ca5a23e637847979c0f2b7e9a9a239b5a8c909bf347fa08b403a81349cd2e21283ffcfcd923d1de0af1a8de607d9e0f346c14d41d89988cfc0669747;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2860673a942c56e4d0b62d667287502878ca9b16250e07cb2abbdd17a14c0df58af2fa1421231925b27d5218e77eeb9255fe6874e61aac0fe16b8724fc30500fd82beab433e7a05cff26b3b6f88ce7b7ab92b92f996584c21304d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105a5763a47344aea7465d0fb0a2d635092589877a448f4fadfdf0c5e1c371aec35faef7e516c2ec285291e418b984c7a0619a6999337337a1183dd10d34496d457fd342a4a7fedaf33344e6fd21d35519650322c58af92d1616291;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3f10347f0374073d1b8ff356f1039234a53e4a2db671d8dbf20d00664ffff40d43e82e38d57688ed9e5b522328307c1b4a3897bde79a299d920469556578bacd1db03fec9bc24bd64384d02aaea790beb76ce1127a6f9bd3b4031;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43c7715b800166c6bb07d61d623fbbf5ae3bbc991880f94373a893dee116b1874ffb13e284a7a2dcb4d1590c1d5da8fb49bfa44246c922481dd6a1260b59968c004b09bec7e1219d1ccf66cfa31c7ef2f51342e308d499ba645688;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a5cc814d3d06b3a6592c145ea74364413255ea5472d969c1a44c210c0221d027f57a75800d88ec7b434a798c307476da0bdcf517efd197ecc2332e0ec04e4fb7d95448241641320d1569d20e79ee76b3f6d9b7d4ba5c438171e39;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa71a8fc7aca945074119885f0b31c188f82e13490e7d6cceef0bd1194382f2cc003ebfca205a2477b7ed79c81e7b1640423e48281294ace8f0f2bff89ecd6cd97372bc37f25cb9b8ca714e7bdabc5d8aab1bb78e9c830bbf8b992;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f634ad646856b41b43072918da890f811f54a3759ea1a866c8f4d7710bee680858c9efe516321ad11a3f31d8fbcf96cd9f3fe5c7757b6900048658700b3f93b80c541f8694f2a4b288665f60dc9c44da62549a7bd13bb3b24de1cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b36dbe1d086053021cc8243ac6c611629e0853cdc7a9511d1c8e0edba2aa181d87b7a81408c832236255b75d7ed80e7e87cecd3a597444365dea827f2b69092e2a300fa3d8d81864f5014de0ef2a007599995009c0e23305566582;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13495e63e590fb6de7691d88edbbf4af3d62d55cc4e87a6289ff38d1ed9df4d2c1d74c51f14b9cec66346654ce48202aeaf74759a6e4ea1743f7972fd669fca837e82d1bd3340e8ab81c5b715e24edbb726d66b55dddd8c3568299;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h522604ef033beba1c5527c43b87a92ba64a817f9862a6f487966fa87d2daf7271fcdc44ee22fc603f888f41d46e19647e95685b7848f46295a2b54ce1aec13a03b75ae3aec06cd3d8c20225b5ddbd41971434a675dde2a889f2dd4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c5e3bf3eb663cd82e9616408fa9b905c2092a7b2c0afe7ca42721aadd7feb325c391770928463668f49cadf327fb1a0f4c438dcf79aef7cdf4284bc9f95e7daef1067b801fbcf80a96aba8923615124edc435a12eb744cbf92a21;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1a4ffd9a91aa281b57ea40fcb26cd5e29cefea05ecb0dacba930d36f78a18db4e2b14205be78de3988450511d94b41e60abaa0743a64e80a843c7873620e8424b73541da6ea2981c9e67ad33d9341dc828f233b8ee35f23b0f2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d41360b1d7ee897f2868502d7fae3910dbe6703e16e2d9f39171986cfb89ba47345886a6dfc1ead9d34203b06be5a026fada0c9e54bde213d8b4c24d54421d0182af9a2f2d4d14e9a78f878c2266ef25c5e6d08e2588311a43ea35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf208cc110729d4cfc395702a4046b4ad5ccdad9312dc217dc5f2a4af146dfff8872e7d363f54f4393b54ca08da6c7e5412d02d0427bf5af3a1e8f77ec78ca26d74763f4c160b015dfdfd25114437134972f7fa4815791a649cbd32;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6bc366a39122adee107ce8f2e62f6de845d78fa86cdd56650dc08bc153932f136f76c4d003f75bb1a21bc50037523daf9226976a05e4f6a3dee6bf5d761e50dfb5f879f4e9799aa834951214d8e4ee1730c16df8536f7855542644;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e0781d8c54d0d32df65d6060b362bb8cf053170398c6d7eabac288ca3934ed412ccb102292764f5402c20d95bf0b1ce1135437700ce1f6f62854f0257fb6a062ed1ab1f7a4fc595f093ee56e23a723adba2f0742c882d3610a48;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7a6e2072010043ced60d3313aa8f186b2421e7f40911389e441484f7abe54757b357b526802f6217cc2161b6d13ae98df5337e0e8b44b90802843d9bb216077d2f5b9298e500d21659e6f0d86909029dc998201a0ba5a3994f6df;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6773cf484b4626d5f688736acac05a21d8c71b8b5fb89c5fbb9ca1298144fd70b65a3d4010c577c2443f5e3c101fa747de97b055964ea30bc2db800f33980118ad0cede0719b40ba9d7acd11020f1ea28f787286a79b84ec0dc710;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha77c7df0447d37ee22ee709efa65323a783ce98f8e082f9fc397350b508a78d776567e80bdbedfa77b49d5f255c691b3ad1b6f9b2e728643d24f2c8be0e4547ef48f6fe611328f6c667b29e42f99e0b0295c092cfb64c60ebf6eb8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8e508a7a5e049edb32b3cdaca8c12aa6022b8fa3f90dc4cda7c6161f8f5c0ba101efedde20e3ac33b67bdc1be0a9c074771e493e76bd6465bbe72202c0282a6f550b666ccc677bdeeb0b20d2ace53731618f1d096ab43ab8e54cf8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c24c9e2405b7159e3a084687112a91de61e185ba3c4bd5f699bf89121dbfba4f57b6249739993681d7ce3ac40ccb1d7766393d81cea1e0ee355031a2405a61f0e1b33bc2c074e66faa167bc0c39f61f9707ac429632b4ec595960;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed198eaead3f2891a9db9352590fda21293135984124ad06a713d59b89d523392f10fa314ce147dc42f51cb8687620f398c5299b867dd46e116e03e6cf73b15e91656a7108456e40fc401e2c95325c00dca1219f06eed35725ee54;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b50e063753252bf64ec927d3bcf7947b3e3f7e160dcd3208ee2e0e91b608730fced7897c56fbccebc91145f26e18a5193f7ceaf5434bc74c5d25f81ec1e283e089f0bc0f672f5ed26d12ff4a0d1c4868a47c6a3a49b3c8e1c3e401;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d935bf8e7b9e7229691218f55255470e238e6245c1951624bdf76a42e6e452e3084efca944a1e9401e3cd3e663abc5b51b01fa32225c2f0981ee8613d28b88ce8f76747d995eca231967246ff0d9f13677ff2258f086c7e71d623a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8599563df1634201c88b971a05dbf06b54a68d9a9c84712197d3cebe62ecca0972ebda5ad1018ab153e8a85d26a76e765ac76b9d3105bd566c017f2ddaa57b1b644cc58614808ede1927fceb3c9a93f9e5b65710a5e1cebbb04d04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h977f4b6c639cf1417eb4056fd1d54b46ef8e88b76850dc58e2dcfaab4b354b1e5f94a875c581929f8159490bcc673b21eed04abde697d5bfb070fa806e44845816c104b220242b939d54167dafc7de2dcbbc107eed72705c561a52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3d63481dd45ad39e8a62d94877fdb4f5d1a5c81094f47de9d78bc2ad0446ec988e0232ed5f5617af898b6e3201295c71b8ac6039365df344e2bad88995f7d713cfe5d91584dd60921311c046fb09a91f1bf192ece9881c70686da;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f2598e2315501113f2df3d51a0c520a0672d4fce40cc3b4d95c1fb31463e5c2e902a9168e220aa412c5dda6fb0e17390197db23a28642af00e70ee50006f89809eda2b4bbf17fd719d643c52065e1fd8c4d23a8f62991f113ee4b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d1db953d173d7030046fd6f5f8ed9046c2c46f651368ea1c48633bb9c6d250eba0c57f693ccb1114621b62bd772c176d3cbcc3ea08a1af0595357dd29ac2b3a2f2ff944a74950c24e7dd44f49c7c5f41fd6cb5f1aea2d71c4b63fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h132f904e43e605ea28662f6e91801f1f67f3450fb8e2f74da6332055e71b16b03d04e0411d618bf7ef48ce20086bd6e4229215e36ced56fecdc4bc331a24a7b1ce8598168fadd2d340196ee6c16dc0daacc75e4562dd5de5edf84d2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180962f62b3281f1c0e4798fbe5b9cf9e7599eaf845e96a23552feeb2110bd899b3c3b49808e82a498f95dc08b61d6b46f94bf0c260fe466213198ad7b0a0c2557ede387ba5a6eb54395c1bd9b76be7b2874569c586215b905bbc7b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f3718e42416090ec162fc8ca8e522344d974528aacaf72af994772eb4e89fcf912d89dade851ebcb266ae668f988136e5c412898f4cf8f9cdda1d5d95fefce974c2fbe94dd2d0514d040996a2b69fadb8b44563b6d84d5e09f8f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e1e2db8fac0980807e58d9be31f251d8061fe9ffa91ef59fc3e9d0f2c5048ed7410dad9ebc04defc6b39c0ce6bd6ffd394fd6903db1c84da4096b01d5a124b3a05c063b362467c2848c1cdc89a5a3bc54f28873f4b520eebbb5d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11109b35b9a755d304c5a7478cde6683f3f073a64ef04329d4d4cd393a4f215e2411589e38103ea1261a7def271256aac7494340cc10ae03f81e88b489c1e31408b4ab28c1f896a72bbf1e352a40bfb8ef2eee4835e1baff3baf1c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1067d22d1948818200fabd62bd4ff943b403c4e6faf4bb6608f173b8b586a577a25f15a07b7a502123ce15aaf2e6cf1f03aa0b768dbf9dfeeee7a94ae1010e5d6fa1d690b90e62cc3f06fbbf05e9bb1b6ccbd7100b3b3a349c1de09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h558c34853426431dfa3b96b10b0374f77ca325835527391806ffd6793a6b861ad66fdac401bd78ac9e089af3c89a4d79e4db3cd90f1d2142438ec8acd4bea1367d0ce57c1f402bea44565798a3fdf53f51b9c34060d54743b8f0d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100d93a24e9d8dd9aac9d9108f9fdfae9afba2b20f01cf4f4c74a89daed50c9fc8e5a79792da7d700543e367d8ee792f2b70280ba1271b6c0c341ef221a2396b5dd040de06dd0044d13f45ae2e84a1c9999284cbf219d4218126663;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167bbf39476a60cebd4f54dd781c55ed24e8ae137693cec446d2748bbb6c7980d158964b492c6e2ec6cf5560221a31a114dbf8d80d16cd3d2ca5e8066c0bc8b44fb1ff47aed1464631a47fd41c6cb96df8662e02f0db29af18a6dcd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb81512b131dbab7dfc34ce0a76851530a242f51c0f608daa45e19409b72eee2b1d75e3da27b437a8229be2cb20dc76520431fcf0ec32e9a71c954fc8a8668f42311ebe6de2d89feb77e2ee74e00a337d24b8f0db89bc1e9eb2f6c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec590412c1f156486238e033851b9ea8f465a05ae8728cec6765f20755ce08ca07f9aaf8692d598ed30da0b790e5f4b6d9d8ced379c30130aa3b74a3530f68dbb541f345f4238dac50542479ce824ac6ff5e93d8b20827073a027b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1ccd6f27810e87fe5923e1660c44d9a768232e69a8ae0120b8458dc4ee61682307ee849d4562c7e496a12a706f83c5c59cec0e68229b5f0cfc5f5fbbdbad59266003a840d8e1136f3c0b27ff9a4e426c4de441ed70240d26c2c40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5e465c50a2b2e34642ed0b397b1a54c6ba2435e6dd1a66eb42fca601bd57cfadc1569cc975918ef16cb76844c05e1d5254e45c245e7158cb26bc5c59157b99612236762b205f1ecd12a3cd940c155c4938486cb429bc2abb25e08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131344685c575d3c37c14e48e25b4772604a691e2e9ce121fa854da9fa3d9a9953665b013fed4060bd62cff9e80cf0310af5853188c9422379b4791504ce9c06d6184ce3d1534855ccba3bd617d69e5bef461911b8caee7d814e0e2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83c4e48eb8cb0015a9bea3e1c162d2e3cdf340707a243d6ae10a3e6744a4be700f1b76ac2b58de68fd9bc2ebb17b60b3eb0b6a892b976a77d013d84a1efe6b26c481fdc0913d4769116af8589d5d038526b7a8041d9cfbc154603c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a236f33c856fc55f0d8a18d7cc9276407dc149fa3eeac535d833f92fc05e2e30660140e7d520c11608d45473621ade53d9fa4a58ee0af69c2ba70541dcace0628ae03290796da8237e22c6c85f3cfeee3b81a399df11e5ea4f8067;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172294a7ded0a26af8cdefee5c83f5f24bd722c305ad9b768f3e774e44ac2c63becda7c388192520a72e4c59461008ef9580e3b8d5d539df5080b0591338554bf13e876c588c1ca3a3629ebb0b23f1856120762deaf8eaa5f5d9445;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4851b465f61f51bec71ac116a77cf278fb6790926ac4efdedeaacd0c193237ec2c3ca2ad2b4085cece1761e6b83b4b7444516cb7c7abd325f08a5d0604b014c65a9d531d4daa7273c086cb9ff6a529b416acf979c42c34bdb6f83a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171f6591a2ecc9d6ffbb7b161b347ffeb0ec99195c395aebdbb58cd630e78b15921e14f00a408e2706e610b359635c5cfdc495081023005b1607d3f36ad20fc6af7434ce7f431294f1bb0a95aaaaf1067e8c89ca898623418aee92f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'habb8599becf560b275071cb65bc4036fec589fcc29f889b9660f92bdc999dbe0c1556619e94ade762c65c6c761cc45218a5aea12d7ed2e73122cb87423c41e9311a55b17e4453ff46fb1c4f5947218a7855f682a5a2902028e1412;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7a3f1ed620503f2c22786948ff28544bb3cdf4c487f065be755151f65e573b97d8d2751a466cb348af894c120d27ff04a21f517f9905b8881278f69bfcb39e6704a23d57d87dcc64c4d1fd4a2c91178aa7d07aa49f0845cc125a9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce422aae6d906a4f88acbfe41af21542dfd7dc6bf6d82781233c7a79a6cf4ac8b42b04593804b2ca838603af6668aa169630a7d96d8d5a36da5dc02bedc8714875c6b633206abf142dcb1a437edad7c754fb20255d9884169c64f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ddcba54243ffcd2003c34af8b6df70cd8e1e23f27556e63677b518cd6bdbd83807041ec6f7b8eaaf6e062075d47071221424e681cc08d4a728249a272082f418c808869d5a33bffafa906e6ca894d2e5b0f6e6319615f08d231a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50280717edbb7c0864cebe65f2d396379cc20ca15899a9595034b812b1b5f25083fcc7fe1dbe30d70b26cec5419c074b7d9b7a72dc160459db5268ffdf3f1bc3ce443564fd49071b7a1e79adc27b5a1612568eae7355c25304eded;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177dafdf4481e10ff4768d927e959f91afb7be1befa7787b58ff90b70544c5d7db63b4e3e57dfee1677dfe73a3c12fe91cb6ae9c428138b90ef23cbf1d0221e100bbf97655b4c8e75c732f6e7c284fb972c80cb5e37daac0ffab9ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7939b2f6551250f4c6cb4b36690de39305b44c8a9bf8c5fd74547c4bc133c4baad3baa1001aac42bee7a8704ad2196de4beafdbf366a0e453f85a75efefed98dfbff01334630f4364df7134eac0d6fb2bc205e79cc13220c1b69b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1e8824beaeb2834b8d8d0c527b6d415dde12f232e9664c61b40f63d18763a79624f70b64ae13c390f60b1873d6d71617189f45fcfe2dea089195653a43f0cae5c863d0cb45e4f80671e6fc6d6e1f512e275e260ff5e9d4de72298;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad0bcb19ad51176222e61ce034a66244238b5d000eb69cc68619c9ac31fa0b28f212263c3526811652989581ffc155ab0b6014b53157729322a863426963d8e2e724bff740f4ab3d052e38942cfb53d1704a86a40cb0f6be5766ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188415a5f8ac84700160e2b172f96dfc0364662e0773374bcb0e10c8e275854c5724ad684ee21cde0efaaa8167f60609b8da1e9341d8ba386ac374c5f7c06b42383c81c69d0d0195cc23b85f3783ced975b022463cb6f2e0a3809f3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140ad7dc2d2b570b664cbd83b5f6f681df64e56d66ef974f3fc8269dc9d0ed5aed25a7c52994a04ba96ea0b68e7c9560353fb7f623c8a39c9a371e281f14aba805df8f8bd9e4b380703893bf8744eac3b1971b50f05e2801a40c2fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5db7e0c522acf18c4230594972f70c60ec0f7f702a229308ffe366b9bbf82685b4d865b7361baee7f07f6a7eb665da57fe9a5eb387709bcb08cab3c06f47cf37ee475f7b196303e0cc6befbcd7e80d4857525972b457b94e826cee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63ad1607b4cb7739c70ca6bc11fdbde2c7053415ca0d15fed3c8121b1eba026524895262681b3879204117d8620d1d8d24c7bc78de9fc640f75404d00766883696cb21bd6ab79e4876f8213718491a2a746a76e2681241a8ddcaeb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cce4a1bd3b46438277a3d6bc58e27a1d29503ccb853abcf31f05903c64ecb1e1b3e1afe656bfaed6ad6da12bacd32672002f849e32ddf286ef3715f622293d6115a75bda5d43795acbd8eda9b13b06c646c9ba92be430aadc8af2c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he10fd960d12b08d9226c9697413ae0b1c2f0496de7dcb3dc9906e199847e7da5a40a43c7ea277176a8c6e3fd0cadb011e13a0268421de696bcf672495537fff591a5d368291c98e194a34f7422fdcaef1eeeb7f6063131a654188b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h126122208420055edbe364e98e685a0201e7c417a8043eafaf441eaaf5280d34571418c2de8fec25d6ff633a5b723c3c4f5dc373b9a018897d2d7d81c22fe93353baddafb2648329ee129f7d8270e16d2394f552ff7bfd708cae2ef;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4a8242483edb4df67f161008ad00fa319da89c2f874f220d785276097f900d252c82e56d45c79ccc7a6b24137c4420a34f5a1e7e41983eda251bae6977349f2a8462362f346fbc35d8bf647147e1794553b5772189eadcc135736;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h477dcf68989168289d720ecd5e99b01b4fb95b4c330e6e9fd747635c825bdb258da46c54637fda68e72afe45026d9c023ed17627f8a71d13e03259b489aebd968c592ad78efaddfb239a63e103e533b11a0b90391d4fa3bde21004;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef748515572b92047173ad62d56d1cc1503de9c2aebb98b2467efb6e405fbe86627c01b6f259c201dc9e1e9ad7bb9bbd50dc1425f93755f46da8c54b74749d8dcb7327e1e52f9faefdc47f52cd714c65fdb22e95ba98cd5d3238a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89f9c79406091138e88e8bfd3e6e9537e12a4ae685bff1329d6bd3fde45ddad86fc0d698ad0de94a76b027bf408c8a328ec92b0ca5dd633885f4cc85d902b4d171a925d25527860c4f60a14df24262dbd036da822be711a899670;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d39004f20c301aaddf25b22b4e490f9382a68de1a7af9011dbaf1f47142b639d90abaaf5a3d5fe29a6ebd36e895dfaeb474ee53b9d9568153997a069fb93c78878df11814a9f1a039694f3e46a71119618bf95f5cbd172ca0f05e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b453c68eb5321e44b4617dc46e55660f40e9d13ca2f27cf1e0c72b6de0b05823d957e75d7a21f3c8c4d8bea6ed721751fab736c65992f8822bbc4033d290f75eceb029e26a657c62969e66f19ef9f36a01ac728775611c0a18179;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcc4a67f935c3d5e661cfe2a3e868c77a296c8d4980c8066d231fe89d0dd189b6e23dd3f41b228c01ef51750e10b02ceacb189778ebd6f6ece2fc4b533aad493654bd70e9475253a82f0f32efa3dd503d437b77ad5fab9bc73e19a2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b833c7aa5151632851a19d25ec88eda55d8657b1dfbf311ee3d8e10cb86354d08a0706aef99d346b4c29810a8b402a0fff2a9ec3e617c96b8c027d543a2866188ad6ff461b316873d2facc1def19e822efb15b16decabbcc61c037;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1548d1c9143c6de352765f19d7fab15cf038c517aa95d8b569a7e716f3cded2de2e00b199b40e172e8eb30a92365c827ea3a7331fe6fa778a1decd6d284daa1c6568bc274f97e0616fe897fcc4276e6b2646cd33771c440ba98d182;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2c4b5e16fc285cac89a1eb94966ea5a7fa6a320797071e085fbede9a86c27a8a6a4d83f43179a994a7bd461ff7539501c8d74d1d5c71583973405b16c2dd19665d473f989e0abda9638407fbc6616ea7fdaf0a12032b0444b720c8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbf15c5d98a6a9b3d7fb97145b27902f7d1191267e3e9fa1ed082b8d994102ab3d787a16fb29571c3f95e79d912769a4476b6f9602dd246e49146590d0bf98a78af9a1841ed3906b3b2404f955f7e8ba05af752a781e642b37adb8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c907924c1f98abea02abc87e2822193cc30ea54152008cc80be0e98d6261e780aab102cb2fcf9fd3f42db35232e255ea85e342096e310c3b141733f6563d61694ab3ff87979ebd2f7c7a095e273b230b21502c0d31c5421b12c71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f045c63e961be0ab72434cb436bf13dfc7c48d1d40db3dc2c77f30fcf602b0a1e9a9d89788986db82dcaa9aa51ba1b16c294ca79a16cfb3cc0e1f6eaac61cbe46c96402bf41486f2a76bf1bc44ee5a07c4838a0934d0d8dcbd6b5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4d872ce6d27e0e420245dd80213449a741173d74e3adb464595321098286f707ebf6258afb28dc438ef16f045c6c49add02f57117175c868990977c236bac216c8a77895a9b6a7d65f38f5778f183da1efd1b4267bce3ca15efbe9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163097ebf789445fecd13f8f1962fb82589f9a2c797cb70a1edc52fce9f39ee3fa74c458955083d71a6e69e2dee65ca281c2533d53088a32039da735799f02833d53925812119d15f57cb228638ea0d65e123351e119b5b7d62f8f0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20283f2094e5d64701dd047b2c3e81c4d1789df656f2c4a1a416245acc46ba92665814816ef8796fef37eeb691728263b46f789c7dda54731d0c63da78b01b470a2ae5a1314c50e13560072332c2094bed6630dd32ce3a9d9d7afb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4407525ce8a453df337ecd7e5d726444e32b1eab61fb9623a5003ac12bee99c8781b9e67abb1ccee8cd39432a0c5dc5b304b0d482160ca34ed144e03b9b6b59b241423c0d5221e0e880d156b4a1299f98f0745681359d261deff86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17160d03ce2c66f6e3d36636598bac942d85cacc3a62f891beb498fbd921cd05b7929896fcc601c71e1e9613e3804ff19316f42e296f3738e6ac65f0b7028fe4c0c7096ee4e6fe79b618a7653842dec885c360b1f2629772319ee01;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab7197bcf88eab2cdf75fbb48024231acf3afb6e5608078584b4042e807c55276e2f53918b062279bdc23c626742e7b3df3b7982023e97d73c1c02234dc7c152a8c93aba0ee7db5b075431e075a2cb7bd25eccd9798601fa9620e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd501c3ee24130ba1484fe0f2eaffcba2abc607758cfbe7d8d0fdc8e2e85672ceff824a523f398f330d4974a076e23dbfbf1a5412ef414522ddfd6dbc5f5e55861c0c673df06464c1806501f3ccd8e433d59a56ea0186e4d1ecc86;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c9ea70f506b875ce1ebf9670a1ac919d6f601c7ed2ff14c2be43d1ade3975731f925e316e8fa42d0f0b65fc045a568d4f309527e058cf33b712fc20f06819b1010a76d8d080edad4fe1ab7d99fb9e3ae19072f7e9315cfedead30;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164a31e6f9556ade608f1ea2d4e7d83eb328855965a6b2128e117278dd13c0e284ea91b0358edd83b698b784e8ca12ef6212ce4dc0f3215bd714ff2b26abff38001cfcafa8a441d72d4bb014b36f5ec16cc8cdbef98496243ac5d4d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0fde8b6dff418bf9b083981f11ac6fbc67c06af3608b4673b2ca1c50003c8abd7031db1e532a081bf5efeb018bf41be8f4e29c06eeffea816cc6079fc37c548f94d0d80a48b631f50599aed84bebd9509a97f4ceebe61eac8abe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h595e790946a98fa7f5e680751ab4418f3eedc174feeb5c4279ccc0c7dbc57d42121b46d4e647fe62c072f15bd76ffc7531b2957126ab0245b949a1c078dcf0625d570e18c29bbd1de19c7867ebf9c2686f8cb9775b0b9084abe8b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c73f67a148686dbb2d0d383779c7879471922a5aa622b76b438873af9e9b6c00eda946617318dd81303ef1d9e22f70c212b6d6a1a8b8ba4a370440c8058e39e47dbe1c27ebf552d142a1478be8b78bdb4baab349bb7d1963235a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c32dfbda3afff1009666756d6948bca8ea35e6ba6d2d4adf1236b2a37f05a9a4b248dfd321429ce51117a81fe9a2123b74efc9031d29008a1ad42143cb2fdc2dc9cf7ce71c1f23b4b4f980ea4d5549964ca8ee8661a25eb042ea1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd197d6b73d91aab0232228237c8dc4c18f2f8a28c108795b8d1ece31f510a35d48e10708cb66826e4fd489ea659cd43d600fb3e1dc21b3bbbddfe5d2298f5aa44962a8df985525414dbbf40421e12bbd6e4e597a4f952e53bd1846;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7a91a0984844f11b47fd8da71c0c6e913467f8230608b75f3f1adc14bf6ec37748e5e41faad8a9eb62a94efac48b1384f75bf29759e0d1c2a6775f42d89916f24c2881788dbea63b1739addb4d276dae0d42c63dd9357f96f31620;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac5ff230fdea663a69039a0394b674798f16178f2059d176f7a925dc9e741df06d7f8a4e38f4c847456a89e256e129a7485a2250da285967098e23f7109fd8005a44e61b60ae5fde04a2400f8d429c59fb9027d97268b5b0cc2786;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e325c50f9ad4c1c81215f750cb3aae9cc86a581beb8c791ebac6a613f486aa66d3213e397de3208fb8f8b324c3cca5e8a89dc7db4a28cfe417994ea2a9dc44ba5baba1dfb40ff729695207b3f4b777e1d0f7d415d552613e0f3f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c498b8e7dffff09e330df5296ae71644ad7c7bc1ac6aa4c3602a5395a102eab6d2b30eaf355f261ae34d1aa8ccc26ed0991d8e7190926331f7cd5544da898aaa25c510c07f0a2faa64797ee02016c5ef5079f26ae9cae175f03d98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbeda10c92c8848283fd62bc7c05588426a784b7938c2e483f169b99562a68858ee136ef0b77686c6a468e424cf26033652789a62a096678e09bf2f46d8cf8c0316f3c54d9197d359c14310aead53f9c75c951c641fa6d5997b39e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2f991db67d1a199c2c50a449954f072b64f192165aa092f5e9e1513af708e79040260f47b70494270b541d8ee44eae6140ad86a5bc5d7b45d150b070ce98cfbc770301808dae9edfd738106ceae7c67a1c49a03e6d54a2d75423;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aa7639d21bd6fe26b5038a4465ee4dd9c48aca45f8622cfa541d0af91548ade50930f2b37d32a5a9b7d9d9601a1b00b9d838951dc004ec3774e342b1ec66b954e751d543528a557f33d5f76e5d19e4866e9bebebf30eae051afbe4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h44ab0073c8cebf408d33bfa6f8c309f1b49bfe8a96f145a242a7fc7fd1e2e3aafed2c899c891e81daf7264ec22d80b2e90433f3a22e275ac50e7b47674aae773b932b8c951305c604ba6983a20cb4e3106fde43ba84e08f434b248;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127fcf42d276389d80cd6cdd871518ef2cda0a116e0490cff25774784b30d319c45bfeb0a84bbab54aa9fdadcf9550b7b684ace8946c19b21510231e4e3f2bcbe9910001cc22c3a9bce50651b30fca77469d237330633067dc3c49b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he38526dfacb1ddde615f35afba14188e6b5ce2c477d0e35b9348cb9709e186025bcf10f461e651b0fb02eb090ba806e7015b068e0abba9db96f5af0972bfc6d67dcc29cb148b21f548d77a4b1a611d66cb47f07e3b64c355dd01e4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h150996bb3f4bf24e892e75b32b85adbf3e561ff7af22120a53006a0f89b5236eb45f99ccd83fe1a8b02f995d61a9e71d0b66a76a455725883ff0f8530c44e66be77d2a0254bac182383fd5e1c4bbb1b1d79af2d3e953bf30da1ea7d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157eba4305d6eec68b30a98b0f90fff1779255dfe0989fbda477141f62b7cdfedf70fb0d19f79b51985a490bf6029e5d9b89b19e5196421e06d9beb9bbd81d0deb343fe06576359c08e48605f5062c1c21f6f7906c938e642e788f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11205424a2858c1a78dd1bd7c7c5b86c4ac0e57d96f2bcee7250cbb0381ccb3b471a9c1b5528a322574596facce35e1f6c67a41fea2927bef867860b736d220941791655443469c4f420c99f8c4ed51553a432b69142cb57bc9f078;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4aac4a0ffcf6e56f0b3579f87952b195817cbe791fdac15145a0e1b6e723437d68b42bf05c2564f350e73dc72ecae00268cd7946e1dc9059de8d496b95be253a5825f76faf994287a32a64426545789e2990a3db11e3598e31f06;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h795c382bc06a3fb51cbadf348c19fe8c7038484398eed12f962059f71c9d5574cbc038db19847bc17d240edcf08d29e7929f592ffee3b3c461b04e06f5952310430449fbbfd11481439c56e14c2596e0ff41c11b4fd98dba714759;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h192a06eeed005c47202ea61e9688bb31a8732397bfe62097211bd37e9d9b15c73317c39251c009d4962b48c3a12ba67c68325c23e06b20477459bd4c6943872b944a30527d7d258c2bd5829f9c1f674a306516678bd830c876a1cdd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce74e213daa7dfcac91450c7631a596aa74978351384203a236070c5fb8ad39d0093466a02190065aef28d9b0a3676cc2589389dfefe0d31b64773526c7c099702ae46e45305fb292129ab71dd3fb2439bae68467080a0187ffe54;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1097ac07e9774bb33b7162adeb9bd04c4446cee74d6f5f0f86add6150ed8d37c49e2fcf6d48b499f0dde88af9544bc9e7883c2df396599356a518371504b5d308574884e069c0c8a01b86da10dd3c66bff59a81ef2d09a51be0fbf4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86daecc7e78387aca8b28e10f5d44aff03824934eb47cf7ec8e75a927730e706dbb912a57b813dbf2aea4b21f0af8fb52b874c8f778f6b26ede5791c7c5737d8f99282c58b87e92753177ea86a977f0e89af718c360c958ebfcd0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a5ff2e9b05f57554545ee92bf745f7e08e8e7535692e7ecc396dcf43758c3b567fa90798600b9aca9f82cf7a3388a5426930e2877700602874052be0eb196211668a4375f3dce4ee8151748e5292564a1d3f214847acc8da0436c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he293224d6bc3454982e6b43830e211e8813e8afb774bb33c22cc2a0d4461f00fae849a9c5ea0569d1b9feae627c85598c8980b15a078b082b0aa4afb42f56af3087f8caace52931d28eb23874d48802265a7144612cb1ecd0bdbcd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1376d4b10452264513f980686c5099f82dcfbcac1ac6045778c5a7e8abf304113b7fdf8b1b310bef1e3c6a412093d55f6bfa80dfdd0da0b5d13f398bfcac1283b1a9c45416da3d27f4fc3704a9085d6651d924b9073f03884bfb1b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5924b11a108211d26f15193f17dfed1a94fd973b9aa3fe7beac0bd5402cafdcbc17b060df9fc07dbdea75b41d28f8b630880009365eb5623a34dedb797572a35b747ebc3351096b7c56cd1e4d356b0270be93735a12174e276d26;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1965dc01567064d29eae10741709a39e48bb8329c8382fbc39d06f563a406cd2e31143b92939fcf94fa7cfba3e3f3f88321cee8886d123d87d0a562251d712d0739630ee8ef5b7bc2ec3ae8881644dfd946cc3effff1f79c6f0af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156a98a32ae113d6e0b983aca32f456fa2e9c771b4fbc1c5f8db94fd81699526f070ae8f3dce8bc911018afba3fd3f468ceafc543f12559cdbc72248104fa7b5eb1149be030b713881cdee3659fcaaa6d17d4d66637c78ac54d88ec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14386157356d2d7b5e6c9fcc3cbbacb4093f0684f914d44696f3012900b20056ad5bb4bd58a9c5f08704f0a61bf361ae3c865a07174157e59a2ed8feb3767a99a7c694db2d62c90f54114b12233683e985497102ac240a1be5dc011;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c7552d0f38e62cb8644b4a066f27501e8e09ebbdadfa1460dbff875912bebade03be59a77ba92694b6ca4dd0abf180f7b47f14f374e568ed84dd36a0260c1e6e50bd1a42cbd8492f50b9743bc2f6c3d3b79a1a8134e25ac0ac84c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6accb5fe2539e5abe5f49f3bd7ecf71d07251374c0970e11e0a2daa211b70629c290064a10d8dd850a9e182e6732a7697c2bd374764f8816536289c0652fe550363c9878269b1f923fbdafd8eacd113f4c88431732959e85acc05;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10e9d15283dafa1cdb94eaa06957ed535d50513acf8246be7f8d36676a6fe2aa27144e698a351ce6ea7f118bb70d123a995da4eea448867bfbbc167f0918c168a949080a54181bbd13a308fa45c3290385e33e9a58997ed50dffda3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11bfa7fd0ba626f7f0b3842b7203e13e45628da19d51459b8e2bece3569181dca48b99df0679ac9105215c7228b937fe6a2effd3f3067d97ba97d6182961467e9690864d0c3170e87051bd5d9d0364fdd9c8e5cd2ea314d45f9c18b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197997ecfc881284990192cebf69cda27ae215b16f7f9a3a09ea6ea872d263a41f84ed4eeb1c129f23a15a1dfca7b5ec73160a951aa366c6de333dd74cb1bc4b0138e8c36bd88f65fdd818c1e5500dab3121f378c6cb8faf7368efd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10250bc57159c31b15fbc263e19fbe8ec87f85e28bb632dfa3e83c29075c3749d7d4ba82de87efd1ca6500966c3d77549a7581ba539cdd8b32aa3b73a2d4e79f1e6d734f94db895b87f218cefabf48f51152be6b963f411827dd42a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c76322cf03e44ae9246bb530699b904c13c65f33d606e7c5d4534e0c08549f8e4105b3ab3dc2d541c02042976f3aeedf0230cd6ae17010a18784ac099206f95a830d159c7cc3d5749b7f396cae1e6e081f958764e55a92d6d94336;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96edc0547024c0e98eb0eaeb29a4fa65aed2d28d58a1ac0d741deb0e2377c5535acc9a0df17c3767ace9a0e6bc91bbb9834d986272f4c3c2e90c31dc94d24003096431e5e6658019573f1ba3db1c002eb83889986c30e75b515074;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce90557c123b87d48cfb70a3e8b5b79194a27c95f68205dc5a4d906936266965d6784c0fd61cddbbbd7900ecd4f65e0b515c9aeafca52a25a372742a3df8f604a189da6f9a4675517b83d0614b42de6cadf35eaecf5483a34cca5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2ee1b7e0c58825b1a76e355c5febe360789b370ec05c4bd18efe6aa251d6d2b7faabae31b7f78b7613b2ebb4b634f5faf78547ea06209049d6c1d63cf43e82c131c3108ad9adcda792e7002aa4257315caf957e86ee14457b0a13;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b1b9132545792a48c6fa574fb2c94e0507e5de45eeddfdbdbb0c9939278f8cb26090e33f8ffaa793e42e271fc793c415b7b2c3d9e9581a025b88bf4be35aaa3f7300c09182d3e83c7871f41ed47ef450c20779d2d5138f7d6abea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d364251a83e836aa1bd2edc0234664f791724d9f3b8bde14e3af24b3b1bdf39552f60b41c0d6cf3cbfdfd7b4ba8c1cb834f0ef4e67d9d5a0214d02d0e96e67c6454decca4a8e5a7988abc7e3545082b773d652667a192183b734d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha06cdef76c861eaec9a0e89abb52993008d623cc272307866367ef81f9d1492d100f4551888f300857fd8f2ba0ede07509b932052ffc60fb59c2bfffdc1788104a375861c2aeb345f056aeb317072fc01a4cd8709969871e8a54d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1445b50d734b8aabff852d20f2090f0c313eb8af90cb4bc77c2000f6fae27caf0d7c7bbb4a54008016a6ff07fd71267149d06cdf68f583a3ad994c0a1e2994a693e1a7166af092573ca07e7412159f3c98a68bf07238ca3cf693420;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1daadc6b14deb17c1d2b68a2fba5a916fefe1398b3fa2a7195792595d9416ca9ec3931438662883a2d2203bd2b378a919491c888f2cbe7ac4784421c212d472c4215b888c3d9e9ee0b4acc8a7bdfdd7c462771d50cba96fc9273bcc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72f96e3126a499c4ad2ebbcbb9ab676cfd772101a146be50385289880e16815f516ca78f8d1a33ab39126d8f0d5abf4c2bb2075243b47e323605af07112e8f3f8ab84b66aba701595c5e4285cca72792f233851f56f136947a09fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2bfb3cb7244a17043be7aab7c740501c45635edc1c2ced991a4ac44a370aeaaefe6c8e7764997910450fa0b9750086f9e0c26ec362e38d1bd17ef5c17b2050e597ac95648af746ecbf760be8e21822d206b4fea42f8f18b231e05d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140627fce4a92faeb331edbcd26e190d0c064c80bb0c5c84c389ed9f638d68e230d5dd8bbcd66c4da9768bd91b15f1c33e2a5a9f2eaf74dc84509db87ca112883fa1a2547c89bd47798e2314e046d2ea1883194dc6ae55de8500c9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0bce5be8496a4ff2d04fbf6b6825404f0025d74e3bc0d6fc459181b548fe4c3673954d4ad36d4addab1b96e31a50d60eaa71f2ee82d01c656f63111eb2e80b147fc557dcf6f937dded542ff6c6ce8df25c8610ba93bfae082aa30;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110c73a5804028a59a1fafc9e35157af721b3b2d60ff2292392290b6edd3ddb0d4b619fff9497c27178011ef750d6bd313a50fe933269c5035eac6410cd0afc55ce525d5880f5044335451b490a1f1b25d33916966268703bf7194a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14421ba15117b799d38b7639e27d15c68ccb0ceb87ab36657b22261f5c7d7ea47a5ba4ec200192fe6a50f0c476bf3ab4291b4de7a4be7e798d9462259e9fb5ca2393b7bea739c04d650dde935ac7a99d16e3b698ebdbf7c5237e4bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113f6eed2de8bf9024e311ee646ded7dc6cecbed9fef72c04f61995ff26e72435e7970757a2d84dbcdfed6ab2a281cab3380d97ce93ae57d761fd6c28a0856416c822ede449d20d3e3b59756c9e7ccc8dad8b051d834075508120eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcbbe379cb7119f4f868a51d67f17914161224f591f1a779f386481b84061b3e6ee215301bb23951de57fe0524b094f37d512432654c3baedac17919a06ec2e71c5264178f0d0553596de0f2a5224006d1914710eb71598aec60622;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9239f4ddbfab9a118f16838bb857b1a5cbda034a7764c635f4a05ce119cdf16e96fd5d709f2ea2946373e493d9116c221f08803597c2ed5be062cce842ed43c4575a6f27a5efdf8dbbb383e8cfdfeac1453d3385c037c16d570fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35ab2ff76ad132bd1cc9421399e325e6fd7fa0ec1983883a010204da525851e13c81536452dce4ee0c08eb9ca0bb76adc7326e0733cd59c9cdca678a51c19ae84b63fb28f7f535e06485085a83ceb9a793239991313eeefb9ba536;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h135272d64c28db7d5db53bff372fc64b0259d560a33818878979d01e6f366f5dc521ddd827e5c8454703e963266aa7c39b5c864cb355fb0046d5d0c98bf6a800e3cc431e1a96bcbf6e55b118a7d0466f3a070af0e3ac086533acb35;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hddfa5cea09094b0fe0260764273a23992207fdaad78e638a4132df65510e915e8498f6281e212b47860734089a0e0d92b3fa346ef12557b1d01d7a7b8ea1521207ce1bf9101b85ca42b63380bcf5e0e95e507a31231c4ceaff8529;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104a05968db976b8f7f4e387bd0479cbc2a07f7d72de56c9587f43d13a60133cc9d3a90a3eaecf7040d22042be9c5c34ac2661486b6c3863d7987c335525d234f078adcae4ee1757cbed7c2158841f5d65feb353a2654d2efbb2a09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfcfb1be706cf384ba0971da6a894167b6d2a1067837384eca8cd7afa4783604ce3b8eab594cf33d2ac49eb811ad9c56474be10a94d8afa970ba91d521f7945167bca274e2ad18306976b35ca9db65fdad53b9a48bc775f38ca955;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ac90de432f91a426e602e50debb798d103ff94147a3ecd5a7cc7aaca9b09b0887a5c8f541f97b122bd97b202b9eb6396238782eb88194c71d7aa86eee01adcbf535ea3a2e5dc88a1a79ec2c1c5eda6a76efc340045c35cd15869a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he52714ea83f8f9718a94ec6f16ed87529140428688c0c141bff48f490971f99f53b9641e49f9c66787b915aee32034de3be60cd49ff2677bf593e43f50e6889513dd3d1ad2575482a1bf57d560025c9d6f6e602aec26d3feb84530;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1adfc9504c5bcdc2538f10d4aae1147eaaf85698e15dde0c2306cc9e97d69984010fa521aa7a049efa1e8138f00edbdfeefbb47f50cdc29d7eb15f1b91f850f93c04e4d42854be52d0d095bbfe8287f2d7a9b6f4de5f9acb6e1a97b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ef52dca246d6fedc4c901c0e82244bf4f9ca1814eaa2908a48842eebc4848e5a3b7bd9547ff34bdfbb350b87597ec8fb5d7e02a0622cd83ffb58e6e70135970ebea8b044af1c63dc380fb2f7678ab137da1a37e943adedf89e42a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3e27c86e6549ebf9f261736bdaf213f518e3ef62c835560f619338c142832be02e3cfb38931d338b5df7ab14f446d33005812a369036124b6a229f1243ba25672c84d4b87cf278f071eb9ef838b8a40fcd7c8578e36b478435828;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf37c4a0d0acbcd36112f0468edd5748f234392d2f3a07526b389e51628df89656a33fc597712eb3e32aeb57a12f14a2fe87c5dff6521634853bb92b0e45ae11cd243304a38dbb0a69618c13d50db0319e4231ff9e9572af1d792b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e09ebb468cbeb80a043a895264b6894c3b1812c9a37e09b7e8ebc10e7511141b2f66a9e7b504ef0a13c81c5a2f7764fd640fa2644754919aeff2203079a7ddd5296e1e0916d5262e2fbf38527fc474d6af13f5606f17dd909ebe27;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1947806dd56ac33c5354f9b05a7fa352a862aa5204e533dff0e6591f013285291fa6825740521e1185db5d0eb0587a26f37010522fca8be0f5d7d31c712bcc9c41786212417b0292f7aa97dcc2bf28befaeabc836404f6f10d86123;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184bb0e4b335d016f007840b998290987eb390c1b7b77ed6b3f197da61090b4b75cd14338afeac7e15c0bed193b8258db90aa0c6970db90b439a0fa8aafaa54f42ed4d96b1aa2686f4d2f03d1716d24698d08471d47d40c3ec958ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha9046f648c349035fe02ce556cf5287519db1f59e5e5313943a92688d1b0085db680437c0935ae3f94fc36b58409c0f84bddd798539793704ba68db25d1b81ca1a299089c27396efbca6e9546587f51bca0644c1a94c51fb55bd65;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4a6c73074c46c39f233635d42615cc0d813e8acd50c9c9b13f0d65aec74518b7755ba7dcd4955755e1a3b692b80b62d35e31d0d96a4cd257e8c8f2c3700a72b574633c2769a2f4b7bb0d35cf279dd4f2c022ab6f961a4a9f6ce5f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be63a6c6c3e4ca90f1a5374dd1e90035d271184b9d1ec6f4ce759a680607a094b4ba01157c2112318fb6cc1236b22fb644e4f63d69623be7919a84b5e925b50f88456edf8a2aab3200e37bc1d67d3e28bd4a0410afefa367dee147;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c771e461d20feea4e3ec3268951cf690f374c864f887a3cf3002b24ff8e12247ba58ee226a3aa71352e0ece6a3769c88f4b154dccb25268114642fee51f78c68f09c865a1714ba9d49b2b9b05acbf05a21b6e9ea39ee23f5950196;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6f8d587ef6e3babd5559fac57f9ea9706b022111efebb7909296c22fd66d9f9fa00365c6589f34ecf13513e94cc35a05af9026e5df48018871ef23372785b8f70e26bec9f0d1eac0115bcedf0874b8d8ceed1207dfd89e7518071;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b58f0383489de371f051d10f806f569598501fb4a51ac4bb9203b7c3804906728cd9cd305b67ecd44f814a394b95f996c6b99e2bbdb8a32723df0e4583ec85397c3bba4c81d78c367dc8f981738e7d4339f562ccfb377c2b404dc5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15a6b1f5646f5dfe05a5f7ae738ae65a2588bdeb2f21e2a79f75e2e415c9631f54b4ad869ad4cdd96d15cf7547d976785c7d89fcbe5dc39286a33f7973499fff46039d29aac369e11249d928a56be1f2bf4c984fba6267fb220376a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3732eeab37e4cbd32e740e9d68f01b8a517eabdbaf63af1aa02743b802ef06f37553568c6b4c97b197852f30a5a253f9aaa987b3ac70b2ff8c9fb762356fbe130cb49e575750b0cd8bd3ba1bd2fb30415cc0b02ff2c91c44618384;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b8f0eb8cf7dde8777656bd1a01efadd9081a6f2f5824c676f0486005000c428dec355ab1996635088e99f6b1c0f6418a94ece6485d39d0771687d1955cb9fbabf7aba8c207a6bfda522d550f034da7b72dfaedd09f5f6eb6424c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168e0a49b5bc815fb99c09cf6655ebd7d2f3e620871172ffb7bf961e6608dc83cf0f9740f0ad4cd3bad570c2321861ef73ddf5e86ee50c7649ce22e76a4edf190391f919ffdb0d688db10a35f72eca592754010ec2e53f80eb8818;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8dad71952f1a0862ba4c4b365a86e92ae8b3188d1f25eeefe60aa475bc05a67d5600b27c1cab0f7d0de43be04dad8a03d22583b1add20ee64645b1ff320142b0efde4efbd9695479d09474f54321551321754ad6c4c9046c3c1ee;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d845e101e4d16ededc36ad0b353efb5229a1df507f317ac1d1a4363d8a3076da1e6f02d56b91a0c19a15327e883ec43f6d3b44751bf4a3e565cfbca48883f390b7a1dc2a1e0b4716f17a7ce470f201d97f4f761adcaacb4a7f922;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h818d71a4f044e234f4fb1333e30adeaeb2f3f2e2eb9a07d80e2fabc4118c73aa286d41b58faabb7086ec333cfa695208aeef67b2d659008aaca0ba2a99869ffb777e756accd3e220fb341ed266acbdd04a0fc040de9cfd940c62db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cae2cb0d3a279b65b31abfd91fb5ab9e4bb0dfef46e2f535ac1806c66fb7065396123db420d2b0c21b7e56b023901fe8188a2ad63895048f8210685a2e7f69a86a0b259af4649a92570a1eb9e1867cbe1da45ec593bb2ac67f532;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b63a0057af3f585ac5a3397adfb8de5a974470c4cea99f1c7b02022d1cf13f04ebdb67559e64b03407050a47ea8974f790b1cb8b664ae63ce895a978a1f5f6fe74928929cbbe973ebe15119bce874275f87f5e467e72b703c6df9d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cb9357e0a220a75b6ad09fc8fe6cd51658452088256646ab29182d5b95f9566564c6e8edc6868d770e29b0e9a8643e55a6d7231156dcf2e05fb9709e8e2bc1ae6a505d547462b7a41df81ec9a4556fcd71a4b81a78345bdb76cea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10bfe3d037797d0fabb75ff54100b64e42511e8040dbb43993391a32612e584dc613ef064573f6eb853a2972c57159d2b55b7b84190027a89de2bc65bef8221a9ad18a2624090f27f26aec9497ab1e038ff909ebdcd82e1e46cc24b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd66cb46d6e3a07578c876127d9ce0a910cb0409f831305dec2fc066a1d15acc8deae5c65ce9b09c071241efe94553c0a8f46bd55494253d390ac1630cc900321f25339bdb8e1679102cfaaaf40c9d3c528b84c76c709a1ba83636d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ded6cde141504c69e2d270ec6f3317270b650b6f08d7a422242db02b978848f8dffe53c5b4140e64bf63f5fa734c334aebabb4b1ea3c32fe0b6990d36a7a89dede4451ba1ef99cab2cf08c8fce87585a64e4e1aba2264485adc9bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he74cf11e6d7c66b76bd3b784c780873ceee8cfe7afc5d8c307c52451593f45f168cf00d2e9787a0eba37a1390d77e51c42a082ee8ffc88399d2c5b0a78e286d0df6a0a5e08b00b9be25252cefa614e205d9e718e09bee732783f9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h642e9900ab47b2372d224747fd481ca9b862b41e6ef760bfe8b2a40ac34c51b85d58d7a214a88cc9137aa21514173ef65143e90dca798282ea2ecf68468821c7b637a8dd7c87d50aa3a7e93c5ee5ebde6ec5b4dd279caf16ad7dd1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba846bce63afc3e66b7c62d23e6c2053b656ba4062449e9a28b2a38bdb45a8e917b75a03b3f6e16cf2127dbbd929203acb65fea371183b9ccd9b11c7ec5e75956bf176b793590e2f735f01928e6d5aed5ce0193461a2806521cb19;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155334a506b829636e74a954b71dedc68047d5d491e239f5634a4a804c7aa38d18d0db4a0d2a4a7b20162c354e41956f3dd57cedabe229fa828791fbea562766a9637c4c81fcb39ab962a0405ae5da6240b973b439f2231c175e8f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171c6e91bd446f2f8612eba7f6f37bd48f35f15eda7940bf3ff1fbf8b75165d4a5f40c6bd6e4010bccbd2be7eba1ecbaaf63fb26d66f09210aef93c4b30bca83e014fa32b56d31e9c9751ed9ad6ff4803b638cc2bf7283f8d1f4fad;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha82c1d13d839f14aa7288af56760c1941b87c24fbebc979f4970e74dd08900fa8dd94b4a1a864ccfcfb2104dbad64a1ea93c06c65eed3fc6f3c128d8734ddbf0c26c08ebfae3262c565f6679d14b15782372064c78d267865098fa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h44b218d26e5fd77d9f5e3c5248247e7b560d07b0e9cebe0a427b10b8bdaaf0b1b6c821c85c94b415937539b82556b2a2570a658e3978806f8f760f56f04adcf7b78d72f11de2e2058b32f9d3eaf56b1475de2c662a9e21b9db99c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36dec98bfc87738384b7ec7fad2f491a97b32e67f41138be5c170516ff559ce6cc155c3fc3ffa90cfd48972b4a28c4dd0d3d6cdf9004200b44fa8aec28024ad0f98d707c7d575c66e2328078fea782e9199fe1ff986aaba3e9c3ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8dc4b0ae40f23261837ce1703b42dd7f645ef98b5ea9499ac17ce97b3cbaf7545e19dbd366941c5492dae47a897551bd8557ff443982bb024a135f37253c1b687773eb178a87839f55b4a0af353499691a28f8ae22218ac7e2a69e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7c04d090e7e42053dca6581a100757b5b661a1ed656d41e27b6bf666d5023f05b4cd5d5ae27d74d1cb78724740e38e68fd5de742298d19373aefd295136631d7233a796485c83c15f5a0c35d63ef595037b6bb7e615f2ca08229f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h408ba8e6e60ed6c9fa6f0602d57e6925f2ff638ac6c0efa1535524799d0025d079fdca38b6dd9528509bdd0cefa9ab909d8d5629e1866add17adbc9382b3b87bd6fbebeb1d1367b99eaa190d9ee5bea951b354524bded646570ec6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fe3411f3476f312fa8f7b70750ae875b22a4223f2b74e1c2a0b0917f9d2f33573052ddcbd07fc258c9a379a7e85a128538b657c75c2c0d3c869bdb5d6a9fc51078873689e78be0c9126af1095cd6cc301da8aa32e69d43bd86af43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd97a47662fd2317b0307f664539127a8983e8f8c2fb012d06b12a7839751ebdb0ddfc8918f3e2dd871403e76d45e318801270da1a96dac1f337de842f59cfefa31f839e712ac112b59df08c402f74bb112e2846880308de5b5c43;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14be6cfd8d501e39ba2f3b603112eaf7fe582eca83dd5f8fe6db4411e6fc246e148c8f8fd14f8409ee7b4b684f3b8ad0bf01d4e308bb3b6ff5fb71922005acb8725c777cf669f0f305872382a7111fee43bc22a116ee12bedd4484e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d34239bc0cf6c1521ed02af73f999c59555bb102083f39297b38ac186d16cba7cc5c9255cb0b7365013cc5ac6fbbc7eda810804ade9c82a45f7dbb4945c355ef715605dcb1145e3e71149046cdb208ff5545230105b38836ec4b4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6bad66a6ad6a092ba245e860db48a4bd3d079fb50e565fd3deafc50c9e01fe43c2f626088a2cf3c84fc2e3d8ad79f331343324d8a4cf3aa5ca64f9b6326831b4fe2cff175b2a796fb44bb7437d8887715ea5067e2c747d134cba7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6ae19f46a6f51216e07fd159891e8bc124f1e8df3abf90583d75e7b3e313926e9eb091c5e6a43ec31c642ba37a8bdf1265817d6c5c271d99bb0034fe176e4fdced7878d8bbe61a36c051ae41cc13ae43add933eb84573aeb80aab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ffa0d19ac1c435026e3b5057cde189d2f9f91be2d15bc27473d9924b994155a20acf9af74e1ef03b251dda553aaa2b39f913ea9205ca3d9e0f836ebce8b9c78b0bd2075534bcb9b1cb305098b1ba61eae3b8d146acc6494933fa1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde034f12fbe6ca92d28ec38955321503fce402f107f37a902c2817bfc592140e57d91733317a9e8063f46afc762cf61bdc9d507acb28f7907361aba58ee9c677c76a4ce4e00037c2b784155ac9f31f19cca7cbdaebf5d82f2d297c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e132cfdbf36bc496997053d74df3d82c7ed247dff5d1a1b4a34602dc970320545c1f7805dbc7ed163868797dad4c0425ed4cd2a811f8f3060603114c72dbf368a918afe7cfddb82afdb9e86a224bd072a095798852b6c7836a69c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78b027b47ea12a1a5be83ec25e61fdf5b8608ff5df0572d44d58609d92c4f1d76f469d99418fea7edc05240f6159e8ef1152239654bfbcaf2bb34efd573c8993eb5d3613961194536890388795561e907ea34793f35bcfb56a7165;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1863064319742b4d7490cf8a950e28aed4c35925ea45a556fdf59d85ec53d47a654592d0e149b764313e6b8d941a90459c4c7081f96cdaf968cfbcd9de6a6855f5c3f116f14e435e68fbc9c2cb309c13636d5e70b0666bf6ae324cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3bbc93bce3bf297d876e7dc35dc9791db2998d919ef38942b1348f84b4595d5f813a485ce81e4e9d9408cd829279c1759e93a61a7faeb135be7195aefa2a09b917eca95f751188f85b5a06fa6c80fb1ffd6b52e42efa165662f1f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fed859f698119d6861dfe017aa4d20367580b368bad19f40c5f1fa31aab50a460f0e2e7f3c36c190be18af0e1d47883bd24665cc8eea1fcb495dde66f97a22b5ffe4e73d9b5255baf8100408ba65252c143e9dea4916beb64e61d6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4abafb5809a29a7d84d03855c1c89270c0cf05d604fbcf71ec0bd88237d9f03466f52cbdf85fc214e712a22b5587ba062f4c78ea350c0fcd7fe2ccbdb6dd257e45ec219075d3180ab59f0ed011333a348d420714aeda480673b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1763ff240d524210745a832d82442e6b2f42bf16fe2a08c6bba5bd7869b22ef223e8bb7ab225fcf5103ac7baacb618e976d13bb41b036bd7ee25edea13382f51dc225e89181ea1136eae47563178b1900b2040d1dffe4c134bbbfae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1160a5c4fdb3240c55a4449ba17e60eac94ee8ce267a8a2d75189a81866481484981a1f88aae46aa3871dfe046abae0135fdf7bfba93304fd4671a25722863a3ae48136c1b445dde51c21cd8333268013790ece0ee33f9f3224179f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bf4521e3fc541763388223ab525ccf59603cad5a744d5086bcb9a45878cf54e326dd728828e8ad82dcbc510186ca1344ffa96277c42721ec01afc2823f475409e1fea53afe05e02adfea90cac8e18573bab643522f3510b4c9860b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11483a97a1563f0339f4f39979d474c0e129c847fd5e840c76b88a98074a1d6ba56bf664964b9dab4915be71759b47c571a25d0dbee1b061936f072dac235ce75813e4ba5c8c7925fd00756c18dc9e86980f3989119475c5ca92fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1999877e0c39928d18fa7cf62b90c6e814d9799b01a1eb66ea4ea9af54fe9252b99d66490f28c367f25d1e9eb7c5b36f9fd5d9de34c592db6c0a4b2538991750bdf85c515cf4808a1a71fab8f7e483d471e6dd81f627f3d06dabcb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12986b6f8f5630df566bb54e2fc61c090f77267cd93e5ca4f7865a2fe38450ade20bedb4ca3f0b29b0bad9be6b43d61ab85027b8b0028ec4005e9d81eea3858fc2805ab5782cd7a4e2480e1205e23fdd9a273a772df00c1de96cd78;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5c2ebabd65bbb1f58a6b7921e2bb85db038b5a0a663452b75de491fed906d0eade7a9b58909680097fe094b362f64aee2d1fbc690db14421509053f4228fa9e0a5e4e24719f0bc7d9966568ce9127427b355f45a9c766753bc7e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cacc42ca908b8d213fc0de23f3d2ee1ec04389e4c7c3cd38ced9be91dc9df48e0d4379dddf5e3b0bf5e5de60b48c2e1465ebe4a22bbfa0eb5d9a73aa729ad37c12b71e96639c1f10c85f7aea399ef82d9bca7f117da294b26413a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16055422a345fc6067bcdabd7c88cf99504745674992b2c557e9673644708f8d2c44842764b6b2f187180e37660aeb24e39026c64190af1ee0d2cb511a864adaebc6a922f80d5507c5f8fecb1583ff19002f8815ab5d97b5e59a353;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185f7d456661548e40203dd03dd05aeb07d29caf21f310a852fcaa314074d01ab4c9f915561cd9a8925bb99f9200511d94da55b54671a4a06e3183673c7d17d8279497bdedfc2b66fe7bcb117539781766e8d8c65a32eb8876f3029;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8bc84e12cec9378e7158d3a8e18c61916fc9b8272f9a7d151372b4e8976aee995299869aae359b9e8ea6f438f236e1e5fd35ba5744681c793de0a22132e67b359673b7622217e6a150b871441e4f6ccc4119b4fd865f2e3916ea5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he757feeb03c962aa141d3ed31872f9926d5685c1c39b6fff89f9be466a97b7bb97cc4463c107eb8c5ba3314bebed90ec0a4d59592baa095ce78bd48921064623b12937b5d1085e7d0ad36fb17f29e8d68f9cc1ff0705042d44fde7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af1499f507db941fa8baac2de97be67a410046f183687087ecd0108cc35553515620edd7bfb489813735b2da710f09eeb01d5b4b90749ae7ab097c1e454bb848be9bde2d0155f0e98fa25f622fb0c0b22604602190024a802ccd7e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ac0eb2f3399d16acbcb213116d73cf5f4bef807e4415f395727c3300489b76a2ca07fc62000849a18dd0af8f7259eb7499c44308b6dbd3a5877dad8d6a50df8cc8bcb1cd18fb05c2f23fcb94ae320bf093f35a1239cfc20f44003;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h174f9545b82cdd3b2001752f6b80bbdc9eba1c168026c2e866c228301a4ab6b9642e0881bfd3dc31082e1e7c5ed3d6e0e7b61db013a6120cb9d589a36d83af84d2521a7ca64cd68a6e3b1859f2d53e399e0327600fbe94d3e106892;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b485ae429e95d9cc3b6415ba0f0b57f0d3d354979eb56ee0f4904ab26ed834f0ce243278e842d081e56036d57611b5c53408f13fece23472298539cb11857457991a9f1593cf9870fb6cde464962e0a2778a34ccbd3e01c44a1868;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b7f92ffe458b96c7c869c354ddc8bc5ea8ad55a7392ac2334ff491b96a5dae0706e918f25b98a7913be5cc866c56a67592a28e20060bd488085cebbf0d8c19695c784d5803375ea9fc0b2aee9c8303e890936f320c098606519bf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc3468793f028d591fb9aa0ca225dfdeb4722a5eb04d14b671448a44dae308bf3ee3cd571d90f2bbb10f508725797be91695285bcc292655f7673051025f5174726193a5a5bbb593ddea35e778cbfaf54233f6d32710b7eb5bcadd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6a6b391e5678162f27b4b6eb1fac74dc04104087c075d9e6f718b9c787e2d341d9d4fc8cc45c122b25541a304eac053fbf8650b79df0c1c76def07b431e281f1a679cf32178971a03e5692ed7127eabf33c197c0c29b11297d8c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1f2c3f12230ca6a0f5deae249bcc535d6d80307072a51ecd353012980f682881898e145319b1e58cf486a8c4da5edff6de08fc6e80c8a49b2d54ebe44fe30f3428fb268a509f7ac453db2b3a2ee7ffd4b6fe26e190a4fc3ee24d3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c9ac1f9fd2b9c2dbbee218594ac17f3f50292c9f9c3d2ee1b9f48462952a6df0e0608e162dbf797e5f757c2102125354aadc7c21dad831a6967bd6153e3ce6ca5a3a861954c19c5e4b87e6ccb2c65ac8f843ae87e78fd13b71ff0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h57bd16d481ec628527451d0a403c84b63b4ca5aef9b5fc5aa8bce5b8cf9513f11bf8e33d220456dcc59fcddf3ae70c3c8fc1d53a671438b8c2008c9b0b8d9cb57871c40485e1786b43c8b20ccd58bb3374daa8280f5b7efc644c6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95019012879b432d88a4abdb3c8e39d9b5b90f14242006baed65bb14ad415127e9cbb7575d420ee6737a46b53513a06cea9ddf8a6f481ab95251a42290311b0cda536d22686cb0effe1d553d3967aac79c44221638326b6de48420;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h462dfd40d45b624fad488518f11b26cd45950161b1a71d61c307691171eb76c94c8c3a5c255d7016086fcca7bb321c6527870ba49a0e3580f28d1fbcef13f17bb478f8c14a3f84c3b0dd1e4c9fd434d1c0d9ec66bb31453c51f0ae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e5d79ea2952cacaf9dae2a9a1be96509f6f72f28b865c8c424afadbe2eec3f8be4b6a785a6d88e6e6168062214d5ec9ec3f7eda9a8ee588c8ec88619c626d4f61b5c1eb5cddc902a1c3c15d2ea40f5e612c2fd37c26cd62a866b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf74c29c9562fc27c1428d5af54fea60989cdd8421f93a63413cc97c2c8813506d842caf90fac38c421ed6f9122633e136e86cae37c9fad9f71db2b2e8a6965ad134a6329322c7758ede6d2d3c10ac16e9a2ffa786731dba5b92aed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c84167fb73b4f36e7459c170214b071dc7dd3d2c04e5c73b473bedee7583649889dc476bae9965de4c753081187b7f4153fe594bf9882e05ae455bfe8bbc4f8d547bf815eee4fe86bd1d793c4bf5c2f83281ce747089ed2e5faf4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166c21108d333588fbc93057e2987e6408fdb380669db6aaf0ff8739571eae3727c27f056d90ba2a48149f35e5ff70783efa674d9575586928ac0820f10f36f5a958b500bbd09f22f4ca75db2ae6ee3c6a2189eb92288e2e706e85f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0eafe3fe5be9df6b590824c539e3d9a207a951c72481f70ecae1940787205221651c041797007e5f5f0c71a2d4e71e73f04ea45fc35941d5a9e7173053e52d1f20d1b0383cadc50b397ae22dd2a42e1d85a0c9e9ab058e697ec2b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha828f03e7315d1ee4f26430d56097e966e7c7db51ece8c8f19c0fca596caad3d9c50347d15097269ac626351d5c5bad9374f4bdf760748fd9e2f7cc4622424240b4f43bd3f9599ab637f09ab299871837559077fc483e242153f6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6095d62aa201b180e1b0b5a5da17e6512d48bd296b03b68b3c12a8b7ab77117cda212bfa7091c003674991d4f5134d99c2a51a3133331b46183fc847aff421cdcef721110e2bbe0d0eeba15bc3b05e7f43d382731e822ceb27e278;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14378cc9d881d24ef30fe451c230e093fbbe4c72d4eaa60ce94dd9af834a24865e5b799746375328836a9fd6e8f955b913c37498b39a4ba26ec8011665fe8743b5f6b304c665e1f8a06c5bc2eeccd50561d32cc6640a36c9c6ea389;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h812a6898c9adf89f20f8055337d390ff0a699c3fc554d0208693f041074d472860a7f683623d1d3017556763e615322f3c36e939018391e6033c37ab877ac1b2a34ae562926c346a6b8bfeaa27b46cf0d751bee7baba359bf749ba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193820d672d4850fd1994492812cb9cd2c4118a9e688979a107628d15ece6c22528634d7be68663e24b1efc329e02e5b195a862452ff60d56e0af8580d191cf7a0f1f0f47f7021c26aa8c0ff5c75493c80042d07c4207e760b1a0e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11202a5e5371c832fea66a65233b89a058d6e9d26240c945dcec2f1d7e4fc497c812afb56fea870232388c82143b35d94396545109a1808e6b0c05833339e83b6f536128bc31433913097fc1bdbc21336f69332c442e8b972c2bd66;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156bc277c653dccd3e1fc54c97b35655243114411680da135e0deb3114dafcd9241f4d29d2bd68dfee32d485862d9f87c00464f483cb8fd7f2f84a761a6026f512f00340bc2abb905cbdd2a3b32a103dd31e2248a1f636198c170f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121339e5b89cde5e449f7f8181199f2ca0ed4ef1934d90daeed0a18ece9c92375f9b85a41af617328e24262320d49cdcccf935b6221ef7c3017a27bb651f90bc130f710a5174f552bd8742f05884aff0c429590001c7c2bab0f96f8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h166d340321ab402e1b4cbaaee9612376c39ac84498be6eea42bcfbc0a486929fce7c6f599c0a7738662d878e049b7fea360fa4d97d28a247bcb950ee9df757dc4cbd4fb1dc3e2fda4aadd9f7255eb3e0c0543caf89ee4ca477986b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b9e4d5a432177247f1c7901f57b32b61728a42d6a7ee78964f0a3d7a13b0b48576b9113e7767ed8f029baa7ce9816942d994293e62094da9bd8d53a0938704e85381d64543c5965f1985dbc8de170bad2774e321178cc85a3fe64;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10d7cd3b884e1f1d0401e9bdac0d0559ff0d26e0aa365edbef447d29c202287a11b5156554321a74def958ad965862ee70942e337f70b30e4493b4a16476b02c5dee34cde89eb8ef01982d3dc5904b26343ca3051179d852112199a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb578c1799f03797e8743c99a5669ef8be1cf714f1745e36b0d32940e73947b60fb6dbc78ec9aebbe8b5c1955df4aaa2955149afc3d1ee95d166935f2e73f33ed36b1883902228fdcd8becfda13d22ce36bcb27d0c4bb8db9fb909;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1517509ac540fbb3d82888d927be90333f96d42c5690ff198ec0f53b4a25ee0857d9d7885ac7cb98ee8e41d9902b4dd1e7b7df18eeda39de1f5fe91391134070a9a0cf217c69a0b3d4d2ce2945dd80f1504af27b5f27d846dcf4252;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d4cefcbb44ebe7ea622dff662899e639c0732323991ecbd1a37e07c5f171d810921cba7fde33218516126428233f0365199601896be16cf7ceb69c60d5852bcea9588fc7bdb4d9850d03f9cf792ecb2edd3ca55352397535dc5c4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc0dd2d77017ad0832155e2db5d8ee4f908376551e272a27b8d648a4205e59daa9a57b390cd911e07062039207bc1fa63bcf4c11f9000417f14f35bd3f44967abec512fa1fa6e1acb2822c1eac3426dda803b5e5fa548f7633756c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf4727dcd3a1dfa881d60945e8f8d4548eb90128b0dd731f7b1e72dc8fc5f54d0734d7f2e340dd51aa275f268145d67033a9b7ca2884e569484f57105bced65cd9538aefa49e59fe3fc319030df35af56bde81af0ac17d0d609ddc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h894b5d9d951690cacaa83d987e8b62e613fad9cdcb42e01b9092ac790019cf054b804b8c8daba8de3ff510b519bea9083fa366a778617472420e95d59216da55a35df4f8a32a8c8e5ee7cc1257add5adce3b6e6c4cf6dcc96f3082;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde3bc56d9a9ba337fd23d56c92127d3b9abaaca5da5cf02c77194a33d4bfbfc7dcc3145bb67da7ad223c08bae059513c69140d059029768fa5a2374502e661232e65b6e6e843c4017c650dbc82222ec821a5ebc9115d125f1cca97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha63406b52a5738a608344507516f7f49d2e37f9bff4ae6e66b0ffe6ed651eff0a7cf9740685d90f3cfc077a645440c9f5c3a4418d94d1ac4d1e4f83c84cbb1191f7ece7295a5366977059f218ae4146b625da6f4433502af370af6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c9b088ef35ae6e9a1e77ee0d40bb23513852fa91b25193c1c2657682e62b63fc67a8bb3a7afe5cb6876c5da158690953b257b7930a6432c5037be2112e4fa58a2a546cfda451d625404c965b78c187fa4c7b8381905f4b9b0e083;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19658ed975c863b35bff0ec98bd4c078794bd686f471463215ad395961d879f439208804f1f0388be6fd4a4a85b22c0ed84330fa18e6601af06991fb422310947da1bd73ca88a802fd74822681a053b311efce0bea8a8aedef5740;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4e6a86556251fd8594a92fb9fb6d663ba34bd78ab620911111d6ac7606e0367381cd1f3a67be79bbde7a10560b6e06a4d4613407111c9f05b73b0b35406f7cf4cc78fcda7ffbb46ef9720ed4b455f7c4d1fffba8318815df271e3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1235386d3d5908ab2e7c3615f193af7ce72479ed4f9356418967b79af585f3133b4331f9b43fca724766cdd12442258d4dca9cdfb8a403b85b0a7d7d82481343aea9d99743c946261ab9f94bd287e7b17a381deb6cec43473bf2a71;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce81369c45a6b110487396518a7875bb3adb620c09a9c77ae4a0b444e964b34ed892f490b5ee2ea6535ef6e6d1d293691486f69cdb1f80e1e7ef19433f368660d8b7cae51d3036b138812b1d3e229291c1f6d754c531dfd55acba2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1163187aa823f672f950510442e22b3f58e9c5ae426108afd4f9f169dcc2552a822f2a64d1cc215e099b000ba0d82dd464a183bd57e12d8a5b7e965291643f35e9e1721947f0edcd3717f8c0fce1d172571773b26c678325c089ebd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d749663ef33e5b0097706b2769f6c83f0c408e7280649ee1b9e76716162f9ef4f4d81eadec6624fe699f28af560cd26110eef4e68615de763cbbd69a574b6d5e52bcf304eb3679a7dddcd5f5557695a4c72679bfb697db2d4b759;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f6e3e7e185e0d203ff852bf4cbc873acce342f09d5d2e7fc185c74d66be7bcbc9c251f7e0478d8c63fbd47ec58e68513f1f923c874cd319ac4f73abc62f17cf4facaf898f87b3745d80fdd99a9e0c9bdb0664ad33153755462b5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h482ec068f000a144d371ff06d8c9429e568c6eefc5718db706abeb5e1521452521bd3e0c516bab22b7447a389fd203aba02870e84579dd07c15d896bbfd66eeab0fcf7052dae9881d353348c96e56732924f8d2815450c5c87d8ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1245149e01f00a70b740027e00ab249cfd482cac3555ef3766b528f3957a9c2f6d636e34a64c2664734f259162a3376c018b1c78f6354939f98439f9d4d5071ad03c83d4a7d787336c15b9d471513ef1a21b4f2cafca5a6a6922101;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h173e3b1032c3fa42ef1daf5ef88102de56c90773e88dd3b4e0f94c313101591d837442e6f980d5ece380cad5b3b0ba08a0493f540275eb6dc15d0a53161254eca0ba665a5a27b2eb146f6d6b7de1a137b58daf479ca6a82f629e6d4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfdd0678bd0e19b4e1baa90fb26ed9e95b8d511528fc3553c949ec4df4075c8c9973984e48ea6b5286d931ffe720f9529b267205dcd57378050ede606436ea0c0cf23fa725eb1327cc3875dc707650c1b80480d4e0617b135519edc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7303d0eafc296c0cc7a8b5405ac4f994771ac8df05d02dbe8c144cba6f87a6ffec5801f63e9ecade8e373ba602e94dfb995b1c9ed2b39a3bf86ce4b408aef05f12c55af74177b0921bd9c0beecd8d6a70c87221bde63b2c4ff4a62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e76bb28dc0242bde9897ad624c7529d5c0ce92c73a5edf4a20bf0aa39e0951aa293b48a4c791dab931a5b1d4b4bb30304e6c31d56f0edc399a84bfc56f7a0381dc25f0d6d2a7e6e55793f6a9badb2376b44e01a2c6323dcbcf911;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ce1b93a4c08248bcff304c2aeb5dc801a400d6060ea967842234031621a609dae372dcf75e44f49a39b060c48b4a5243130de420496c7ac051db794afce5cc6f7ed852a979716cfa9509846bee7a31857f2035107aeac073dd987;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbe8286a32be295bb56cf0d0c41dda6719a954c9b8983252f08106ad46a56d92f193890e365aac6e199ca02934758f568acce1ff44fa3bac95482d9d9894133ec1c723ff04662466e5d788d31577b7e6605f95752e209d18c07513;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h805af408bb1eedc44abefcfbe84512427a59b67dd153d881b2a92766cf4f1504b3c1b4dcddf85499ab34c6c1c798686b6a4b3c35d254f11add9adc578c362d5265526062b8c371b2f7e8a3a7cbbdc89c91c43274caa28b7321a129;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b8e5b24dc2b9416b67f14c1ee21ed5f17aef2e68a2d6bdf4afdaf65a17c6dd8e75ff6a8534c4ebd57ce3fb7959556bd9b6687e5efaec4d84953d6d9cfce6853e3f03e46d213dd4ecd0999e1ca55118f52bbc1d10fcf5c7f50f78fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed517623de0a3bcda60968941bcbb38577c84582964be56dfda2576e2b0a71f635c0b720540b90f5c5b8e8841cdce09a0dfb72f65a2e970cb14f64d05be04da863acf6849ecfd185c27939c492a556ef9353ed4abdc13bebb8278e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h113a317d383f1ec23321ab4f2aa5038a29d1fa284bff391df805a93bb766c5ac1feed72ef39ac0a8f69a85ccd8afb8171a30bd089ee745616f8a9cf1e8ae642b5348424d0c335ca5edb1b1b1688cb4940f024bf83324f8d37dac41e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf3772b2d0156ac39989569f1fea90be8b32f7780bef28bfd46cb030ef624af4b4a219f6cd820fa7814b51ec8d1adf7869ee2da40382a04b6225b2ce325f35c406224b4098e171b1acc4b3619c80b62d61a11e4a41ef740d870fe08;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b7a656df7aa14f67d8b4fe44251f8bee61f304ad3b72de78abfbaa5cde9afe4a8a54562c3b3bf06317e4c353101c87e8867442b9d3aba01766bbc6b3cd12454d7ad9ac359fd5a45e731b057f21a5019017a21567ddb74a5fe6f2d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141db12d9e81c96c2170edebe8d0db13690eee90aa4343319293e0f392c4e1459a3f12db476c5a6d0778bd21b336e7c554615698ebd6a662b21e315d804b04671c38bab2ea31925f6debba56937231ea6de18171bc322bad67f6f98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h49905df1a61bd1b15c5f2d920785ef704a5ef16aeb60749d4ec9a7068b736118df1d531c82e61b6c16d1ec8a5590520146061a1743529a657a10f96a11a62696046da99b9fe66c9f35154c8426cd5a8e7f135aa766f1bbda53219c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce85085d4ac182f303b6f93f2537d037e037232126cf15c7ddc45657d3bca12a36991f1cfe923e55cd2b56c721d973fdc20758a8ac1df2ad33f44defde74ae89728c5defe80b64df7f76c02596f3b1ccf59bfad2622fe3fe8474a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d999341d7b3b83631848254062b7f7eb21d2f87dc723276ad422d44b78d2b935929d89a575ba2e7adfa132083f4dadecc3a6bd22d0d2364a2872c67da289be0e006e74bc6e862348215cd38cfcfc40357d013f76270efa26fda4d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h39a0699240c9c9dac2a7d017e5ea076930d0eb38e505898c0aa9447a6a767b51aedf5122f560953f24f61671cea7293dd75f1d6c563febee2fe0b2ca5054c020c9c8ba6f9014ac41643a971ec33ca382a4e0ded498736e1a3e88c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15eafb58a691f808e1f500db4f016cb096980febf1afba88d78daa51ae0ad70ec2244b0007b52a4d8f026f1982ba3682d7c1e7486a904bb67803773cd1bac0a266731b891040c6171925fa6595ea8cc23fbe904d42b1c4d48ea546e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17553e3bdadc1feeab2c01ff16210e4fa9a98b102442839571a5b8aee51b1f7b7e979fb02eafba3eee559b77f1dbd0e576215900a968210f513a8afc6609824e4c162ba43598635b9aafca6411bf722991459f0dee12455bc821e10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c481cc8855ad8a2ac678cd44c9f300cf9c8c40484965c0ad8e87abfa9aceddb2dc6f7e81c60122d5fd5065aafcdd431233b68630438d934f6a8e5771a5b6ec6b8d9ff486b49e86524f61d15f2cc5f5a32cb438091e55dcfbfdcc6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ec0489e57125d6b4060636c7b05d66ce520d51e1034177fd4ff40ab1292cb777bd6c4bb82f406e9137dcf745366b6f639e97ad7624bddffa77efb88981b4ee469c81e0654a1c8da4adcd8922666c5b6dafc43647922066fb5cb42;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b69281d9d1c197d2078736dddfccba3d7f8341424dc56a7ef2a2a242b8ea7fc8bef697bb34612648cd64dfdb85365a2a2d56e2cbced2b42535c0604d65034e028b684d2ba34bd161792ff02f4d8bbb590694dfe2b6877b4a7f3de;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he84f8aeb5dbe6cbd2c8a22a227deb6841739287411164ac03a6696527aafb2d0a856a2bd8fefc443c245414190d5a63770b7f04eb7a5968d0beceeb28777c52d785574dd48ebdec81f09db6a0c7abfe4c9a2ab5d00e1e50935a831;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17f44658e37d3f7a3a6a3f0aa8a4ef6b32060f21bd6c9d4f81f002a6a886871f1e00231e2ee2f9230f60115265c7e616e85bde0ef8cf02f122da7fa9939b64697f20f56f2195fab3d506209c436ab34fc58c7857997f3217a72e7c2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8ef1577322c417fb02c4315c3753532917c31feff059d7fb6d220f426263af234a527b378a96e38bd78c0a1e0e25eb99d0aa516a1608d7680f9c20d3218c86694467614670a74d3050969dfe99606bbfff6c2917f31b9db1d28a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc4dbdb1cf4d56b033dfcfeed3a9b742a5efdd4fe0f2ad7854ef63977d0d789b484e21325d2ddaee1788ee11a4daacbf2bd023109c9e6d0afdc86d79abda81e8a15d7255e74d5bebff6c3867f2df9523adbe76770788f16eab802;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148746db2883a2276c6eb45b688a16e85e94daef853aa86e687425ab23e0154407ae2505cc8d200fae782a6d6036b72b5283d0f39021f385af78a75962b82a2557f257b556724aa7536ec22461d4f09c168f3fa137bccd50974295c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb633dc6c73ee1dff3c8ed5edacd8ca9e42ec34b5bdbcb39968c8dcdec71a94670fb6dc2730f0c9cb8ad2ca00b74d67192765c6e237d602590173d6046097e982c63754b0b852f4a2c87c7eea49cb68edc098e60ec87e4c71836d79;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a908db2ea532853775259cc7661d0183ec33935f687ad99a3859108e0599cf686da0f3a60e1f7bd2775e2e5af4e90fc550bc7f429a28d95dcddabd9d1c0d2832455dceb299bf7b9111e0f100fe9658d634810964dfebfd2ac4f00;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f37356a316299719457994e1af322ee06aa73e3b51673f588053bb0c0670c6754006f1bf627dba2b087f0b66aea6d9b278a8284e44afd09579846fb597097b89ff44a726c2788bdd0b56f8b9a9a81cd0f1c71d149bb311d4fcff96;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb093e3599bbc6e5e3a67163a2863200c5d8112f362ddbc58758d5fc26f76ecfb480e4d1a2573978ce75af72cce0d9a9c0b100e2ef753a404c06b58eb5413ca21892fb645a5cecc7bdccc768471ee9aaa6604e6ad35c5e890a7ebd6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188d6d8d26fb0819bf8e48fab5fea09db0a422997b3b8c6cc1a2cf3442a66ba31ef61c15261f333f62375d0d5d9b596218970bbd22827c147db9cf8bc72ce7efd69207bd5217cdee6c027f377923925b21c243bb87dd70850b4b038;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cce14c1ae9e0e0461307830946cc619230bbeb7f7dc9f62843de3ca2f1017bf8ad49231a9ff2e4b6bd96886d714798d65b4f69197e956bc32314f5746acd78d28e72795f9bfaa923fceb603af7bac07adae11c514b7c30c19e0aa4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1032230f9a1b2aa47e7e88d7ca0a61ad5fc14100ab88dc6b91077dd31bb16972697ac217875c1b7a8e03baae09f0007695b8ef41bb138cad790eb8f0e6f4e7460fa2057f218c63ad7ae9d888439a2b570bd8e7706cce2c808464c6c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f092b6e042ca92905b06de495230ff7449eef0086a87ea06015a818ea6c93e90c1dc1f9dba2ac953245758a3978404db35954b0fa8137e54412206b4201f3434ed020c3f071791e32a853885bf83d25db1d983b2ec795eaeb8e0d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h859c56ac864f3363e2293c673d1d31d208cf6a76fe2c9bd06b2eef4f166123a570e1d87d11de84a445a2101b09cae1ed2e20e7adda19086f7665cdc1474159597a4b038d0a3aaf0841c51b9882e2951f3d708b9c84d286179bcdec;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b42c8071cc596bf1f9e6e66e68ce6a97d7a53b12b17e41d3b335355d7e9c6548c8d9e8e00b1d72a1c1569e4685af44e2a9f78ff094ce196e591e16cc96c529f462242268e4cc25510bdafe0690c2b8655e5f566f60ba3b70e9164;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d893073465cedbb9e275a657510f2517e7a729b22bee5f4e0a05fae5c2420549738fa6a9b2fac04926c752d59a049554da048d9c24b20013c960f2664b6844b01da32db71454968a043d0c7b4faf750c5587a05a7df8ad1d65373;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3f36dbbda1258a13f4ce295bd856c3981e10398eb869af80676ac2fe346cc8f34bac08ddb8879af53ae4b6f1662dc6280ac258e83c377f37687209961e768ae81e656bab89a6cbaf52a6a92baa034da8c90b32ce93d9c486b91b7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17eba63e3921d87179fdf5478f2251ecc49333bc1b5b50f137daef25f268c43bc3409916720cd796814e6cb16c89f57e4748c5b8d245a803daa7de39d8c2ca477308b5ce5b8fb9aa88bfe56d3046a6b74309d972547847b15cca2a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35c0291d4771bbe2b727dbacac570bd8175126c19c5656fde57ff937d344b60dcb2228076a6fc57643e2bdab450c096510d6afa0c32b4953ff405feaf6a0128a6a6aa4ae15427ca8f11d7bed1d8b8de6270e0bd72ba60ede21ec25;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd95afa91e84862e82074b8f0d4d1842c11b5c1a83d99e47841bb28e9273eb428789d57a9fcaba1c838fc757a5e02ee6e9754892285809530313df9575e4ebb6f9eee24e11a4c7e2ca6122eb0b291e165ef40b5b8d7478e72e7201d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a7540703f0bd977d0712b892145eee50b913e391e357b7d2621b9e62cfcd11d6238a2c0a904b10a1f61080c6b5a1d31f55dd493a9c1e9c2eef62e05bc4c4d8b738032e3e1086b813423579e8a5096b202614562ae24cca967df8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e0dcc5098ad0fe538a32c68bd2d9b8d3c56d1b728b649318e63ff0ce50a029f5d07e00e3f51ed6a0fd5d876bb065c955c55b4b350238d71b7f4d12d587f740a80bcf57391b75f883580cc3c678bd5a76409efd96f5fa2d50f951a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb724cb4f5acfe1e3dbf6c6ed45ece7c7f499bf2434e5b9516bffcd9c95ab9d7aa62f088903a2098115ab8b675420a42b6e30b80feb3cd0c5542a902917e1691893f9557f1b10527a5a76ca2527a77d5177cfb2aef88cbb60d68791;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a01c4a0c8b7177438add4c17b1aa033b83915d1aaee6bda2e6b306c129d0100b1ac9e050676653c3b724b1f5ebdcfc4c26dd5750098e17089c75c1c82c58dd116eb4f569333ec4a38c177b943ffc85cd156a8e057787ba3ce7b5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c76833efc4d2790712d6a327fae9bbf4d5d6de5c06db206d52f9f1c0e6e0a0772dcb451ab55be5454a68ca56ab2ecff8f238e58e6e10984d6f3dbba760a7bff4205f949b5015011d6f75692758b0177ceac901e027f9abec4a8692;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e43b5db2117475f962c8e797a1ca52485319407957c17c9b24fd3b5c7e3e106d2049d1f28f1b51b3e70eb871c6cb7bd4f0771f6eec6c1495f0af62fe9bb167ad7f7aa8d733b26b2fc5e060d545f09ddaa07daca945815b3ff8d7e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11ea12fec43c76792ec28f01090e8f53335de0597c06fa013bf93ac6cf164fbca682d81b483ba6e41c2aaacb717294b8a0639b0595f5f3158ee7b4b9769dd3908996fa0d05f56401654c2f9ea0c0942dce01a8af686f66c2109b174;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1addca181e937eaa8edb2cc54a921e718fb69ecf29ea2e078ed02ef6f0e0c2d5a3859547928cc797cf303b52486bd7c6a4f2eab1b009e900586cbba6bf49f6a07627bf245992473552b1c41fba1c8b0c3c810e0b26129a03eb017f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16141d54d1b580dc1a96afbaeb2aa4c66bdda1aaedf5ac75a41020dbc08cdb2325a338cd9f62ec4211578980fa56c68969688fa4fa48a4a2bd29f7d12550574a89081a26764f53c3456fe558e49e875f6de8287dd817913ed61e425;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134d1fd9d7fc69688cf7a1a44bfc81695d7e40f1a39841bb833aabf51ab325a414899b16055ec17ff686b3b217db5b0b97cb143b30a8f2928b8f76d057ef96c30c20a6fc357780efa0a123a39c9bdcc7a776c73be37ad28a20b234b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d278de9ae875a6c571f80fc2bb0364eae98716ea60350057dd15e16f4fc61c9d7f6c20d8566c24607cd80b2691fd3f189105a3792852e3bc51c10d54ab1933e6bb0298d6a516eaccf8bd442199eb58ae56dc846152f68dcda52cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4f403f3853f807a64da20344c7ef55cbf50974ead53c555caf2bccf3ca1878268f0d196d56aa9bbbc1eafb270719959bfff1c0e244fb3754f2d5f57f6fb1081e911335360efbddbccec6298ee10c9a451d43df0096447484f3117;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha778b232f2fde9da9d94fab219d4fa2966b5c68ceb2fd7dcadec9f23c2df632aece3a242a9da3323d2e9c71adcf48765df0eb8213f07b5f8d046b53a0706db68a618c05cf5ebbe5c840e46c39a8577878dfcc55d7365b7affba3c5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d6dc8a2a75677d7f054abaece4435534720a0d107ce4c5f965323d409599e747ab9dab3876e8f74d9b6eb57097650bbf6622d2199b2c93f71fdcda70f23fd662078abd1a9588aaf60224671d19b071ebdb2628f60384fabb3c0adb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184e202bf0b6b310218424313f78f3ca3f9cccb4d0f90262d8654a1ae1db9e83db11461fc09d2057bbf65e7714863ea260fa3a8b20d89460fb97bd00b2026f8d1d770d5ab4ba205992cc740b923d5759c0928a221e8ad92cc37cc3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2faad03fab8482b422b88132133bdc81d63c5179bb793404c99bae279dcc9a3e01e0a831011c6a859fc9eb87770ebacd483952acf378d1a9a38b1f34e41054ab090694813e01410164801dd8703fcad30900cb0275a7c8c9188a5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce19612cd42ec660f77d04de3e8041dbd03c916478aa8025257cacb5bcd427c130e757517c9d52e926f4a70557cf7277211d1d4bdfa6e0138fcde65b48b9cebb929392d6e0ab950807430efa0eedce94ebe25011047d2cdec42f10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5da15ff6a15e1bd4aa4f79ae429f453f11c787ce4cd4097ce0f764d0ee8e6c96d5adeadc3b9474419e5175d325e08c33bacb9457c02c27f256f3ff965e08b3f634a654b8484edb41e6962cf5cebb8668cbb9114b7e01d84526d420;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc35c9ce49782e767d6b50d15776de7e455651b94ed3e23f351db26a5b1bd1eea77bbf5546b2a5caa883f54100b945ade33872c158e4fea517e2768b6cda39f58cb79184e7e67be459e5ee045ea4e8bf9d5297f34b319a72ea48906;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10ac0b054209d32927b445d9c42fa09ab11f31c22c96ee326dd680b548fe4819a53a209b8067ef983b762ee77757971c1bf3a3777088d3ff48303180f066ff9c863ecca8b2afc5ce1dd7732fb0cc4cd5475008f9a93acfb4f6a9822;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haab0599ff5b77d81706a57e01f40bc321c75cd655ac6a3913f9a4367e47416f2e7541352f4e87bd36620ea72e0ef3a9a570b8118b29e167bcd278a819c4cef22db4adaca57b1f94dedec928a73fe6f306334c01f6080779d6aa296;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7aa9ba107328c01523a2995d1ff28d2d27806a4d9bdd3d495bed54af8f13f00be9f5bf17b451f548baa673202b2002303e1ee3d4c8e889669893f2fc48e8a78620424374f56bdd540c42f9880e67c998cc28927bb78fd36e91a16;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce4cf2b2ad9db3c3f1f55509b33c4fa80effaeec5e064713dc45424a71a352eb255e4d1208ea4d3b3b0f8759ca07cf8cc39c6f5c43f35fa7c746b3d7bd2c6b882ce2374fbe8a602c3540f7f25729cfa0c66562081d3919b017ba93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f1f6d0020a30bb338e66032dfc59bc660b2f9cc61bc758dc3f75b8b9eb00611af8ee0cf3eaac4dbd4ff42add73b0f6eb584c42bbef160ebdd83f6cf65b4d68ee1aa88c0b7a5c2410e33f0ec3f8ef27a84c3879f364ae2f4396249;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f2631efc9d77d7de454858939647f5ac11269f95a1b11803bf0a3ecab960ca54ad4f96890dbc91f773e65392a151c496d2ec76997883fdf80a3d045e5054050c4cd53b32708a56efcfb9c7de7b4da8fb341a5616dc9a4f6457a00c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h112cbc9b28e7aebb73b104b93ee421cd180269a232e3e4e311c5a009e751cc7a50486f85f2c277331a6d113bb847f4209a10f50a3e443d293b2d169da4882dd403cf8e9f64f43b2a052782f3007a1cce0fa6721fb37e9867f3274a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadd3117a3d2d5d190809c2ffa56d0766dac366918afef145faf605fde5675d5fb5cf572a3a037e2c012096100324163cde6585b297182a8ec1f35a7ceb03479f2f55b5cbbe81367288dc6cd2ca4905606f84fe819e67e0dbc68ab5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f61933c4634e520291de73559e6f59f6b9afd44f77ca8211d423204c3640f6038dbc2dbc89a3acd70ecb7795c44d62cf9fa5eb24234ed18898fcc67fe6df9ca4f888d8c498f4560ac7d3518029209b05ddb3fbf43b0961207c6f76;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcd2247b014790b0bd054d0e9c1fa037a5e3648d773af3ecc4d73754894a0255953df328c4742d3500545a22fb69e13af5ef371e918c8e22396f3e65d9804fbe86dfb977ed36a1e5663d01709e88465bf64d71b02aa865dc47aa85a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3607aa17083d3d92b955c25a07d1dcbc345054239e3d9b60019b382fdcedfdc3f9a19a88e724d76194cf7959c546b40b0d899ea3d5dc90e3692f7e60944386fbf8ddf88ba35473e4e9a8bb2655bc54ab4925b45096167a15710cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7b24d5aced38237eb8fa16e8033350808e5ce1e040d0bbcf763826e857d523a13a48fa9b4371818b5743f7f27487e22c838ac79cc14987a53fe2d6bab7921ab4c8a595ff8fa49fa220c5cf35b0db5d153d076afbd0973567af6e37;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6dd64add32be22768344fecc1448a816576783d44502b395a5e542508ede5fe48a8a0e98062416bac05db3a67c4ee09a63be84832079f0920d5c4ae2e7dfe0a46d433b27d7e84dc00975d97d9b8b91dde7d76db9a77fb5a21faf9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c7403dfcd9ec282620083b87d067f48d921c06ea8bad17bff9dbbb40f434a93e0adb7189ac0dae70571e072e6f108b0821865692ca503e5ba53b27510f55447ae9bf3c1fc5a300705b3af827917bb8766e4fba051fd3065b7328a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h414adedb3be86acde5e5b558b73f0fb45f18e12ec9075aec722feacf556793444a00f949a2ccdc1ea7a017aa126cc7dddc041ff29bc044aa7bb0787e2b3284f61b29344996a80ebe0c6b726344ae1d3c16efe33d3a98968644938f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22cdcdfd8be27929c9b2eb9519a182b16ed100db388ffd2431f62f3ce80922260d17d4d1b217549536dad6d6e9de29e0583be6bda2d62ba7fb18430f7f0c70c5af528343324aaf6b2f5f9bca00c3d50fa9ce057f4a77de3f383b09;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11bff82ef99277202904d01f6574cabce367fffc64ac9e2e21695c8a67817dcbd54d7d1cdc35b9de252308a3e0f73d8c5a1d563a7e44fdc3f7558687b324921bc1d361263d36adef25aeb2337dde8f30ce8843cae5a528920b2ce02;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d2503dd6dcfd351906f0cb43443e36c848f3632ced5a8b8c492477731f7b170bc1d8f46d9cf70259903d4e27b1aff1f727196e322b0271f79989eaa472b639093385986d31afc82d53a6272d1e6b0515e210f625c2d4d9ec45cb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h675eed9212c0d156d6cdee51a0c858a89c0ed1459764ca94a41ca1103dbdd9159f540231a9e4754febd883afd576aebdec034efc54a0729523ab51ec0fe1e6d09ee02b157de79dd634567b26061534cda16c9604b95ef8c2e443e1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1783ecae6e17143cafb89a2cd8e84c6d05226b0c828aa15408c23a7b6beb23af8476bc107f0e3059d3ad069f7a68ef323c55616dbc27512009f93b677fcffaab8c55b2e520405376545a66fb0eaafbbb84b4533e162ae5103300057;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a3038a483b0419f61f3f9ae273148be8a306c3386e548f493a92cf703ecdec68da18b1289ba756680a84c2096ff3ca2f1620d46fd4c6324bf6a2478ca8ef526c1adea2161be5b7cd1e2c1f5ff01c0006d841bb36be4a47d727285;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fd9fae9f0d638b905ac3d7d87a1d72549b09e9b59e2a049691d34ca6c17b3572af20d2fee79b4b77477cb6140745584fc069b5d84c280f894a7d2c4b005825162a255c1c0e7b2783558d17fd83421f0c7981edb9ebd65bb03121f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h253b62500b5450c0355c4f8603069348774ae83dd5f2e2e3a93c8310e6b3a24b2846bd1a57486e6a44e5fbe3370f11970f0d2dc1d988a9008eca25d1c1a39efd394038d99fd14918cc475360fae79e56d10a1b1b9c017a546e3701;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6610e988805bd50f33ffaf497184f8db0efc7fe8b440224980433bd5b7bad0ff4835662f2dbaa7c8d77a414b355a393980b4c721dd670224f2cdcd4d64a84897cd0a3a6b9272c9adb712c037fbd45b84e7a8107bd2e44b40941a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4d835639754a3b2fc3b21350d54b5f5d04735720ce70467a35a571146033bc7ddb52ba6db3d4510d808b0515393e7ee48ba6139bf6479be25fba19dacdb3101bac0bd7dc64700453f3c3c007a7c606034e1230737b2f4f7938d60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h178bd1756f414bf955439ba70726128e75764ebd14fd053ccb38c9f32b44ac568c7348121c67ef0e4489b031da2311bda10ba49760f6dd8d3a851857ec70eb9d8d475054ce816017620fcc580cf6cdf817b17d43d706efaf7e50629;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4aa63ce1d6eddbbdad3e828e101ceb423b1f5af849535e01e8f88e904a7d20e2c6fd76bbbe580795bcbc14d56530bd021966f4e81eb24cd7339ed111a685700a980c82bb248cd942288c965770e7caa20a92c4ac3c9e4a118b44b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16bb446085a53573847dbc0cce8ef226e7abbee9ff2dfdd1bcb9be2f0cc27042fe2b2aa2d8ab9fb1a0969c73f6f6681511a68dea8fb756ad00181d75199248bd73c004fe08daf5a7896c424bb92f7821175999fc875183b50af6218;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h633c953b31b4ad4c4944eddc5911e0244c1d770697448983cd80e52ee68548379a1d5017c6ce4c1b2ac6ccb1736a06068be30e97c44f3845dd326872a956f5222ffc4495fc6b56778bfee912e21ce14769969ee6cec235a1ab5727;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18b31107e69cf1a484f43f744f13563be75df62c9abb44e76683af05feb440854eafaa152bda880ea76043816863275afbb0cf13dedcae5b88fb4b95e369ecd8f2e6d6d929409ccf1d7372da5c6106c505bd635639c316b352bcaed;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1884c276af19daf3d9a1f873cbc3d7e424c3677d32a27844a44e7aed70dc5cb76a9f8254472244233934d00f43c09ed37de48a5b068fcbde5b3e6d558b6fe3cc128b3c2d9e035dcf04dfa51dba1f9decf485c7efc3cdb0ed13ca7c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111c2ef14d87e1982bdc580fb78d9dad1f3f872c7cfe11698188fab5dbd347f5b9199688d82cb47fbf3eac2b398b88119cedf9f42780f40049a65f084b6c20b66c485294f2afe1c0cc3332f5d0788b14077cc6023a99b4d9a267c3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd84c921fcf5e44a6b34f046cd22162548026885a1fac68c4b734dc91ba295ec25f47a7261ec98b855e6fc8fe3fc0f23fb0f19c6f3599f34266d8b24f22ad1d12de69f022395ee5da51b02963e9eae483f4440bd49c455a80e0c9cd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h878fc44545b176261a3d518ee0a2acaaf64f080a2a9279e07c2e42f4311671f13334d021b5c07d36978f975fa03f60cdcd18202b7676c885f6656100499fb61830651bc49b368a9bdd2155edbb5c9f0757f8ed44702cbf23e40f92;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f0c1ed0ba55cb129dbd673023f262ab7dfbf571055ca710baf562ac71efe97fdd2e937a2c3713b0c3a2f589103920a389de58c56dc723d47dae4628dce5d23ffb6ed59eab2f3bff92bcaf22fe6dbe1d9069437e20097c75b35217;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fbe915c2001d2d91cdd605f82618462961612abeef4c24dbd1513294bf24ad2469a3ef55cd83630ac250bd330e9e72e2773d42bc0d2cbe18675f3751b2138f545bbe8a204f230b8ac5cbcd43b5ee9616d6bd47b608bd41a358b60;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b40325178af64e32ed85a44a6bb58ecaad304e3b2e2493ff2ff1fd291a9fdc77a05a5b1fde2e70d795ea1d0021820e851be803622fe1b456012c8e7e8c6bf6f8966bc50db0916d7bd1be978cbdb34958ce6038537e569ae62838c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17fc86533a34a5ac1afcad5a19b5a0d0d84d09b081405b18510f350fb5df34955306d408dfb1351675af99f877574020c3d0610eaca8fcc47c73c7ed61907cc8b641bc1d004183e8179b932edbc1fee6bf1f4c277b8fe80501f016;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h146d29d68c01a9177b27830a38b6923939d94beab75b8b56659b374b8c1225a93542ccb8d74c2ab68fea1a1ab128ca4fde43800d5cb547a1fdc2340fa438dcbdfe6f4f2267771ae417572998b26f0303c68e1459f10dc74fdc61adb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d681530bd3bae265988d2152c586096fc1a5e441e70be799f1af16025df4b610acf75027718a1c491f8cf9ecb690dddeb3e1d7c3149130052c69f1ea7c043251891470fe99b7b6eee77b375905f650f32df0afed41109279d82f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4a9efc6600cf90d934027e1c44773980c74d3e37707d5d1caa7c4ddfda11decf85f09aa7f6354369d6f2433cd7362b54347591ce4b7a7a3d3315ec7b7f24d2ed2ffa418af9714ed339b253b21f866a6d4949320f54b56a2ff29e03;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7945f8ad8e4e0d25c7a515bc6bf120a64dcfe4615017b748aafd2f5b329d30643afcb512eee056bfad86f9226759a147b747c385e3be87a849ba4b18e54337dbd09e4ee2ad36886d047fa0b8e1147ce1c0037d37ffad7ec43b1bba;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7195a8f22c1a67866c37bae1fd5c38d6f2ab11227906ecd19c50ab9b3d386e6f32a35b90e778fc8d157a096d3ea9fb4076db7774717d400321927a596c61542608c15b9b3273c7f9f8f37eef489abb5d941b1834c4a05c3b3a79f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1415ab266c2886a60c6ba1ced700953d683bf89011cd089c19c798f5ed4fae0157a51d41c384dc1deea219c2cbef99b95394b9393131e6c032b0923db09530e7b2232804171d491e63ce1fc619f47ffa97310ff7ceaff806c71e90a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9ff1d92519131774cd20e30b9879eeba18e12c364ce735b0df2ffee601ca83c48dc8e96b77d29022e058bb5c9ce8c8de73454f7810b4f14611313a55543e5b4602dc3b09e7e3b1cde3b93841df0d43fcdc682e967340ed329c3d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c45f2993471b86e24ce2a8de05163666c16b81d27160fc6c667624cb2e4eda2ca708711f531f69179e2d7b50c04551f836ac354958eb0ccb7c976a897e1ca3c8228b1f8a71cd9739f5c0ecc0711faf44b4e3837092a64717d5f7f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1913d5796dac2b28fc73cdce449834e1d2498b9a3e239cbb03eb487272904cbf05a51b115869b515234ba9c17ace2e65b1964b920bf1dce9d5489e3cabadd6f94850db77d43178e36d4b0da5e3bc436c78499b5d8af1a22d29228a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185c9b4ca1df494f12fa7afd64ee4c9d3b5d25e9eaee912a9acddf9013538b89166c089f5d3ec5cd08be712195ffa700828a5034db781c8b8f3cdf8ad75af9ed0a6f5049e5a10aeff6ce836d58dfefd2d9e3c6f1c76d78aff09ed74;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hde8720db25da8d03669b9922eeecde2c9bb610b0386a2f3be15c6a3b36c160549e15158c9b50f8d5383ffcbcaf2cacbfadb8addd32625505ccce3c8fed3f947b506195467f492911070a5fc8dc415e1e4ca1ed7839ab2dc7cb2e29;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72646ca7d8ccb084afe8adde2625c82f795186b1ae20cdb1b56f9e9bfa7324c4e958a9e94bc8c64166ad5769d8798a8ef73f2775a1fe1e65653771b0f350e59eb04a084284f6ccaad6a98915088da3ff5ec0d9a7056fa332c59f1a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h108734ea15c80717b63137af72d96c2fcae81020e22a61cd401deeb322cb364ae09d3503266616910716201ca2dcd69dceba5e061843cc1ddee8a03cc12cddd8de0940669f1585e0a15a55e2a2f539e70664b2cddc8095dd173a250;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13395e5a505e67152a88dbd3fc2688b66f19313e73a59196c6c1c5115a6615dacb28c73f1729a38b91bb51d1f6a398b1fd77a803fdefcc06fc474f6e3d16c5c165abf06ab7ff920fe8838ee5d08454702e7beb839d67dad8d8ae675;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e17ec7b8041d3d64caaed86400c445f25a12d519763f0c465ead50dd0939fe1982da2477ab55d947a998ec499715ecbf7b0687a63f6ffb6105871b0f0e7f55a812a79f1947078207dce35d7b438da0481b47775d605f1c8e11c3c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h65eb4ed72fc99db5ea212d94224595b475bad94dcd69d4e0d9f965fdcde435472b7410a827c365764b6072512b265f422d54d31e62f4aa7e6e10270c09d398cd44e623f532c76dfca91c109272a62ff17c7bfa765822f37d8a4bb5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb4deff2165d32b8244b493d3ef8db8fde1981f6eb4d299186c2101d81447fdc548d6b62ab25ba8194596e51f69113028d757abe51317f7141b2f2d205785e94e5e2f9bea2b521670293f44c8d51219969f70f2b447ce3acb3e8afa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd2eb7e7efb0f0a50085e7bd6393aa6dd5b3913d255c4e086a50d1c0e2d7159358bf59e41d4cf96917e0cce4809fc7c4afadd502878eff870e93278c10e4353d3538f05a6207debce2095fa636ec1a60f3cb40b23474128a6eab5b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b9b7802cc5e7e777ef7e98f80ca32065d12cce755e2224b3d94a1c46da1be5f560061efe57dc4fb0bd340ec5d38bcadb46abf4f15611537ecf63e2e460074764f5e44213d09656380eaf5cb36fc373f2f0b5c8e8058069d4210bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d2986395924842df048188aff9ac80ea01adf817cd0024d226882b8043144f42eef8029e65bbfd476a9b26ea28d43f92d8b14b7e17c5ea90838324cf92eab3726236d012d36e532197b8e5d9d597df32683f3c4a55163e0488050;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c1e1ef5c55d147caf1b997d85d2297c3932344033c38e814785e9dcd0d45466fc8cc989d662f59abcfdd720953a49f26ca92105b75995dadcab5f362c637fcb5dcda63426351d586c8dd363d47a87a3f9a632adb4a0bbff99e082f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78c8c752089aa5b861fb066e983ad83a5d719eac0c6cd610151e1b7ac1211381d0a15ae8cee47a1606d1245d7d98c2d1d1baa7eb9f5e10fd15052aeb3f83c0c29b051185a8f79b96b96cf69857100acd13725308633c8a7371484;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38014b4c2f568acf12c80d03a8db7ad9287cfc0469d069d1a933fd2a470df32cd669f47ee7196cf83ed040c8b5492f89ba1498d6a392f5a5c3f858c751ff9e6004a05383cd555c62f279921f1c2a7b76408157a31b6da4e485df7e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he570d7f9e26e173f3fde823bb480b7a5aa17283723b3ffe1fcee04bd8fff30fb26dfaa5ca0f0d438dc17ec206a4a453641659250b009d17672597cc3e222a1ccf966b99fc6cd0f3125f3d6e761abc1cfd85e72e46dda2b2d80e815;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4435581b6efa01e0c7b0076b1c666b5a80367f969041be8fe040f002e5e0d2cbc74fa5c3a22146159af8f94f1a07f1e5ec214206fb8018cbc92c3ecefc43b39df7147db881d425f889ea848abab704b3598b43ee93a42b6ce663a3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf18eea59361c5295b60fa5f68b3b5947c1037ec8c0047b69d2734593224c435cbb523e07b5b66d205f215ece1723cc8fb26502c1a0f776bbf34a047ee86e21aafc92560fc38d5dcbedcb62a466d7ae50ed4f56c75c637ccd4df513;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha462ac938714352133fa8b2ddd9e52ca46ac0c18ee795f0b4e3ad7fa8bad858e2dd26bfe624d0ccfd36e07854e3bef056f26631be2f0f3bfe8b2ce7e11a6bc4c38674ee587fb3fb46589ebb5e9d1d36b1159488497e831433743a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8a8385099eaac54610b1276b6d42f0d25f96edcf1b6d42e30bac91fd76df22f010b6b4543b49db3effa3f4569cef2a04592ec25e9eb7fdc63bb131724aed64cb72bdafb63e9c9571584406b64e0b0c334ee2a2cd8ce10b6e3742a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9c17ee07ff9be7250940440bfddee786c4f974a0f968fbcca9f6205de030ed8c56f4fbd6cb1112af95b43a70e2392216ac8f2319ac0fd2ff1b0fcabe388f379c7ce0851f4fa553008149c427275fca91aeee92eec83c9222cd307d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193f5ac2cd2d26e58d68d1ec0aad4b42f920f9c551d83248f3104948032cb286a2a8a475717f74c7f9b00779e5196c6d5cf668b2ddbdc8392b14deaa6e3a8f52e61821996feb69639f838c16d64b51955f69374a130f026fed8a32a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h81b88268e849ec2bbbe296a2983563a5fd42bdbdfedf8982f0a9d1353afbcb9bc5fa6eda3ab93f5a0e692ac7ff88f9489c4a224cd400022807a41bac1ee18725bf6cec3120c4d17d91a5f1439240f03bf7da7cbe27b8de909477fe;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19304d601661b8859cada92bb5baeea119476451bf2ef76bd0f2c03e4af96f952facc701145b36a1be16c875446d8ae68b79893eeb8070fe27253b3b593be4a77442d13216221b928e1209f83d8e2bfdb1d2453eae94267309d8c10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18aa5e098fa7cf74e372a09583fb58ef024ae6a85246881b743cc1fea2b9fd63a9219b2b20c606d163ab304388db8d1f0c51468cdc82e9c6a29310906fc2ed14ef9ab7f223430f41141a7be07a427137faa2b9ef0d036bc51a94d98;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19341cfd8d569edc562273a549adb9041f9f8716c4508b15042ad9d1781b5dce5cb79ba3e9a3cf9c6491476a73d7431fd708039b0c9b1231bfebf7f39f5134cdc0d0a4d8886ec115d8612b2b45d7e4301bf78d87f9a52298c0262ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h897a42560c043039148776858479bbfb4713807ad3b98e415372a89c71af3b37fcd5c5b31712e46a3fed16804a7da0c9a5a5a0518dcd93ccd9ab4f1d6d5e49814d889de6e875e80d4ae2484bd5ac34c4f5b4dd7a71bdcbc3d32130;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e31c7f8ef4e7c0cfa22c9707a02277897e93eaca10ba5e3ecce948b42fd0ca37b366e5b376d32a84529813c697ad6cd72d7c2cff6a01bc81387cbcbffb6b8cc4e36be20155103e328b189dea2096564221c15b6923fbc72a25d4b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d9e13f57841c2ea646e7dfa4eb87fff5669c23193c132775558044a5998d24cf670777d618e5223f306908f9dc656bb510a37550efb0967e2f612e5931a807087e3680e47bb4f210945728fa74c08fdef62df180479adc0873c4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7802ca9576c968c2af8b2eac6c5baa59b41c563e2ca22c516abfaf012175ff388dbf39bce4acdd397be1aeea6bb0225dc6f3c125cf265425df2229d055b765c02104753f171e7cf27133d220a21fa21306b54fa71d03e363de057b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cdd335f1bbeb88395e8acf84b2e6cc09bd1a239950ac9622b7f0286ae55dbbd28af935bc29c1ac1ce283e434b561b87a5f575018cb004c82060527a66a15a6b84ae206dc6c2fefe23976f67f27540dac6cdfd9aac4b952d78036c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha410e050b56f4224a0249d6d5a826f18e864f560d72485d5ac81d09c0f9cd03987c79c76b12115062311cc2d310a94b4b9c6441f690b9409705428c45588e5231a51c454d8ac4218d816d13b6ee45aa532bc8e4cf11a005f84602c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a82180dea5c291cf3e8556b980c6531528c7bd7471c36cc4773a659844639ccd9a5ddb69f7b7bc320cbf86e625a81b45d330148522dfd365ec82db7a7167f349da22f1c53cfc0164ccdb1cf2ce244229b117d1f50de2da0124ce9c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7eca2b995656c6c42e300ce1bffaac03f7711a77153d53f884e4c548b0a0c20f696b1992b387f94e34a5e4ed4eac8bf714d6377180ac3b24f1cc1b6a8a0074ac230c5a643f9652be37e65b06a87b107120611c2b4a820ecafef3cb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79b0bbb04ca583368d21e201c8b3f73508f2485be21b7b3ddb90af3613f2cfc3a7c89aa864eb05bad41a09310ebdc5864afc32c9f6cbe0acf7ef316ef8f3ae5dbede73d1cea0de08aaae84ed1b00d42265e0c42af791f9b99810fd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bce31870ecdfe7419e00d423fe84e8e8ae13189c98ff47e1447ca21a452ef45068e357d65b6c10de61e09b031eb2376ca8fc405437626e179acc2bbfb91b498d26d56584207cdf987b8652f201af3446a3a87bc20915d15c15cc54;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5518d9b9abe96ce47173498d9023b8f181997ff6530e64559c9aa2b7b90cc4cafa53592b2d31a8365640691d4ac0049594b0b3ca8bebd1aa1022d283049351c582d5e1fc764ec04ac84336d9b060f38ca8293978711a2fb97a55b2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8eca2838d0cb5183a36151daf98df179c31a0abda7ea596ed760f67e64fa5057bcd094a8b9b8da9133eb9e5de8526208b1a35c0076a1b413f71172408db8110d8419b0c8d557fa962dd6800e04ab05766893fd98c93726c7ff295f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha7b7b04b038a2c6fd51cba3c4b00329fb99a8f410df72aa7bd1143a23ed49c10ec24aa307dbe616e9a26a70968ea45a66de6f2f6983c3dfcc653bde8ba6c083c88c527c9f04f96fee3adf01970318c8acbbf9d69fc97f9c2c80585;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c43242985f361490063e03112a93d645e85ed8264221b9fd76d3d77dbf810c471376292a10d967c49782e414a8629f52966816b28113aa7a7c9cc15282c16341f1865b74721bf136db83e1826372df4b70b6e9bf67e69a59b48b3b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha552f4a91476f6a6471e7bc49146442c59837c986361252dfa88ab953175692d26173a69f123571ec83f554f8bad331ebe772ba496112488617f5a8a88a23c43e0eeaf8d1c7527639f8f07317995bdca5cdd1c9aa1ec3893f26f7c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1958987a2b800dfaddf449373ef38371260e6f10c2ef8027a387d71843805b77c3cb8e55246ea2625edb18a65a8753187146f2d1f49de8ae07b59ecf020e875a1a0a07a9b9ce85164b28c7b72f562bbded13663d1808a5ed1d68e93;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd58e401e0c0555b0b976233e1beb2fc2d1d630f9a4abf2a2cd27908e8c7a95b2dd77b14605d45a9b339cfdd0564382d71d7d0f6fdce99e5601df7c34d290e25d7b89264c093c747246a6382cad472c634dc2ebec0b3efc98edb3d5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3859f7ac87e1c7313b03a31a14f150ef8c0af1c13b0f4e877a5e9aaabb075fdb3e9b0ffc953dd1cf90942c2ec30cacc30a8080aa04701db0bcfacb1014ee593d37beb2c6c51090953e051fa80236f4261129687e8a66ea5c1150;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158ad73f68bf0d232937d1852e74403e75feec53f5b17fbafdb5723e351facf204037a362258979d8df86fc42ff78fd871d8033e320a3b476c75954a6253f5673eca049ce163d09f1428828168ecea3ebadf47834999cefefa0e426;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73aae83d28a4dcb310473abdd574c63ad0943d9dd240e35258f7e8070b92e8129bae0eff413d2f2fe1bffb56ede9f1977eb62e5b46e86b14f93101ab31dbdac17a18a07716b765fe4df8e8dbf5c4beae2c5a5f371d9c56a8d7105;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd3c2bd0d5f38d98183d593bf9867a40a0762f752fb67ef12b91321b5a53e451cff5fbec0b9c46de133472ec2be7a899d3bac18a2ed78b424730ca4501a458656627245b7186d64f13cd23e5923dbbba09f40c6e6a21ecb9b08529d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f09189426c3ee511fd21adc5a737b76a998a520cb8917d274acaa7c2011c256cbbf045523ef9dbbcf632fd9fe84c88382e952fd241790dd18455dfdccad9912917472f9a8731012e892f320ef88a97d06ee42e0811d224e577e07;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16da31ddc62e4b55e41568aa56153366e39f6bfb854d366cea77b50f1f4568914ba40cebba9f6fac35d39e8ded97d56f30671537ad624b046cae21e2ee4ca1a58de8d5d3f6513ca86ec4454f73952d266dc8d97ded0bb2a239bc07c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c2af5a0c9eb060a0cb1838edd7359c7cf10552ada8f1cd427c9c7187f6ee9269e39869546a0a4d09a7a1242bf004c27a1a9652b85de0ec9d90eb6fc3288e35c2c4c86d4cb77ed679a2bebf2ed81e88af305d9d788765f4a07c48d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a3b32cf0e14883121abdffe922c14afd62e0a7f370873732555d17e451744c70a152c1cb5f4dbeb3b9ad91ab58f890ace631bea4f54fe57211e83bab448f3ac75968400ab2590660ecae1f0eff6c1c5d8812da69f4c74b524776d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4c2f2434c118ae88cb3b45b3605e94b755eb0a27bc1310c0bcb65570ef11f3c1c87e9327e8aa3cd6fe4483a1c31988147af5838a5092881fa6595e04c17040a2bd5e24f01f57240d48fae9a71f5cec380ca997eccff26dbb6a15d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa9aee87e3e4dde37d374b2d6d4ce3a305d0a437172023908bd01afdc3ba778ae0df5e0e76f77038adf7254054d8ed646929bbe73aae2da8e7121f2d2a38fbb3a0352509de29401310748dfe0ef6872399d9fb75a29272fffd61c0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae5e03948fbe2b821ad664cade3683b18f009e4aa089a337f8386047fa523039412a9e30313325c54956702e767d284a6c5b22f784bd27d8561b76906e59db0cd48e6c60936dbe1140115166f6d8e627224ff2196e267cecb1123;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5e759c73dfaefd74a35714cfa0c6e9c49b414ffdddb3bdf990c0f2c828657b9a8b8c5f3bf8dcfd5bd5609ed5c70dce3fb57317817b0e45ce0af12e2ae62e739b9eadeeeeacaf6cdbc454e60ad971127e38e08cef507f7c17844b0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h879f65712460db1a983c5fa2d30d92618b1a59b8b069f9988bb9ad36bbb04942fd40d47491a20b229e74cf0a668d7b26fae0fe7c1b41d8c7837bb47bf41ff1fae3cec698a28e0d0f1fea1b6032c77919ce3cb52e6b6db91488979c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139ad468d38890d9dc2dba4793be84fec2c4d6981fdc9b635189ce9b50b1d12b005d76be26340d0d8fc1474ecb64f01c81175fe72167022cfd8675749a421d8b1c3f4f2655d4a7f7133d9bdb41684820dfa36fad3eb4dac5d91d271;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14262560d7a290704956394948c491283a3e052c882efac43733101b9484323ae7cc78306d7d7b32f6f230ca4cd9d9ddd1c4f5a63e17f6d2414a9b81cd1bb0d086d63a3f604ec5bba30369ec075263d89cd5448c5c12f9180b721a1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd2b154ae43ec575ed0a3001e8accb4870eadce504f121f072966454ce35c1c4aa6610c29a02fce9b04a72e4d0cdc2fabc00a0b4e6e0c77a5bbbc8bd83e5afbd463fa41dd8733716dcca671334f03fb44f6b7c4f4d6dbd28693c99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h604d5e874c7967755a280a08d4513255d69fcb9ce8121b5f828016bf7ef4eeb134cb59302947d8219ce9c4147bab6108e717118cd4a9cc8910aeeb6531046070a75a09133d99e84314b6fb8535f211970a71bfb0a3b34361b3dab;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f1f127c71ee7308c06323e91f8e4e840a9c1ae94d7686bf509297a1a807ab59d52471a2e9fc6eec045f66eaf93f434a90f4af433f68f15e96098ef5c34b1af14cbd0c90b4538eee5c78fa357669b3878816564ec08afce72f5ea;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15bc0c16224234f108dfe21378cbe07d8ce371455001c44a1bf333d5a3ee85635f9de9eab376e279db4faa2ccdad210c86777a57018f88e2c1ca45d023309fa69e285fb1cdeda15cb471ae322d29057251a8632df9adfc86cdcbe9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c29540a7019615e207966b2c1f5a7a9fe9bde5b691d6b9da84f5dce2a7050c574e38fc53aca3b5dc360eec71ff15fe802c2508598765f9c9831bad8d37cbc0bfb6ba114779e9cdf7e28455c231a2aa6324e84231b043c96b5dbe5d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe94e20868b77db78a97b909fc0fcc05bd2e2bd9d95902a4e218bb11c5d9f251195665bae2d9cbe1ad06aec92af8964b4fb1d7cb29c09c213a3e9b84ace20d351fd2d69096af1ed6f2e808a28f27ea2b40fa0458ed894e2b08cc99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h167036ab2175e227b5c4b8c1843ab28cf9eaea022583dac094a1678849f896266890bd2e81035accff95e87cb73421799f7dd28dd6bfc279368a545dbbacf5698410871140103854ec94cc3c3e0e19d9b99980a6413c3abc39bf7ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e31331388ac5e7cfaf0acad92eb343c21c5eda511b172fdccb5c4594d1ed5efcf487799ac4ff0f194d014f240753999b4105c582ecf4fd40a0ee9e1f2308c351fcdc94e321e0e18b2483673f05caaadd3ae9fe78193e0bebb2a9a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1187d5501d91f748a55d1026bee862b54a2cc1dfc0772f300c5302c8e1e3a1fc201d43985660187b033d66997cc8508eb19578d9f8bdaab58298407225c2eaf44c764c5efaa829b4aad35d76db31da709a9d486e21d7400e46b33a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1015e8466eefd1eb5096059366d397105576caa88173bf2ec545318ad1f1b8da57c221b5a45066698a1d113ffc3731f3aeabe22317d5068a24ee65492710f79bd197a325ccd61a40c140d9550de56441ee478fe850ff887fd5e414;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15b04030d327e5a0b9939a450ef1fae3cc57571fc9caf6dce659e184f6251baae4a80c87c73d4f65c9364279f46a0934574d648e7d15b7099b34c3b8a7cf5a2c6713f845314ab053486ec3722d7bf78ca84e2a5c91f461b30377820;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12ae5f1c24fa1efce4ed6790749e9750accbc717e063d43fff01efde84a0c29ccbfe9d73046fc7ad15403c49e29e07f9ce7673ec7c85d8b004310196a052b5f4d8ade4255d4fcf263738b93359c71b0a50383d07d2fc1b1eeb7d942;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec1bfde488428fb03d7dfce47e3fe0745d403a16af415e8be965c6636f4cde3c5623ea5b5f988562fead7d9a30f17d751057458206dcef3ef4b04660331adc1725ef54c2ea213e3be64c33fe50724003c4a0458ccd87d0a3614270;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h592891e107e1a25af0954d133481f2b419a952ca372f97dd7f94c7b720208a6b7db8e1fd14a7a83e47a7c4f52bb0ac573c110f5803a29ee9bf3bc92421d4bf5c392da5176208115ea6124c026e238740ececd1a9699ea5f18d214b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35baf5b0d656e841e2e5e3dd4663a12f0bb39939c77e523393bfba822cd5a43641140de1f3411ce8c42bf99e9d77e057ab216f9f55ecb1c85aa763b465d20c7ae71a3ddbaf5b592958957bdadd6109c04f091e184addb8b78fdfa2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7e7218e1bd372c41d2b23d207fdc87da885b34ebdcad631d0acd3cea60b9bc8a3d2eee0558d1b8be1e808ce9e390c8ceda09ac1eb16e0e2c194cf08dbe84553acd91511c33a1a276d8c25cd8c196da808f62563170b413bef46d6f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a64c379ddf22d0bd8dabf6407b503ed6c549b12d5ce9b76cb5078db554d79f40616a3bb688c0f0515b4b7f3750e3238c8ab73b1c3ff0cf5758ab53b2e648a962d1e078edc5cdef658473ae97205b903d8503dc52a67b3901074f3e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ba931f01fb53ebc4727a68b13b61f35fa9fb232fe06c18b9126081d91cef8e16367a664359fe61396de0bdefbca32a3f7a69bd9f3610943f207cab4eda684eb50f02174fbc89ea60e897b5efd3c8fa02cc6e7265f2b72378890d1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128ec47544091ed21c1c5415709e7f7fea9387bb877147b50170cd2ba3e514d69495e716c6ca1b56d4608e7c83b0d950fbbb034249a337a64a0f07e4e18773893ce20ccc00aa4c3de8282c4d6f137bc0b56aaf82f09888716d26d0c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbba07006f26c6930dd1fabb7778c1344fd7ba2d4491b802ecb464ca0898117e6d6982606726b13c786a9976b8abd69513ac5ce63bbe51269b66799b13edc7ba61bbb6fa7e0dab5e748dc1a9bf9cf9f6da4d632ff0f5d38c5d4769;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h40b74c9884d6a238bec03b9bbc268bb258ffc6a0ccff223c36a5611ac24758d32f07b800a255feae7b2a908a754e99a48dae4c1718c865883d424a26986d72292eb55d3bfca676d204239f7272d41007ebea30797fb5ab224b936e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80b2e8eba4d2bdce7f4ff0d06e640aaf365807eda32b5c0c02c8cbf363fa3f378fed1144b4263c351d7c6af1efff7346443357585e40d867b8198229885c37a9ead77663962e36a1d26659b1de4dd21ab5a268cf825d9eea931ec8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3f49641d581a658b659bfda4f24ceb6884ed79ffdf8837dbdcfcc76943e358aa967e608e78c402058adc26900f3b3c8af10d610e5241ccd516dde75d499f408b95f43c4af8d62c5194d6e647f63bc95940a679eb7552393f21f5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e3acbda3ee906888bd71cc039d3b4f84cf52e8a32967896d6232c360b081581903718a955b10c93ec601a563db40f5e0dbfbd4c3ed748e5cd83ce0f01aa11ef28436d0f4e65b31fbc7a66acdcf96c75760c40a72653795e5b343c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67cbd731af67153a3b3852e0dde52fcbc0e85142948621c8b268ddaffbfb55c4e8050d49dfc953285d27609d91c69f56209ecc825c6f6686fb3f60e1dd9ab0aca3c2077fda891a283c80a7e0c1f97e0f402a559b43c284a1f43e3f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h782299125752435e1ad0d5e927391583d4b7ea7d8de1ba93ba7b5f9d0c81cb6d09453046c62d9e209082b08f0f4ee27a1206d6f7d2395b6f15a020dd78d08e65587e73d1d7cb4659cb60c3474049b42699ae7a61aa866b1c2e787f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6b1e986c66d0f22adbd7fa238a243191696ee734057353ffa500db53d77f9bda29d6de045092d9466e454ee2c02630210989a8f61f9ce09b4dbe6482d47b2ef1bb47d043e5b4a810200ab9c8aade698215092071e612523b6d92d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h34336b4a57ff56f3f917fa39c191f5963bb265bdbb80d3774b4c68f96cdea6fcfa043c3070777cce7ad7a3ac3f9c7ac3dace6bfef5085106ec3919e75c7cae6341bdf9aff81dee376fe90a7400a7b1a0e1a4b07f0a0933083d99bc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadcb44c2136bb9954e365eebbb1bcadeaa50f9e54d3085673425bd06228f6350c3c3e1ae6a49833241a3b3ac771e82cabaf384e01a9c7bb06e37e1ec83718eb7009d0722083adf8f196959df8d205bb4698e5f626db4fef6606e82;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7841eebfa6d30439064e9259a6fedcb03fdc89ad6574a63ec24c74537174a3893dce0b1945335b22621515bc092fd9e0695a374ce87aef56f360b254bdd3b2fafccbfeca0c77036c02a287a2ad1c466c933e68358b4c0b62c1b176;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110bf193bd9a6c7bc292ab72c1d9138d3e134cef4eb6f047adc900b7b0fe591cc9dde23e6822f8fc3674d02c9b64eb0ab0af960cbf2e9330a161be10275135da0b7bfaec9b4ac3db104f8fc4dd7ffabac8b711a7e3ea554ef406af0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f7fa887c6f58e95035745b7e392beb06e1336371d29e3a06319203ef8f67f86a8f167857bc214b19d5a2c6f80300aa362e3750687108bc12d5e2d01432f0dfad028311bce0a672a757c9237e15b936885e98657688fe269e5f21a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b16d8c5add29fd2bf8b3e8695d26d7d38420012609a69555ebaf322fd56640bf402b06ba5d6fe5f18b9cc566d0d767988bdd1a602e60f63c2c2978cdf44b75af47a8beb14af3166a754e76324c13b6a6c726d10e2e2b8f0bfc2288;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1919cd172c7a9b8b91cd8f5e7a52dac3f248e68d7bee0607d56a2cac189e957e3589747fae77bf293df125fd1f728f19d1ff8b96f437b30da0e547a4acd7a7c4f05103c6c853433243d4aea2a930271ed6585847542cff13f584352;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8a5df855824464a6c40d3e6394a0fd708ce84b2ed3a8cb18b2815055f6613dcfede4790ca2d3a5f8e8212ec4bce062f0188a65cc8acf16e817962efb4f2b00e27354bfbf8e75c7169894fa1c23cc27733402800666f403e224c7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d9c8cd71b854e95261427a928acad5b1fa3d3469a6b506dd2f63dfa0427e8eb4af1000149e72b79d2a9adf7cc7a14a242d916df925405b8cc53c8e0812fd1852bf7fac9582c904ff8b538f771c13d89d7d72f2517995bbc0dd9eb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73a8be5458019cd91732fdc40b22bffd76c07a701caeaad2995b2472a1497e07402dc1adf9532ec528d42de51c229bc47fe5df897789be4d5b46a3ffae04135bf34a4d6e34f03e16d38e7cdf61524eb4024bdc04a2e7abb810eb9f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50f1d3d2f17806e51044c3d2bb7e8e427f59b3c2f3462111ddd86a489373ca8e8111f0ac7caa744579695ff0485ef75ad657d44ffdeca743e96b7a3a514781a494a0b3411db860857505ab91d4891976edad8dccd33375669f076;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cb2702d7c7900c471fa2024898d595913246e2bf0afbcaa6aef01d7041c1a3b442697e1f66e831f0a8080b44371f1e7c65ada86f2d6a6831257d711ff88a4388495169ab9671b15d854b9b8bb75b281fd1bc93d1aea2bcae81c7cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed0b04dc7abb5ffda043e50323bb0a367b4b615ceedcf6a3d7e7646ff7eabbbf3850d6963b572d783b92211392f5b3f95777e51d3f0f9760efeab83c6af1b564d9d3d0467928582934e6b488ebb5752e9d3c2c982b0c3eecedb8a4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1acf9b623d3f423e900868c22f4594290cce20327e57f904d5aaa184f9c9291b52ce922bd7af6357e715a6fe59f7e7d63f8a4f913fdd4cbae2b6952c783f27cfc22575d8bd0346f752e3f00b7f5f3b8ec41d9ab087ff85f83fa30bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc2c067e7d729dcf79866f98bb42e123bafa401e4be2786f168c9280417629efc1fcf78de2d460c637015e281772ae1622858fb043988c003106ec8995ed0b1d6489fc5f69947ad1c53af2a19ffbfdea3ae831e653866a11f0c19dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bbb68207c0fad0333f3dccbd46795e6c086c6cb587622a8b7ddc3ba6c77be7090aa176b7f1a1f4dcc50a9431be9551145817bf22df32788d3d74a2167a5f55f7bbaf3d215d6893215775aa9df229a3159a9572828a247a01a166f6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h168f4e91e9edf922ad349d9e30e8ca7033e8346b17055972234764912ec2dd32cbb52632c83759a9a2050d9652e23de960a08acb91633a978c877bd902aff1cc8336364a8bd9ee9319721dea8e49e3f43ebd7e743d068f1d67250e5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b3b6ff43b51f71396b09f5d9ce8e2daf680ea32d631eb0279bb3f727112423e7d828f11b472ff78f35daef7335aa3c073666501d74d69159ada29fa538e9e62013f90cfb7de676e9911ead4d5c34bbb2434cb7e539cd330d5bec8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14007899518d8744aa459fa228c9d20eccc0ec0ff0beec91ab01a797f58b2443b424494a4dfe790986f1f4ec56df91fae888da972a57511420ac47928768839dab7da263dcba864ed6dea775623925d2819f0412a84cfea304345f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce204a66d4f808d1e3098e03835695b5d729dad7c0182909b510a44d1029496b648dc1df76c615908e5eda4c8d7c7cbf118b38035ca0457bc64521fe380bb60ebf492bc63460931a36f608d31f6a7d0c434d910ae0236590f47d1d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haea4e2be482f1cd19e9a8c400db20f7431dfc292c5e20e230aca0a2c23df6bcf3228e550d450daa6e2ac00c7515ca0cf857bf81188770be3427fb0edad69edbffb3e025277192722de80a7978b6a1e79f93d82ed7a194463db2357;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h102c3eff27aec0c0ae1d8bb2e4049cd194a90d964f2b5c03ae3d61a5b40e17a8b5a743f17db3883e0ff01ead91389ace7d53b8bf69cf9838aef75187c2e61665cc33ee68185a96b761c2ce8cd62e85c44211158e082c84c9b7838e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8f889cd16d0e79a0284a7e9112d60dcf85dff82cfc3a1fbf41d25c5e6ec0d2a054ece4e946aece488a944840fb53d1bc61081eef1fd0d9b4090d1b55aa9f84285cd56091298169f6abfb96eb073ff8fc4d8f13919b613314ce095;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1041c9745898cf64b5f38fbe70f76aedf7f4b4d2f005557040107591b2e6dbce3925bce5c1a4a25ac4a5faba5cd90e66ec2d5a947e783905619531adf3b6dfe0e4e11a5c1fd4e7bf5bca26ad32a1d83d888b25e571fc8b3f9e03708;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a549fbe450a2678526a9147ef8d7d3d2e156fbfb4d6a0f2e5a883557e8e05740fd8638f6671e3b08ea9b19393e56beb57f28c18d5f30d6fff379bdb2e0c7fbaf2af23d17582bcba963cf634e56dfd1c14fc19980e19b80189beaf3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1139161bf80d7875cd83626314d77aaaf0a6645dc7f0e73ecbdb88f537039f0bdb550875e6a6f05a9e0e87433026775726b0a34fd6a161b8f6ace2ef7e86061d34fba4457b6e8e4e46e7f544a67bb82dce4217c41045ad866f6d6bb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4f43c305f196ff5fd9cbf7226d723f3a61da96fe2f6e99900772dafdf1aef77fa50811f9573142c36c856a9a2667a12814597d50d8ba8f03fb4cece7347db92b25cd6e89424d8f86fa15540d5823069b533842f77421c1bd8813e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ed1521326745703207d32eee456cbe02363722572b4de423fce5ef1a197eee7c8fc38c358f4726fe17f61bd56ee0269dcb05d3d70796b3bcb1b931a779cb7b650e5c22535395c8f2e472f6a2d7d765062b5259bee7330035ed9e2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12df4c1c0b914747c9f516c1372d16225b6dc0cebc1b576832fbb97b2b6300936f8c45d66ba3c5358024ac7cc3cec767077c33ba7a784a4b8b46a89fa54a39b76976d88ae3cff96875e7b2d0f639dd0bdfd802e7578db5d8e904816;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8106ffd3baf7cb1948c9b079004285360c22e558a65c52c1a0c68b051de132c258dba47c17056c494e937c54f187a3fc6b8f8630808f65afe77a830c98a60cfa1467bd7aaf88edd021d105900beb6195cb978a3b05b894ebf6e8b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e728f1932ab21912c89d443901847776188c97d52dbbd502601828e46d20f18c688ccbcfd61df8ab95d5da5cdc88274704bb989974604a0b780684eef288f12e5186c4a77da16f6b850237b5e0f2bdde557989b72f6157d813e7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b9392676600525608f891c1fbef3746b79c1e4959236778e1114bd640633e0290f5763c0ab724b0e1e71088e8e40bb39be8062bf28ac045ed7bcedb426f67c304dfb4168724c3112966613a61aa157318ffe0ad4c63823ea9894d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf830fbe524577c0dfdd816c7c4e82f49b5216e749f90b1f720204761b213021fab6c4a92c670614b54176e43518554aa045129f56752c4543d79438b4ad5acfa73ce00abe7241baa931dc352e3eff5f9c0372e9dc2b39e6ec90a4e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19edffa7a4411e7c38f7c1c78e6ac713beb9ff5c28cd61b468c4fe32f0bfa0fd94b60631e6ebdab21f9e7617ab6c29829db9b6c95247783b029529292aa5a44e5ce86e4c5b1acd38f1e0401f0968bfe8596303e48b8271c25812152;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he99cecdf5721d087564fc9f1ba925a319bac07c0d82bf6602a709ba976354d408f71207ef91549cf5bdddc210bda7d3fe30a343d44ddbfe5a3b96f67f4044ecb6bfb01b0694f480b537b882aca73d5f6acb696f30ddc591f2fb0a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c7025a4e8ded71c8a2ab0fb1b7d93c9c55388a0923f4d6dcaa7771475b1b25c6e930d4058f6b98c1a34755a3e9637184cce825224ffc73fdd388fec0319753600b9e20f6f30880ec8c77284fe9747f2f4be3280021c91336bb02;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd54612256bccf4e02c85633fea1671de25ecfefbfa6a88455853eec85a13d8873df17b7270731eaa7157b0462accb7d9bbe7bbc637b5a2c8c8d90840d9e0af57411a60eeb8a58b12999e5ed3d5568020b9e0c22892f6440c8adec6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6ea4c06bcea6b6a4f7d215264da04d2a738b9b6a5bebb8ddd83bc5472604e81914ea70fc987f72ae297d324e093ecc67836498fc852186f245f9bc6e9f410ab826bbf5b3a1e66a82b824a53dc8298aa117cde0928c4a4ae2b953d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2335c364fdd8d7219b9ea41c737d60d1c38fffc92717d4ad3a16b7d16ef953d53112bdedf0e4113dfda316f6d706708f91f0427b3249ed710f361abab4176365b3be643db67f3d472ebf1e6fe2227ddce7deefebbf3fbee1452440;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc279a80eb806010426c7d0096dd62a6505533c3b0962a050f48284d8aa77bfc0a2f0c9d5fda29d34fba679c57be949e299763567fca6d6bd2136099680d5e43464ba5fae46955f86bf952ef143ca6e7bfbf7597f927ac00b3ddaa4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc80ca7a5c88a84fe0601afdde49dba122dced6a924a28a84bd65d82158516689c0c8a84a9c9f47133cfc9019177b8f8d88baf589d61c5721d63e3856cff77844195db5ca3bc5abf393a9321b92abaac32c65fa0c5c071b0d2cc151;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197b7a096cdc6109a6334743dd752079b93ff5fd079b1ed8616caaf20866bf4afc9107cd904cf169cb32e56dcc284fc5d28d4232638c948ea9da012da58ab77c9d71a91eed78f154a8b89b5b58570c8bb15273d28a4b5a6db8631b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd16f0a64917f7390028d9fa9a5a052ff3bd63d01e8231b1c00f7fd6ee69bdd7791a3571bd83bf0f1c6921a2414bce41a7c6e1dc8c41af4d842d0f0f961434aa22eb466f0cc7f809192bbd6a8afcbf59fb704c5395230a2a5e340af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1773a317e00e805080e657b3d5d0acaed74f6ce202a1831e244bec330e25559aa3302eb0446a5634f547f39d50a969b25cd483e06e569d8496fab6d75ab1632897bae04843bbdf4dba5931b834f381f29ca64612064828c5fa765b6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9ef88d0d756c0db2e5ced186d132863c0b35d15dbed0525442fa6a6fe42c5339effa1a01b829363110669a8f5f0956bd8ce2650d3e49a7fee5ae2e0ba67a9eec93464e5d4cf66d148ea937795043903dc0d562b149f32012794e0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d5f7261b9484e9c81942c5dfef9efea41b342798961e744c4da2a8f23cbe7f19b999eabaeb74f3271b7202ec92627d9c34257b920aba66cad603d52ddf3d02912aa4f67cd0968194a6067f6d1fd65c98bf18cb6765f40a4ffc890;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1120fec30e1b99a0bdc5f0c49cd42f91902836f07b75e45840f3f59b0d615275a2ad3c1b2fb03509e1dcd2bd8f4844e0a90df9d7d6e3e225cfd55c739948143b9eb89260a9e022006a84f700bfa9c79ada1a75c96411068e50972d7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfaf8fbfeffa3eaf00d47b7a07e3c390bc85f133bbcf6d610df3192a883e6761049a20b912da15a4fa0e677512e3fd8ea33809d4d95dc6333398277ec56a59f9a94194c0eecbc84018dc58d0eac35a4e5d0e8571488c22155240386;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131531ac614ed6ffa2876ab417496268421568f2c38999ab14b2ed6e396dc867fd3551526265814fba7f8160a57f6e3431c16219904d4f66cd47c6bc3b92effad5b047565ef9ea770e1a22ea0d93a8c3806afcaffc14bbfb5af6f62;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h88de95d6f5388a1d2feea908ccb27c2392b83c04a6a5dc9f167018fe87b4e3dd351849f78115b5f2f7a0c0acf5f28a6cae3c556ce09af64312028f45ab17cede7d81fa9e83e01b43b5a8c5997fd15e8fd37140dd2834eb48a73e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1463db24f81a61622dcee0faf7a0bb287df2f2ce6b8318fe0d69fb32c63106f6b39a9c8725bb85b9189f5928cec7707a70d782271e7f606ef28e52d4afea6cfbcccf9a4c7df1ecbc17ce706bfde4883d388f91d1f22f9be855bcc89;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111a6b31f73c14c0ed2e190fbe413b515116e4f93deec0f55a18f4041fe7b84fcc3ebc74fbae0cd2ca636e7ececbb1655ca116934218a26d415be75ae1b25565996cfdcb0ad46b1693eaa2b594239c4590a4203db3db300d28a6891;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2075485b02c5f1bd8a81d04d41812ae67da02b54db9363407f0bf615756a46c71afe04bc8afbd738ddd6c71a82f588d5be09352599b1f866649716fffd3b39fbefb9887115f2ece6db13598b960a1199f5a7c0114866933cb2aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6cae91dee7a27fe32bef58d1692c9dfd1df892938cb16b834a01fa0e0d49ee08d2468cdd0430f8523da9ba821d13e652b728651c50d1cf75b8a37f56844dae30a71ea4f4ff1babf0f68f784fc6905b39ee61e18b2c7318938ce0d0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1972d488891831d48d0d5b876ee464930f46e0d66131313d1b27d97edc3a1b3d4bae351f7eb66365345f788f57c200f8fd50c35a427397d69996451403fee016a525c56f7ecf775a02e90ec9a937ef0a3087bf93e9809cab899533e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182ab5b636add41e0b3b687fa1b6af7cb3f519e8f920b5dad05391f9d7d6e2872c1c7cb9e2aeb6bac8a130367f2448ce05c43ec3c8ffd3051ba9fc8a63f68f2668f8136bb699bea6db496ed43ebe996730dfe929b44fcc8c746ae7a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c21a56b17168a10d39cbf7ec42e08df099b4dd22c86bf5184d26b1ed415d3d84a6129c4094c9926c39db9de11edde44ae32fd1d017c37d608102258312e2bd474814a255603ac10ee70ad786136301169b303c9fb86dfed2efc40;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c8019474b004ed3ce96c9fd36f7384e5ac643b54e121742c5ad4ee0a4bd24a7118140ec173021bc3f966ea6fe6a8640040e12693ea081a9f4e39438a09626e07e22374c875dd9a45aa9036686d9a264c0f75152a34a13f77736f1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6153a545ecb2d94f2d02e052002437ac43e74f81aee15c456d5011e517ec82e4a4c9bd43a607fe3d32ab8786dde6bc89a3e054559f814e1adc0b26aeeee7262e17f8077938374c5716880a3efb778be6c27ebf72cb5203aa216e45;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a7519eec3875b30971050adfb683d8b01d79bd9a4bfb02c302ea75ba9f0cc0638546c98aaf7f9f9bc5cd34af35af992fbe9c73268b9142b8ff61d55e9c158673f0ec47c50c859672e09a8a0714f05d83180fc4c6b42417216da17;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h494e15d6b779d1379324c13c568308fbceb05c5fbf0edde80ea64932593be99c3a4f058e85e007a633ea0ce7ad37e99c51cb940a07926dc64239675a65c7b2fb183e81a08b65adbf85d1460249f4cf20d75b6a469b3a26a6f35236;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e8f39be25e7398ac0035d67dcb22af73296289ee358aff232e361384268e4a41963c9c94a05016a3cb86babe0fcbb1debb097aeab7efa7e448d3ac8622fed5152e141c37f6af7cc64e5ea0fa0d1559286e335ec9c4da062eb7bd9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ec2f75c478da95a7d64d3fe2d1715f2bad1e8ab8063c27a62e9032b5afdb7c3ab2d8b7e6b3b29d679e2856c8f874b77f49796fd0440d09512b1a85b05d57e5aa5916d1ee244aa038ed22d060314fe501408c46788c6805837ce28;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ebd270bd876ae311a9ccda78dc949ff13541c810c69324a61f6d57d2ac97e9f7976d1fca1db96c3969d5479ac15835b27a96bfe391cec21d9498de081a0b5732b97e7f4e3d9a249e7060b669771c86434efc1e073bb5627224b33f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d0be9ef0a5128f1a7f3a0eb6a9c60b60d1eb81a092c145f64f52a7d6bf6e38beccf56009b07959a8dae1dd2ae7fe190853db481c89d36739e8444613e3cda931d86c2d18fd4ab5f5b21cad68b1894721ca3290b84ff00319d31c12;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e43ef8a624ebe94318bc371c6e25b483a5f2fd8f3e57a4a65976e0dd567c857567862c6450a6600a11ab7636d00c9b6b471b23a053516a342035cf5bb2b320e5a808cea704210db4b3a50d44f777e233cd196ea042316284c1706;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e3903345bf60b90ac5e3d0e868b3c3d1377d4112eb4991c4b79bc13bcdfb5e4a6600d70f29cde6fed4f9364340ed33b20894db29f81ab48ba70e8b8ed52071aee244ebd744f4294e5cb9c5304cfeb455ed1d5057d8dc69b7c15ca;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7bc63fd6a73bdf140b6a7bfedb42cdd6c559b771361158932f3d545aef92ae5245d6a4e6297faa023908d06b7b3428657e75a627fae7460a1cbb1225ab16d1129bb3271fb5e8d356ddaf134db0c5d331a3f09687c39ecfd8f075;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e76962c25772540ba46c66c4ea113e3c9f4a4a90c599aa3611a805699cfe1f1fcacb3feebbd0fa86abe93ac9fad2553ca043335635baaea51a7703ea213b2fe16145ea3f77b42317e49e08ffb0b6d0234ac96a4aa7c7c15bf68da0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd28cd405415b70f62acfbd2085df4b873fc939e8822f3131f3056288fc5615df40252926a717d14beb8311aa01ef40a39e31d73e1aff55370860a6205023bb1fd2612873d5ef2d56458cd4a0f440da56f8b3d0342ab8e754b9b2c1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf00e61f20c2fce206b79dfd5abeb10f1c1b006904844a8d505fe58d7db71a75c0235225bca3f641b368dffd7984e2e37026dffd8ffe87841972162222bc0be08e121fac75498fee4db6d5e2ae8b665b3857ae22f0f4b8e7453608f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2867d8883c3df3412a4a4c1bd1ee15f2fab6b460f116e1ed02e4147ecb9604dbcbe2e516fa2753afe2c11d269fb53e9f0d51d0d2d1b28de843c36f8635d8f7cc54cf078a8ed56e28a6dd33f39d4ab565751f436cba54af145faab4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7ce3e6eb241ab51840d32302b355dcc0809ac18eea4f34663231f22df5f7d810de9cf64405f617ad55a5a44ad25a93c9ccf46243d309dba09e2e5ce0e65774208117d7aedb8cd8a517c413e6b141313af3f247a0ed0dc1ce38a7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba30defd96beb9051a2f466cc90073ff14526808cdb5af84393ab33781ba40028421b523b79f5df16201ae37436fed5ef3b2a15c0242b5281f1c83b6fb3973d11077f42e0afaf96f1233aaf3634de8283cdb6fbd1fb79752dbadc3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf047b6989954a9347a7cdef9f62defe628b00de2a0c605457fdba14d0fc5f4db168a908e5ed76e5c04c845995047383d2849c854cc53c57b40f4a67febc55c536f83b3c24753681ea313e842c5701880bc829b6e822d0dda78cb46;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ef689af1eb5575ae24ce38d85a15c757685fcc812a5be417cdae06f55cab91d4633625a068f50ba6669c13b0708dcb50c1d6e92642ffe1ada99d47f2b4dbbf1f9c1e3839ede8e1e8d13f8541ec3055050b5338d9dfe098f586cb7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf3b42494b74b77073a8793c56731de14c92074e405033c38458c70742303f36ad11ed0de31c3dff2317eb6b9fb9408488f8c5be12dd30ae08c012b192b3bb3ccfb0d1d3bbcb61b031e951ce99e9d1b0586936261a972cbdf5c1573;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h577b6176f60cf65fe80e6ba98df66cb677c155ed2287627949e5652398336cbd344f4c666b31f9d791c3fd5bb21ee938ef08ec63de4433b703c9ae6871b6264ba673ef09b7391b8c22b9028dd1c630a0b59d356df775f5694935ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f98477efc3f72bae5bd073f98d8fc50a0cd47e2076f1cf3cb8474941be0ae7cd20856002149290e0efc84827a340a6578bda8922af6f93c063c1af834c31e9f600e691d1b0c690532c9c423863043af21e64931d70bd57e3a9379;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h133f58bd2175ef3ffeb825bcd6703bbe82e414d362d1ec9adf1499404c33c47a47aa3b708cacbdf5f1719cbee7e14a0f95481fb2da2733f6ee37d683f78f94fd27b218bcba84052db7bd2abcb899a5a3f206a00d070752672d77a8d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b441924ff2ed1a0c73b9f0426102af8147fd5f52d5a28a35d23f92c7d7d1a54f63e31ff18c5dfac6cce25dd53d43b3c2257cf2ab0fde850f4adcbc25f32c9ec60dc4f678bd7111ce44212132413301f135beee30e9b32a5afcff2e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9642f57fa9503777852d458afc3e0603f210ff8866035c34ebc5c5f5c9e37cf7da7eb9024f5d36895fd8bfb013277799c84b02a511dce07432c7f11f4c77a8588898507fb7e7adb09e91908cb944fc25d40514bdb489a93c452ce;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf146b87ec36274dc516b363381aaa216408188352afe078797a217481919f933a0df8bf0c3d7343039e38a23b4c84ffdf6fbc4ca7f9c8a6d329e121c719dcfc42e89e06b334131d3a1c7c2d00182c45c76fd6021c2b4a686dfb68;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h134264777ac78ffad180cbf6fc00ce1c05520b1f91fda25fad7f3c917335241c9f46628a9329707678e139aeab7e48d26266050616fd018933f86a637b4b252ac51a442286c85bca7a741ccb83fce666123753578ccab26c6453912;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1993ff7784aec1db38f8320c9a490d050caf5f08e5457f7218b1f0d32e293a252ad064a3454f23a1fc55788650b62895029e7d0b04d8f03da362477a896033f3dacb5b3ba073029b8b64cc076f437ba460690998bebe3759c472937;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54d62117bab45af17a1bfd1695e4fe9a138b31d53fc0c18f7844ad2f0d1f43ceb34072e76906dbb5456215c9bfd921cfd743e075ba5f6603dc02834bc1ba1ba3fb601149f59f028fd2602356eec59adc59d0183236a8a388332fa4;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b645010fd31865bd3936f1d70038badd3fabc36c0eebbf91972a169c658ef0ea452ba3d0dd03d94d2ad1f8adda8c6fe348f9b442ff29225cffcd64083f6bd56d8123269b5c2538a7e52cdaf37b5605c2ff6960087944c6780f4609;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb91d3ae1378a43163a04c8ac30257c9257751b8e2539baf066bd7da32d30e545862b3dcfc50f309380172b05c60200ad614f4cde19b74aab0e132e80545d189fb4c193b9c106672c4c1faaf74ac6a3f0be2d3c73a9a0245b82372;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8671829123b908ddb1f59d137ee53301a59d594a60810a5a3a7588a7f1639cadfab8bcb126b309f5846c464815d07eccc6d745fda9519a6591f69b661bda10f36be69fcac22987dcfa1b4d246ec4bf6346c5d0b9a1030f44c17d38;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1775e08301173cb823e3c955393fe8fca7fb4b5f06f11ef93a63ad603178db3f71af7d3a4faab0f7d47e5f94aced7533c44f3a4a477fbe7d4ae9b020e5d5907acd25761262d576841819f850213e8cd2ccf1c4616fe329f797ac44e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d29189f812718459e82c9c0ae7c7c12fcf2d88f55d0f995a6a5fdc0e13a3a72583e51f073b1dca496eeb62d8280e371da0b9a795ac0600be04ceb562b353b01f9a14e9b0adf1ddd2ffac54d64808244552566c46cbb9e0866f34a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f67ce9ab4cf33f085b3d4dfd7f4cbbf769c83f5936529f6b787aec1316f309ad3c8bb622730cb3d0bc868d7703ef5b4d8bf2d63aa68a4f7ad63f1286dc3b388debf8a5b0a79f3d6f3d3cf278dae753f975f04997b5b4f4f92f5cc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1e883a7732ec8fca5868d60ed6e2e88fd36f7a34abcbcfb01d71cb7b61250005d3082bb08d63a92d2b57ae19d088a0f807ce9df7aa6ee042ea06d924a893c80502ff9abda2e31e38e2e31b481a66b00014bd168947ba4bb9bd56f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107d86b0586e5dbd5329bd8aec848162e0154bc1cfe2a44586cc09a9e8dd505ad4816d1078a4cea3b4b1959b76c0c6dc9a4866f4946028822729fcf85daf2950461f6baa4a05c8961878b604f88f43fb34d42b849c7d4b0918050dd;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e2ea48dce39eb440f8e9b5de95e2eb8748b082ffd365f0096d16b19d49a66e4b1f3255e0c6f22f95122b65e2d405dcb058f8b5d9145efabef57de161ed2c120bef91b28314d5e47613a9a179130f12515e1545cbe78942655ca30;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a1c6ee6d0f5cc8e0e76e85d09adc6f9ed79043cbd753888aa7c2e8c3d1c4c2fc9b7c0c7deefb19cf7a0dde0a3108bd931649b4d0dd493049a125ff1132023c01f805596389de3666cb0c9ee8f2ea558adf92bb4fb0601015a869a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1566c33104a388f6136e3a5e73c2b649f3fe96f591292bc29a1586676a06de83475c12cda5fb4f830f60b65454ebf9dab57e2237c195d68dab854eb7c692a557948462a6e13a41469cad756c06dd9e8c3ead158a13f07a9e14ee84f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c14e8530d0960f430e82f2bd1c57f293b3f1a07523816ee9ae1c1e7f65804677e83dd24df41fb638bbc0feaf5fd81cb7b59ad817b4f2b78059c8b5ef0a2a933a3b94e5d197c52d226121a32b20541ce671907d62132f9903ff498e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13948cbc1574223e32bfebb11ba57d365cbf2e788a95de397eea7b520a735ac18063ec8499c35d517798de54f7eb1152d7bd65d09fb5e79c4c26d7f7c5771d291043c4e1413eb2f75792a7046d76a0cb7ccd26c21600be42c110d49;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fab0aaaf2343038d2606c17ca9eb02b48322dc2b711f9f4a1f7cc62ffe744f7f02a45d6858329a98cdd64f95bd29e1e16133ee115ca5ea441b0e0634a9c17d70607445cfbddef0f4d54e16f7148146dcd8bacd636b3c1fc6614994;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f55c543e2d2fd4e81d9877cd3dde0d68a3feb5cd5d440495aff5c418cb6e56b777562d5a13f08d7af3024a826c057f3d988e4924c37bfb58d951323b144a33775e0a5ed9f797b9509eeb4d837c7b76ddfc5598eb0ec4077964ac0f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2b302e7b0944eb1d8e5f9a59140808d79a2a68b73bf307f460fba3a4bcb8cd1a1c7467fa190e672f64a78ce7fd9495a2f4ff5f4d82f8ae139bf1634476ff4242d964787c33f623e5d235a62f608d5c9907b71045ea2bf14e0e0c10;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b0fe75e484a0d17df3a5da55378845771005e99c9410b196f9d6d2e2e833c0b59bc42e31db7a290677bcb336428077d206c0837954f5dd0597a7f1058b241c04c53f812e2fd2901742adce26ee1f1601da91e42799e9ffd45e621;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6534339df83729e60e7d3de15fe0e993090efa36341a3d3cc6a26e7c8fa9c604bcba00b432db31e839d767ceb2711fb5d5f73e4d0241882f18b1dca27063cfdee847a734302dcb5a7ca137da0ee8ea7040e1314d7fc5b66ea0fb7f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93812046015c1ef6b3556d839777581261f41095f773496b2d842fceaf98d891d404f033581fcd8cc729209adb564794579c265ecc88a20d27d7475fef7718633a3829999b0e190b3e248480a2b649c677d967f6baacea6ebc0923;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8b401ac0bb6be22eaaefcbaf58e5fc6ce4d018fdf20aecabafb4b13b8891e207e9bbfe8796bd601179d4b2a415f3e2cc4577719514c7e6c037926bc48a14ffc6698f4164f5203216ae713220f514412dbabda9cf8a13edab0170f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19cb8d39a8fa13168a571191aeeaec59a8ab3a86d3e1930c3b4c74b3bcd50e7040cbf552d2add9662ee0ac6db06a4fbba4778d9476eb83a7455120577624db6fec951f6141f790562da64d1adcc4caf73c48afa994beb381005d739;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb8d3775bca8203b971bc7f8bf1f730e41b031011bc7c52473464d412262f887a325318453e7f7388164d13ff35161eaf2640baac759615dc6c0964678468b25c048442d140d5ca94f3bdb4ee3439025cf27eb018b4220f0a50e02;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d152a92d58541672ce10870066774cb7c12170a2520901fb1c15d62b2d39cf85dff154a8ee5dc8b20242b294d26f4d2cb227c88f9f4f3eaf4611106dd0ce487d11ff7c47b6a87d79aa263dac457a94cb1dbe73358fcfa0c346dc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h187453a8e9404e649a7c574006685daa1802635cb17f84d1758a8b5ec4d32c1b2019cf4bb42d95da515a6e52cf2a67ce311f6ca9c41c86f367e62a233e67f63f22e3eff7e67a2db9ba5620513e13177907082f626affd0d9a3831fc;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164d99de6251ff28d869e65a291eb27564a4caae7d4f52cd9f562d351af6b569ca4e123f1909aec4dc22f99bf391ae1d6de5653b407cb82735baf7eccae440b7635ca3f70eaafc744f7630bccc42e04cdd9438bdb290acfbbf4c2a0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7761b91cf08d07acb672b84387c9d92a56f965545c16201660671bf879e207162e96cecbe4faac25abd69b911165c90646a48de2fa66fc28914beec10a21ee3fec465cbb7013ab7e21ddd6acedcea685a12f2b4a3fcfbcbc0dd531;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h95c97dc26edafd2d63a405f1f9c09a337d3e5fdcb5d80fb2dc204e7b21dfa044ccad66b80dc78a8c600ab5258cc063957833a38a0ea535d652c6553d778835bc54848d18664bf6014e4316a1503a6dbe4455368a415752e8a6462e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12d5422dc320b5c86f3f3cdfe84c5aad909052826730fbd2ed3a19e8369e6fc0c71edfc1d4bebac9ebe4463240996ac93f91bc1a25637e3adf17af64eeb05df3cced057882a77f557c67047a281b46890c3f5f5f090dd0f1d09aa41;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h140504c75789f0151ad49909ecca30df4aca84ce6d74a49d13544bfcbdc991b95b46640d0c13b77bb94bd356150e64ab57c7c2551a97fcf432992fb0fa8e93b8ad4a3918116b42d831ca2a0338d0f1f7a5b35388b1802c6ce0877ff;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13597107a45d080590a00e1aac7bf16f2a8d6cc2dc14112e4c566bcb221279b36869609f278917e93454d580feb676dd4facb70df59ee73710131e93bcdcb340e498859b20629533cd0aa3407d9057c50b5d83228139f4023df5006;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84ff5b8ecc1add037f9a2ecdf231dfcba5ac6771c795668e1f1fe7dbe366980f95ba6a9bf97d0e9f74af625336ecc753d563ab9db872b99fa82169e82ed1a59d03b3a165f63f04866f6393c5e4bcc933a819dc2f937f693bdaf931;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1ef29dad8bd72ca3c8fcc190aca4de6a1af0e9bfcbaebeebc482c9bdb2ccd08b1cd5bb8ce89404838de0b32c75dd5bb6ec2189cbad82e9452fb6787a727ac2812a01f53de48bcb8cae46359c6b074971513be85a9bea223236796;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18fc9925f72ee1d55381d479ad8b9812226e98e96bb0d8be4a1dc68eb6911e3d23aa2ae27a50d41e60bf36f8a4768b72d79a3955fe76c5fe36c2eebcd57e39ae00149f353387ebfb4619a3ebeff7e6c7ba88601a2729759dab7a0af;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6fb1b0479d89847290a3aea356566e444f949b802df8217bcf355d16d780129b14de088e9df8ac5ad555a3d438e533768a1913f6aeef8fed8811bcfe44ebcb59be17b20f0dd0484fc0e4500b55712b2c56cf8ae3f91efb2811944;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e1c38c465937c816753f5446473d8d56a0e78a7775931809dc193df878b768b53dc779c7da3bde938677f7d72976fc205692d3230216f6cef34e9ff9292c7242bcd3a3350e63861f016630f367868b1fde2470a8ec3978d99d0a6;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3641af9b3a056bd598f79d2db1c5d94fd6076c9687cbd6c0da70eff05ff86b6a8251fb931c5645001fab9c171214119b85af72b515592cf1c98f208f75679c2d8d1dbab24b65638cdfb78361231fd44247b217629a9841801811c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10c72f15216f883e4825570c52b9f9be6bf84624c98f7735e038a966bcb1de2bb395cc0da74de3aa181ec038716f2f2cb8a3b7e4e3f43b4cbae99e8613bfe637dd887d78176c6c67d18cc48d02965bcada1a02668107321c665a8;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9bf2e541c4a2718725b8d34a08248d0676c6ef490c1f2151c74e7ada6d48dd5f9e7ed4b32e68f7f3a5d4dab08f3f7bd3117e57c6f0974bea40073899e1268dd7c9e4130328faed14cf169eea52a7c69e558daaf5e4ea60ca87bbcb;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h194e7d8771ab0384a313dcea1433b4d9dd501e863c829e5b640de92c5349952634a8248b55ec8f1272ab4943816c3b8dce034fa7774b7086db4c3be7cdbb674fd1b1e25db4c88d551fa70dea6725524e5b40bc1379ee552fce0bb04;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1cc4b06c083db8f1c00a1b0174ccd0dfa076d78733a36c59074b6c2b9ee40af6b4ff733eb5c17de515cd842550522e9790fabf841e853cd9784d4de88ecd62d6cb522b58a6dab078b104c48241308810643389a1047fec2a4fa8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ea0903df0cdeb4dceed250cc1a8544886dfbb4284d793d9e43b9d658d1c93a4f1f9f83eaa0d1d85bc0bd56b2c997723b952c0a060b2b3375c875ccd4af1622c9cb36636bfb4d7b70c3550ca48c0728b430b45ece5b1b7467c27e9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb66d57ad38ed7093e2c776927da40c60ab7951fdf1ccfaab4bf788e508387a303326caad2996e16db6f412df13e3253eb17edcfe045455bd3e44062aa5d4cc43a7f52599f7ec5179a7ccbe92cdaee352b9434948ca86e221dcb6db;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce5eaaa2b7ea5c6af3ecab7832b70ec3ac39fb829e842c477a9789a129c936fdf9680eee008696df7fe7eaae272495f4f33fedb8daf9f957912f8619fd802c480b6a4a7cc0d2b7b14dfc326b50113c8530e3b66067daefb2deaf99;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e925dcbc14cd518ab91c48dbcd1faee479e5ab58ebfdb0764ced16e14b31b5a6decefd21d460981a94586eb3b901cf2012ed1d0161674da11f2e91246ccec508b6ee76b1593b8eb88788a83fad9b04e4b44c6a955f450f15afc770;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha5393da0ae86f181c902146837cc6db7ce14d02dff3cc3c8dc2260188f09c43ec13d4fce0beb7c2344f0f7aa0ab893473357950aa28c92918aa2c003756f13965c0b3c35961eb893fd4074717847ee87154a3f0bd4954ff389169a;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6be603f5085fa493ac7f2127970149b2672dafcb4eac8d4247c0114dbee18a813536d60c848684873ceead8a4f023a90fe26417b01c49c6d95b486d832437ec3bdb68c283d35e511eacc1c17c1295be8fe0a0d1a4767f6771f9032;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1594da3257ac8632fbc48a322354ddd4a8d00661d9423ff3647a117e3ef82a1e1b6ed7a07ecfce22b4ff0e560f46109e9b14917c0aea914b9156445e6df8f451aab7955095eaa9ac433fedd5242e2862dc5633ef8516b6bcb8b60aa;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1919a66b282fc490a7eb24d583521b59581b52e09d198a61af65b28ec5cc0a17e014d8dc580eaccd412efc025555677e740ecdd35a7466508e174a04a769891896993792038d520028155abb0c5638bf72873ff11426d18ecaa97;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f75f1d2a4e7be7c429626fc7949f6e7de8261a862a8da35fe3c60231dea2435bb8d1e93810dffaae049e92d81316dc1fab479316941cbf5dbcf07390b9fc0cf3c2d458206d8487e0baf0692522331eb66b4c76218ce53fa65894e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h346a8fdcfe7a0d59bc63ad2240d12cd77658f864791975a83a2b9a904ac28fb04dfc7eab11b705a28c2782251d3b5796418c3dd4de55d6cab29e5959faed809021cfaa686523321c0994a014522a770a4e3e3d14f8b59f2a256172;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9f46d732db8687b14408ce9e84f7bbf78b35129ce4f2cbed0feefac84e7ea51194b2a09c00a3211ab9eb54a18424dd605956e27c9ef57100242d1b8bb985bc02cec37139c193acd4cef7c04888a37c9fa4629bc329687efa276cf;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5b4dadb7b8f87396c152ff7be824259134072eb3d1180f9d8786c3cb90fdaa1342cf8493d6d46df77110ea6f4f58c590312b7a80e8ac272c5849612a3709b57aca57f5c7aa3fea319aebf9a6c993ce9ca7e493c7c0c651315b6f9;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1152d75bad58cd89de6b13bdc3f0c313760cd9ee2994ff98c2268b44d1a6d6d8a4f95b285bf5d7c5d402110ecba2caf96a1725c01d9e3fadc33f39c2e6c009da7c7b4f7b789ab61813bd4c0f10fb482828ed4c8aa8c7a6eb6be425d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5557f819ee59aeda653b501e0db7c3987765b4ca54c374a95b78890968570e5ed9783d98162ac210be0dd968642256f68b96ad10216495ae9691dfa06aa8b43196de673595547337bd2b79f18153e61eb899d88bd332000a69d82c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9e4c08c2fb6cefccbdb85272d3e2c52cffa0b6c1e164acc19092332bbe0ceaf991f87d6601ba223fa2f81b774001363649fe68fbfd7fae12746abdb1a94c2129def7a7bc461325df122110cc21ade73d286c3e9f53af4de2508f11;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68cda784b5bc0f1ee848c27ebbdbc98048884ca27e15af275c91aff1151bb58d97b7a0e689f77b88c201598eb7ec0c3feafaeee94a6d5a89484bda90d29b751c07b2b321c5750a4c1e4be91003c3bcc3d34a76411790207b09d3b3;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffa58e1909fd4232badeb3d60b346338c5a4b821c2807027a3e2d04d4e6ea75d9b68dbc5194029e3e900af88628668d35ea206dde837084018dced9b693da2026b7ea8ad79bf559d76bb45cf0ae716b7327453cb491ce1d385625d;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1389e78d5bd00510fdc9c3434dd9322a3c39a84c1c8411ad0a431c64b4317287ef031823d9fe33de43f20d74eb63de3e6a89cb197f944b4655022b2ac031c6b68d0f0b017258b409e6d3438265439b00348bf7717ab653e9409eaf1;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h35b73084f618df0324b7824b36a168cecdd266d40180d7e6bfde5b12197dae0a89f1340b1b99706cd86f02b896b162aab8f63aa53d47efcd978aad43f440d93a5fbb89fe0abd8cfa69673f8d7a9c06a84cd78f219b011956e14300;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he12fa08fb09fef08e62e8cb2bd6dc71d49c4ad146b6949baa8a0f44294c3923c3ce45b466f7ef2bf54a58b1319dc0da19ccb3250b79cd8f821c94f4dd88c2696179663c21f2aafd386f8d0b61649449b00e6a3400549eb8307206f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f9cf6bd6ff2eff479ac52883396a66fd5c7007172c76240393b18a0a40fff8567341e918364ede3667f7ee8998e4c8151bb0bf852d21151739a2663f683d61a82522355031ab3aefa33a5c9c28c4fbc23cfc4323a90020135944b;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f0c63f05c30c03c8cc01f73a538303aa5f843bbd08e38faaa19b9e54f9e419c414a19388c55e392a65372ede3b8f4feedd99c612457eb613468cbb62f8b848c8abfb3e55016045bafa72a2068c444f4a2d2ee9407187e5439f214;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1564980828855e7f911ca7dda8ac1947be639f60b68013e73517c509209cf80214a3f1d804d4a5b5851d55c94b2f1030f9488d845bbe475317a955030aa1528dc4c9cb01808bea217ff488d72f6d76780a7fe4d08b03cb366316ff2;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16becd066f7997b1f823b39b06d57456a86127445e785c0964fea704801718b981922fd3d8ab28c4dc954af01d0b09edf1d6505ea79306848f223e780ced9863ee0093e965d8ae04ae7ecaf4b6edf025270c6601d77ec62af6b7fd5;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33c28fe5e39d5100884ec8986140da1ecc3ede3a88381b7013080cbac92e24ea817812efce2a9f2e9044a9f80a15d1ba4fdf30fc339bb3f9b36bd0eb96898eceec2da44c87fc1a9cb0ae00a0d432c34474a59e7a12fdf73cb3e449;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbab438128ca2d24335df52188f75ee70ae2d104adf5666cb0069a925b8395306a24e15908c2e43af076e1a7a3ceb298615efd7d32b3172d0f15fc3ce36744654431e0e5207b7a6990d4f522b21a56b61e101103fdec234dd55af8f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b74eba69e449f5645edf1f3066b7c6835dcc203cc7560e62fecdad46ddb2133cbfe7ff72e64331a12b2b6f556cc72f79cc1c1e4fed18f59d028390b7c31fd2cff899cfe5216d9d82ae047c979302ddf53e990d4860ade56fe38e5c;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he7d5a3941bcfb3831a75049c626224dbc4f0556f5629ba3652d66407eed8791795027869698b538d34b95aca7cc2ddd2e03622bef62f76c01a8b4ea916fdf8e257c8da3e0071f291303a0cdd718a67bc382896b0327f0a6261928f;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70f318459e1447b35eb261c71466e8980cd04e341cf82985c5899eb56b3a04fd2e126e905605a5ea6fe065ed00ca30149d8eca6e4ba4e0f574abeb8f2efaadfac72efe87ea11924eaa1ce9c5ee165e10a53df6b77eb12e3b45ee53;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca6f05f89978d79c701629de780b858389cee8a121ce4f9c2d1a0a5ee86a64fa0adaf7e7f97a28f3bcdb16571b338780c40370583ce82e4eee70838f671e0e59ba18d0651d37946e372bceba315335429fa32dcda520e010ff4781;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a50118940bf98c536f6914e2a80f57454cc2b6d09168dc7cf77ecbb2c4b6d342657a74dde70e705868ca5c28b1c7674b82d87e2f92dd3bd2013500101743ddb7176030c90254e0312e3c8bc422229a553951e62776bdfd7356eae;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92d929ebfab2d0905e807025e599c12534769af040eb069dc1f056ad19d9645b9fb975d48ac08c4b4c9d312c075259079f4d517e645f3133fe47c2ae03cdf6ac3d2929fddb475a16c4b902b29ffd87a9db67307a4e4aaced867d52;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f78a80ad2e6c026085e4f3386086f5ac6062608d4d6416f37ae8e6fc3280287619b4e69eeff4703b1da8e29e0b8c22bea8b2d58295ecaf9e3dba5c08b86c432f9a5b74585e915d7298e3c67f6bb5962ffd190925680f4d93d9e17e;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e9299dc1d129551dd258e75b9a4a7641f8d65bbbfd011226035d2df3864a7cb9ba325a4ea174bd7960a651a886083f80812b5a96769efef6cd7ba438bef5f8f6a66914d5641c7a951d0495c6fc89223af9e3c0ed3aca3f5a709e7;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171e6876363ecd9d1dadac1ba5e7eb61c0f301cdd26622bb28522a489227ae8150ef1b29c7990cdb56093d29b4be4f2ef88572873bca297b306575a0459329213e8bed9afdf5266dc36850571fe534febafc90004b464b5073d4616;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7a3dfe3f06600cedd6ff451e6a9085b54216c18e222bec71930b4fd7a241a54e20ceeb952250009fec10fc168509a6d322ad3f3fac1ff83f432125fb5f59f3062d7b41ecf2bf48933b9fa5da1d3f0c016e60032e9efb11713fde0;
        #1
        {src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6870ba2355a8eba2c8e42ae58cc65f09a63d22913a87a8cea556a3e867fc91041526318d03a2f736408ab31d76eff3ebef57d945b54fc09b6fe83ad793d3ce9edf5953235fe5d9e9563c74508998c362cd76b364373c733ee2d77;
        #1
        $finish();
    end
endmodule
