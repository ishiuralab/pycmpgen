module testbench();
    reg [24:0] src0;
    reg [24:0] src1;
    reg [24:0] src2;
    reg [24:0] src3;
    reg [24:0] src4;
    reg [24:0] src5;
    reg [24:0] src6;
    reg [24:0] src7;
    reg [24:0] src8;
    reg [24:0] src9;
    reg [24:0] src10;
    reg [24:0] src11;
    reg [24:0] src12;
    reg [24:0] src13;
    reg [24:0] src14;
    reg [24:0] src15;
    reg [24:0] src16;
    reg [24:0] src17;
    reg [24:0] src18;
    reg [24:0] src19;
    reg [24:0] src20;
    reg [24:0] src21;
    reg [24:0] src22;
    reg [24:0] src23;
    reg [24:0] src24;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [29:0] srcsum;
    wire [29:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1509d1e208b45adef7464f6c09f6f4617a2394edd3d49060da5067fd8c1136d3532b17102c8fba10eb0cdd5d1c9981d6c1f82bc82fb4e9fba4d8876aefa0e8170726349b7f6b8ef311be286216ea8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1096b7a5f0e489f1cf58f2f59d7df766f98aa609b6dc7231beb7b6f3c1cc0cd6e9f0006e6fbe15f1e509a260393e78a2ad38d27589207ececa456399c1b140ca0e55b927b242c6b5a5ed1a09dc97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197aff95e3d7cb560a9ae844705162a47ef8685a2cb6a1318bc1146cb3241dccce0886c30f7d5479eee9e6a9367f775ede820b2879be635f75b97949b70ce42ee6b43f17054f8b3ac9ee71d6031b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h431d9ab482017e7e419338ba50a6877cfe36ed8efe2dff1278a7e67fc19a1f8d0c86abfe768b75aa997d94161500cbfac1aa9b5403640ac80a6b96e2c998aa2739d2d3a7499785cfed039231656c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h36f6a630b0ec61f752bd2f70cd5638897ecddb18994c5322c2d894e59ffd082ec73beff4c2b6b07e777e77ddd2d4cba011b5f2478933d70343638a1a313407794d5543eea94b90b29682de0c7b97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b5d63fdf613a887ae7be94d65f0951d2cd582ffc45425c61cc7a8a873dc2892cf73daebc998f1232712e0a35eb61d925d258bdb84d0517a37cf5b73cf10aa53829466a0c4768d7d099bf9d98127;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf9719906473416734958c979e664fbde1f642fc940fa21dcfe3d2efb4bc9ff1f6a741d1e31ead9517db924b6d7e6b212698bf40f106eef3ce483297ed56903c17c28a1a93176cf40b9c1dabe0df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0805ffe9afe4e49fe6bcdefcf7c7f332c2fe2b341ba481926c7e79d2e32d024d35f33c77eacf4cbe6ee1829484eead44b9df56cf991c3dcff99c54241f0fab928a8878909676ab8ce48e8b54fde;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f357410150cd5b3df94f418130b8fa63dca251b9df029e4d26484924a47b343e3d2436004a404d37d81519dd48531f68718d3d846e11967ff7198ed5625f17352b63c3a72b86fcfa71a2ba01a62e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he150ad60c0ae3a231f7fb480519b6e68aa6a63e793e6345b4a87a48917c27b2b2e2533113d8fb8d0abccae49a1513630c6a151f60db707417c5c8be68327545be49105f7ee44a2440b87bb66c7d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4fd28b328babfb098bc92c1fa2920915df5b862cc5afbe3274dc75523b84a7add4c522a86f397774b801b55fa8f2ca7b31b8b1ae41cd1d33a0e2604768b8c3535e81b1e4628092699bb165c023;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a86b4f9bb726c065b08d6d24d311005c10bbda3f8530b48eed98502e5a5d9f0fec30efc38bdca510872da9ecf945eb1fbf04680c17ebb3383990c135e12463b572ea7bd3b92fe8ffa27ac90b46b2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb688b061f217f49073d74b208a23d790c9fb45403a249e0d3ee884810a60a975904707d288a85ce078ebac1eeb35d1977dd0865d19df62deb38e65ebd957475258e80d3dd8def735d586a69102a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1186fae9356deb99d852a6a11ef8204d4fbc78cf3a6ae7d0c1e79c68d54a0ccc4f6eedf29761a21d5c6d28b1249cd5f3a20d3c005bc96beccf38dfdf3380df0a4a3e16ff6463241ac144a01c63d97;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41c1cdcac4b9276ecb0b993c724cbb82bc26f0ba0c82f9a0028e85ec0d74e9c3bfcb49ecd975794467a699b2917b156f812d49aa87b0ff7bdd5f3752742d743e1ad590fb9322d53661e71f054ef6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10717bbf340bb5d5c02f0c7ea4d9c2f3b78da859f057f64c967cdc6951da7f01acf6e1865b6b758879f30eae5576729c870423109d0d8009f63e3623b2f57d3cc00be36df5ed68672f19431c1113b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26d368e3c32dea4a14660c45cc214e663b41d856c468f27162af712091e8773fcc40427b3a4fd8852e07bb4e6c54bfc0b2db7c1c6de26e2e5087d32ba4bdd860dd9cf5c0a44aee7b3aaebedd03ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdac07a5558fa437bbc3ed903f4358f4fdbb612949e523264a21aaf178d70365a24c1e7df5ea82b081a714248e74499dce58dd08c1d0c2e6733347aaf395fc8de982c20b5f3c8cf028924c3ef70b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5eea7051d0fe15c1912d2592b37b05d7d90639bc9ca006fc655e6444cc5e22d946dde8e78cc700f682aeed60ce29f51b304bc45c6db21297687e9592fdf6d86a29bc36e123cb5b59cb731d76cfd8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62eca80592dc9bcea19fc60acba8353f3bcd903cb33e5ed9c4a43d5c2e5d18f05271101e00b04095a25a51d7a43835c74b572606118b251115c014c2490d72288bbeee7b9a64782359ea5b0da8ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df63e80a4a3a15ad18ff65a86e44c9b849c2886b91a95213bf4d6604d2347638d7e16432432f613b33254902a0e175bb8123100b4131480d99d5b64b9dab866cabbedff59a27ac43a1175e6d4762;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4651d46fe101053b9c59cf5098de9e0083f90cea861152989d1f1f1bc9fad6e76a17a0e61f94e94042e88ebd0434148f467d37fa94302a5713e0e66d67135578118283607fa9cf314b8e4bf2735;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h58b5c67346f99d5f38898652ce7a8585df47871ec3f6b5ef85a1005581a8dda77c5e7cd148aff5e1d45bb49ba28d6fcf0496b9322b7b1720a84a044ad61b8e4d6ee726a1ffbaa32218b7cfb7df34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha72d0ca2ca368cef7b989a16516dfb7b9873c9e733a1560b8bbc40a724e03f846b93599da11cc32ec4f4b58c1746ae4a2376b663dad4bacfb973249ab568596f335ce335c4609d2808ee7fababe0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e412bf1a059d860ccd0ca15035966d9cbd77f2e4c7050f405a552e9a4bdcdc17e69769dacc4de4591d563ca077ec59fbfe39971e6c57c9b4750ea7d17a977554b33fd8108ef4cfe92f768cb621c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c31f69a895309afebc03b4d22587658b32b9ae7400bb5d32c787ece21a447c02a4f9bb87949a9617591393ccc761a777f1085863fefb095fe40d2d098f9c0d621dbe42b9fd5adee6c22fddc23ea2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa240a1efdadd2808c083cc0e541ca4655c55f76f531976767249825d948b351c19dada87e06d0f06d12ecec623236c8ce8b380ce9e9d1d4e1080f0967bd607aa624964158f3d7f75b93b57c3f5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11583e561ac4c275bf55725c9790b2c522e971e435a2a72da6057a2d3b36eb7d89b1394b5dc7e095add3316c8c71bc9bd3e2aa5c0e41828fd4d62f72b6b8ee8c816c1db83d7e203e6449270a68b33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bcc0371c9796a88d2e96e7f147d3c5ac029b89076c049d9f76c59ae9e86a429548f1776139bce10ca5e36c7ce6a887788d2b44d744fd130716dcdc804c113cbca362570da668b400896901c67ce8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hadd84d2160d867068f016f4f6fb40f67a2284e8c02b1fa581ef25b281f7ad43cc9edbb4fd5ef0f57d9f858cdbfff373e77a72eea06e46cea992e1c08175e3eae1c8e37bd8f91be5b9f0eb187186d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1877807ca480264d0b2cc0cf8a031abd301225ef9a9e350fd9ee5024e8392377de02854adf7404ab2ade136b46bfc729bf3401b9fdfca765d6615e3fff21ed28b3f5b61570bb982251678f52c463f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ed77aecae5f412647452cd8f8306498319b619fc000d32ffe3ec4701ff89ce1c51c84e4c7cb08c94645a584ac26ad3df706ce0d87bf467f9cc7cc331351dd09ab7c03852d4fc8e1716ce253b8d61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc531561fa0a6a99f528b5a53aca7323bf15123e172fc2265b263dd8d828f65d72f1c0a3d0ce5b290bcc3c7174528957724ac8938d6ed194f58f964e03ec9a8f709a2ad11a36c03d6d5bf53099161;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a2197a7d76866604e2f60aed03605d1d18a3ee9e2e4ecc91f6e329310d4fb429b715c54f3f49b97d6c29d009631d6504798e08211653a3a39ccb3a24b75623dc4f0db7aeee3cbc712aacbaf54d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11e1ceb255da53afe24ce0b6a36030edc2125255e91a16b34ba37cababda07a31abc1c9801397986f9c4f19a74ea910d2d2e2564a9882441d190be0b1daed170f46785149048d6d4939730a955f2f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1414b7906562edaf3972af47cf73e267a2a33d31d2c1053fd875896ef333f0be177a20a1eb3b79618eb7a6a902bdbf1b37b4646664955afb7cf029149bca10af6e221fab48ec16ee4099480b9433d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50221d61ea30afcc56962161271255349f87a61244a768de61d861fe1e1b19d490338f15d77c048dcf745cfb42e99c337a481e5c01e6c7405a6480daba6452b638d5fda28dfae04966e0d7f95073;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171c345e7f93ed43a8fc2e66b79ae2aff7789952a8010ed39049c0b75e99f376bc1c30e9def98554a21acf20f7d967a2b2d37a6c50b070d2a38de16f881480195fdc59663042677385b5b98784d3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec5971b5ed1a0e32a73d388baee874825182f12f12b047593d42aa75f0aa0fa335659053070d1f24c4e4579685d5cd36a12898dee7aba42ceb0e50da5d5053cecfb5375c656275a4e54a7353f2e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6469fb0dab26eea00a8ebbf8cd98dd3bcbfe8ee3d74275f66dc33b41b1065c7f90606016b599c7f89f9fc024c0ebeac2afb5def7d5cc9dcdeb2449c8d0d3f5a82dd9aff12aa6c8742c5f0662bdc9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dfbfa6ca0f0b54c55f18ee53d1bdb554bef0c39cdf027a59d60ddbf8bfdfc41ea30c37443b5a0e177632640942d3c5935e97aabeecbba009b0e75225ce4e11b807d21941bcff1b98bf509ad18582;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2013339b1b32c099fb8f9dac9b6705c31173b9f7368b1170c9ec2cd482bdeba893573cbe8114559b39444776ae8b1296ba2d3fc5a8c5bbe5e5d4f3fa3df4efed6462a9eb42337ce341ab841396ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a788bcfa0becbad7e264d97d0b04686e93297ac468f0390924e73a7016b7513c24f7cd2cedc34e8820823222bf2ffdbeba5a35d10201bbb3e3586432f3618b8c13de80ff997f70f5efd9b46ac14;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1b05ffe3d226ebb7731671f8aeadbdc2ba1405e78231933deac94559a5d62430bb8c56510e2b15b4927ab0b256ef324497d8c1447db248c485581019e046434b6cae699845191020b36cce60a34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e997b10a1b8cbc1614fb94489e6b6ec9ed712900f326c9d18e7e5f51fd5303a9f150751346cdb332f772fbfd59ba5324f940a18d5900473acbc83bdbe4903b0db81086b0272bd27ff245bd927541;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c6f103f057775404d13a26b6faef816a4cd724817fb730be1698d8227d3d916bc0dc1d8572b68b01dbdb842b71056a560880de140385e5ee9130290b2a7fc2a1aae1aa23b77a561470d30a53c75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hefab8ebea0df5c5b1c31cd44c69d328ec16b5c6fd36f76a70ab8fc09539b65c38f439e282b25930199a56f867a4da6f3d57091a9111a126a4ecee841c6c8d3ae128a72b2abd1a1069998ea11f6c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57398bf6491c242abbcb38d474df449f6ca7a5af8b537f61e51285420b9011c1a76605eaf888dd5e720d59af4e734c7492afa7a8bc8100775b4ff06c413c24bad693c2af28100e48e7030e750adc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e132640b8948abcfd5078e1e66248deaf7ef0f6047c131407faa0fe563fb63573f881b996c34ee5f8a6a97a74f1ef35e03ccb9d4fbd2402c7371a49b1514b3ffa3fc3cf146cf3cc2b20676f8dc0c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1cbdd758715f93dc9a73db88bae813f61f78b91ffe7b4867a323208a18ea07afa79f3c384b7a130db534a53e85f7e5f576f1d1a133e836ece065e2afb24d3a7bbf3bc5e7bcd3e44ef1d8ec88fd0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0aefd7c78ba9316af6f62f433f93455f3947acd846ac9b7f9dfa23e4a03432e851991480a284fa23cd62d12b3539c229680f610e5c1cb2429285c0dde838c2cf5c0f31a74683938045f0cb626e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dae975ff0af4bf2276dc3395d1cc5abd52e2c0c02d869cb92c4bde8a0af31e49fa896c66d59c3dbb9788ad9057db4331c4aedff6829a8238951f4ea0aa60ee24ad9427dbd3ce2ad376319d077d7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d88c5b74e8664b32a869d71b422f1c2e5ffeab300a339aac61f09bf77f55bf85b56335324d205891e1b359a9e060a72e42a953c3a7ecd0ccb3d93685acbb011bd55b016f1474722eb33c94b9e51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3d806996bed81172e695640258948bec786a92a7ab5400f995a5a671946b162fb7d174dbfeaad98d23056fd6f6f811b5c245152d106989da433a62b3d0ce15c72ba18e3e1b229c45a05b6d564c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hddf77db54dcb9650dabe2144eccdcb012873c06ee47111c286eeae829af2045140e3a67a2ea1d3f05170dc04ab45af56a7c8d87e3910d586dff8ff1e9071982e35719f1e0c951905569346c0b1f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bf4f7011bb43b73765a82bb9233b6d40fa4fe2b3e4f7202f0f5c19129c70ac51e97895c458d958b3155391797d7e20e6b8a11cb82710f3d81e4d0629d1380779b7f89c28dc3ed5cfec77f781b48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc32ca5193a19a06e33f8b428cf7099c5b955102c9ca595a5469d87c9c86899d4cca35b58298629173ac603aa22e647375071ab5e69471d1fd1795c1f1064cdedd5e944e69fc0d28f5b19cb8939c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8184106e64abaa7c0c43c6b1fe6f3d7180b617e37d07a5937b6ed36cd7bd7edab98adb38a4682555aa5af4ad2697c2cf42ca2f30d11bd05e02da5feea440c24f79c659975029e399eb31aaa89179;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18858c859249559eb07668492ea2d8c9a3fe2f044ce7a217d1e3ab32d1a4db656bd52dc3124ce0eee0c5faa31ad4c707fab770b7b7446b60661b719234428e2c2870d7a4a0456de0319da2c66edf0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d3cc8035f7a6e5fc8a9aad881b66f9dbfdeeb1f7beec97714f22deea06b3c562999afe8638ca49468b6eb1bcf70fb2df5fe4b2af7db1b8ffd27f1ff4553c101968b76b62620fac9d16369fbf358;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13bfb7e4d882160f98fd340df43e8158729f41c89c6f3eeb73ed39f6bb66cb79426062520e84394918f345bbcf25efe2e9824cebc777974470ceb5c224e4b3529ee08e107e46b72b6b60aa140248f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f9228cb2064f127b371884f278a48a8b3afd7ce0c22bd0f666ffbb466e49a75dd3ba45b7cee097e92c4b79c090a51e4b895f04b251f053a7bddb265098e8d5f9298d3d158c6b2bf68bde5454244;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12fcfc564b045d5f162b6ab6fc356dfc14e870e8e8779c2719efe7fd24447d6861fa13b09c7ad2b0501b01b8461de7ec0b5d1146f997dd397128b18d7825062619b86a1cb42f43b106b8344f27a2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fd06f8db86b5c808709c7cc45dbfb9ce796bf99f339035a60662b16b5f2bc648125aa2e98c547486cf6b1351173f7c7a8138f99fca3d31f43dd73e8e8da30334bc3b4c4a835c5e311332158f3be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f47d7ae64ccd1516f428391bc6bed090ec0aa71367b1dc5a88d155bb76abf7af126d687178a2a7f7d7e6c48194f604d80840b78f744b45f19d0366effee6117f71df8743dd39d0a2850fe6626f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha4850963e5672da38f7f15b4d4d069142e60902e78653d02b051ebbdfebccd811b0ad0ace16a7314c1c517bda5c50d080e8406d56709af05be82cfd1f3d163e8bfa35981cf7ad85e1a8e0fe26c77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc07e83d680286579da2443da8ee46b815a0feb8e01e815fef0cbadbe39175979f5325e8fe5392fd9b43792fab718d6b3f9e5fac440e500a7136b71cc0d7c2ee3f1d37cadbd86b801f19dbe269634;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3bf5848955cc429959fdad6c017ddc5a38851f5cee5b15d916543a05b9d49bcabab5fb4de166eeb7b3d24543a9c4899e4bffebb1956b348e36c83dc1213690f96cba9395d4de56d7ad581d966c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cebf72210eab86a0ce15b63df401b797c51c53502bbf596d096ae419e4e5159866d393d53aa82422b2010cd8d49d6f340db54fa9df290cea0e62902ee007c6f36bf0477765ecacdf0cf8b010b32e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86e7b015d6e97a7e0b2d4c7c0af4869810b1f70d8053ef798ac447c6352da95e541ccab8c366d5bf0365de21b3866008d9b1ef28921314b210506e8005ca5d3f9ea601a5be63df8836ddfbeecbc6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d952c7a89c9dfe04cc02587bc7ff10fbee34ade634abcf8f64e949fe79bfad7411cd95bb24e1466818c07113188d42d09b82970b67e9a6411cdab3f70198b9a49be56c6685ed51f486a06108ff34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea673ec736e6cebf3b4192483a2f6315843e8c739196fd34c55b9f5d3b843d8bb5533d20bfee4f69766c7c661fe63da5690b7d4b5715fd30cf9e42c1726ea8b9d6feb9729b394e6316278ee8688e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6fd2aff1e25211231f80a00ff29ac17e8399c321407c2fc6b91b0712c8d01a573e87cc4ee87b3b8d9ad2d4dbbeb0539aa7d7c58c467e9867786b95c765a1a0f1ca04e687b6092dfae0b3ec50767;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1648d530c9d93c78962c7eac82cf624aa67f60cec44253f9ec429ea749998beadde7a0f007cd798fd2970aa182a744782680980bc33ee0a06fd6b8331cbfe2f538156d6e3d42d76adf3d4765b0856;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde416758829b212cafd64822de4d0933ee90f82f8d893732d5c04eeb59799fa5ec323fb159ad93b1b6ae06d16a522cee6642ae7ee537b37c839befac5153389caec29f7002973c152856c0fde3e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bcb8e6e7f4caf9f744f2f85029a72a0a48941498ac0a556c9be99b9808d43b1b24972fb100fdd6edc265994cf7862113e9e5b09ced116416ff5d771c7ad24ea41e510040ec4c3265a10b4add36f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h475a43e9bb57daf35028792daca29c6a77b25041a6f13a5146b225937f201890c7ddfb4f088d4ff740907d220b69532f733d1b1f541827913aeaa3d0a7502a2bddd4bd9233964d8372c3bc8228d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd655ecdf33bbbe01ee47ba9f0fc758a4f6e71ebb69a686d0b5e88ba284b5c4120a8e68ab23558625cc1dd338ae910b3d8d938a75880825d7362789ef8b1d1a2a03c2373dce52fbe2db51b2010994;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1249c5603e0598152df1d11b1ca98a91706114458d7ed0e80bcc359c87debcfc3ab61dd032cadfd1644ea2af7f5cfe7c1256164c61172997f6e37cd0c74f479fa57379e5be4151eda4abd7d981fd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1490fe517f84d6c0ab4e6889ab07dd75bb3ed6ef315d6706f1f6b8a0728149e509b74d6ff5b97339cab53342723d5bc81a3c4fe431828b94468b4689328929347d23270d374c62692a1f9412d59aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16684fc0c39a7bafd73782c85242a621bbd2b0c9b791463f97e023f340d5d153542c1dd91875428be0263b188a59bcda8bee8a6513023faab8751a9db826d9fae0a3eae76e29009484e41f1af6339;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b41c25982cb59f7342ac26fc7be26e8e2fc65046545cef7a3099afe3b485e33e3abb6d1d71aaeebbf9d507581c979fe4762c67891b6b28c6125d20533f9901338fcc3dece10922747cca2a22bc1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1321d68fbf4cf271ca82a9e950b7fd0bd21592e83ea63c41b0f453f890a150ce1b8f29c4239c5876a23652cda347f26104a08ef5895141e2d2b3b7e4bd67ad3f39cbb0250af817608e39d70b149da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45f21a765b5fb1257835795e3476ffba8830616640bdf6031868db895b4c867aea800dcd45c347b138cb19a68f5b24fe42ebf1f28478e3118afcb7e6bb3ee6fdebe04715664a2d20cb87ad7aa221;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5a2e75e3ea0ded6ecd9eaf4f97f11c289a07858f8dce6e6738dc989b305c10117ea87cdc575e8ba9a9690f0f67125bbec7906ce07c2283809e74f7d7d0d5fcd44e6aabea08158109aaf424c7d42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea91c0218f9d11947648975c107a2cf87d186c4cba15c258fa5aea5f18b8aa0e94f87c1716ea66a50b6e77e66ab203f2696f2a3aeed50048fbc3458d2e6d833161e16fdcea2e7da149f4eddfec60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10586b5f757847afc1cb30a813c7dd649df132959fb4e8c33559c060885bde27866d9a6301365786ff4fe77bb03512b093696fba94fbf492045186213a00eca67729e84bf43124329dbce4a76c6e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h522e58464519d0fb64696c7a5d1a46b3388f4309261941e252102670f4eb458f20ccc80ddfb7bcfc39c6b6485eccc3a4362f5faaa765d3c1212328969d90f65aa821601a3b3cfc0d87715234e260;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93f255108995a4a44ba62dbfaebe74479f7d7086e467d11e866d51cbe333d8e8009577fab99c5205c03245a0435231af8ad333f6a3f61cf1bfb95da1f4f69020d4008e5acca223b64c00370aa419;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a015b86464fde47ccb4f3eca81fb9fd50e5c1cf1fee285b7ca5351ffed03717f27274469e1813b613fa6b0999228febe1cbc45231150cb13fb69301798a5dc2eeb852b3dfa430c18aaf859c115fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16831e3bfb3db9c9b6facea9ffe0870739f100e511f0383e933d0ff1be30751cf8efd722ff6c7432b5e5578bf38fe6176ad83bfd9ca19b462c47ca482d577bb26b790266d836474f320a8b41b6a9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fb56c186613034765365118bece0f69c1305de91a8d957d8f2d87f8038e8f1905f20c5fdd8f17fe6e3b923c74b11527cb02268c60818f9a60a5c2df643f5456e40d04a1576eabec8e745488007e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1776281c644ccc6bb791fbecbaa2fa0c2a8a70c12b88f87639d2d89280ea0f5c8b1429a0625f23a811a8f33c5da5c3a4d7c236b892b1af4c87532b6cdd7ae56a28047e24c42887499d7957856af51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64490419eeba39931a3feff6c04e0aafa6e3280279a91f4d087b5bdee89e7ad640e837184f7e58a0e10c434828c504386b052e916751647dd22270b7bfa292141184fda9595ab0fc306a0d3ba0e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3314e6713dbc28e03169b17b082b4172363f1bb298aae96d1f2d83a1da4a5ea74e0fdec1195dba38cf2b0d0564be066032c835d37412fdaf8fc54fead2ba18f8426a0eed72fbec4532fd5040bae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d6ec7724dc0a4c4ce7ba733a88a14c48f81fea2d87bc451526e83ddfaff1a9f56c2ca4277969d088ceeb9261d7bd20e3e77b616e05b67c5ee77ec05848bdf77a65315f45fe96b73c72f38352dba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77d9da92706b441575fafd0688a17ea39287bb18be73100e5c3eee622b5aeaa26550c2118085ac7a0f03e3404923db02bd7f5166f70b6c8db0f85e763aaeb9424de82c3c87c65ecc47671ea17514;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0d9f1c9dd298ce53d39b1d8905c68c4e56ff4dcc0679aab2e3fc59e246b404ad747cc8992669b99268f1424d1a8edc6cd9d00edfedd7f06216df7445c8d562297d9517c8517dd4fef66cfc6f9a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb418d77066014b11d618cf881e7baaa3513b46a963cf16873796d66bc82eeb2e7cae8e7255aced5b4a058df0b44fe5c21f9dfebc3a3ebb06157a7eeb6f15201fe4f4a23deb488629e0b40772dc5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162dbff6aebacc8f5a2ce8454aadc74cb2be9045444f8a1d4256c2cc26efd995ec599439c770b95ff6603547f289ff12cd26fae25c9d3b5eeaf58002c924ef53614cf8b63348a6bf94a4da0e49d7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7b1a842fc769e06cde3affc3ab6239bf6bbcbcfaeba64e0db7c714864c7643d54c7e15ab29fb6dea4414e6c6822ba4cbf46ecfee154bdb2eb233ac08d92f57ee4fec52e06d725b55b23760923c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ecbed3d32dc2584789c8f71c31f9c45b20745731bcc4fc44ad593b87c04641c033c82140abefa98c447e7ccda6a2dc0a11b240ac4c3453ad67ad024011808fbaaffaf08e5b3e0321ae6a1bb2928b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h401a1a67b8d70f904befb71547059c9f8e765ba17b0982289cd517f6efceb7f76421a1d6f204adcf2b6e5d5cebcaedc270193238bb7ea9278d6a40287d3c8c294f62b198d29602f6c57212bebe9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h493e08848839a052a466af1eee48de815e023d32aa8445bafb0d8989cd0a9ade8725e48321db0c9ccf6eb234dd30537ab7655dbe3c1ec4b30f101e1e106b9ecbe98fbc91df24d42f090e841c0f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ef84c481f32a2cf3abb38a2d1f980477b82308f9af640126a5ed6b4cb2042d3b73457870e43b82defe79f66afbbc4c756522ebd8e5acb654cbb54199ac65ec0d2b44000d9b2f1d2d140617ff2e90;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d2ac5e9c7979b527228e49c4a861b177d292594b847ee8991ba0055aabbf9afa689798be32cf328beb40592e0cca56a5fe100eef885e7bf27cea6d70ed8fe2320772ba40a37c6efa1485f4be2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca8b863fc013dcf1e5177d8f4be3681f31ab1279ed0922938cae43c451258224dd1b93e4bd2898663f772ca7f81c1f2803aa70e3462a78e3cd861ccc74fdc592f9acd11e6dbf7bc91dc36e96679c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138c66a03bbec453023d4a5cdcf3d9b40af223e2180cb1fad84a4131a3c20bab2c6ca326b95e7e9443285c773b0f03ef0987495edd8d426c717966932450d8accefedb08e9a1192c6a4d2cea8892;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c163f19c553073464d33234d4afeb2cc9b3e35cfc281e39916a1858dfb4eed4210076599e6d2735af06f779b833b293651872581eb56842afafabfcd4d4722fefa626052910d0ac6c91fa80dc9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8f27379b0dc037dea1e2b1b1eedb5e4aa0e68993c1e191c2ff61f62ab6c056edc743dedb4d12b1491fa5b215bd85c030225c2e310d0b95f3a01f82e569ae2224d6bb03bc7bdd04034ea5eb53e63;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1787bf8b8d618c2103fa392ac902c2d6537c4cdb78fbcd1b64378d608535ccaebb1d45b86c474576b25602b72df4a0b6148d88b3c2a16b46e5eb89f0f7bdb9a403d784ce78ed2527fdce22bf311b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa68f006cc0a42eba5677da525539990fcf90f6076bbd8ae72a4246cbd6aa32cb136ad92dd2ec090d525af59ede7988e726bb011a42f96893ea76089e79b9a49f22fda505ce83a5ba8a7942314ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf11ee3468dd47274abe631efdc8801b71592440384e175fce7e36a217247e376f181c710bb7b13f7970d3181c5ed6cf7c321ac2d12584fb8efb3cfab3ce571371efb48f3fd39f5610b220ad0c1ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c79a0e44621dff48510129cf533d061057bc84b3ef56f004cfbad6a4ed9bf9c1d4b31ec376730398c29f32acea6eaa00b2037189a67207061a724ff59daf723682a7d6ee5ea0c4e49fbc522aa4c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb391453ab63855602276c50d9fa831e049a2614e1c540f9bc64be21ec2cea0de70705ba0757b1078b84bf4ce57d35d2ec659c055d17d8bb4df6322a24037294bc7096948132fd2694384adc328f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56a1a9723254ab08fb57987641e3f472a25f205722a06681c6f22c9b55bc5d649b62e690092c79f64ecbaec1a49e3803b74a60179bbaa7b35c8163d6c55350e95fb1ead428addfae7c8eb73aa834;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb63462c4f945faa6a6837817424bc3770ce582c3796871482597d45de7f70797a1a635d796ce63b89cc908cd22577906ed29bf42dbaa245ec1658275b34f4567ba5c1533ffc337398229e3e59b44;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b64e79709cbe4119ee2030174bd4c8791352184d09946321b96b1f8b76d385a0b512e71e334e06f930a8793a957c0b24e91f6db2b0189f77911083548048e8f1dcbd1f976ac695beae566849e5b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fa7226b4b744ad056a0a3ce75586803c80977cec1c8b1a933265eccd1288f9bd4bdec5fe92604557d43c50f881b5442d89187fda5d2d61e0139de556fda7591c4e500a390a14273b48747d36942;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ce35196b554e9698d45716e3e3067a8585d594ff4be7804c6128ecea1d0f974de50e420e9bffe07e21c1ef9104e81294d701e7a5eb4de20b2eee7ba42986f061cb701d87f62823152aece912407;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6e133e2f45e4c83dadde9e4df19e529003f506c8e785c8f7433f0c7e7a0060b0b3db4ff07c22c39e9af0e1d00f6c4426c42c4218ce4c18a42ffcb64086b37e8f0cb1b622f329a0fdf0922a7d8ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1023fa573ca133257e69524762b60f7dda6cadf63dd4067a527c829d308f2c7d9802d036f7627165fb055f8878fda0cce78b4d6bd66d4ee91d010461e103c5ab76df66e377bbb9dbd7a6ce971df41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d428f272057a4bf90e183d2b208428169b963721a3aa2c4419ac35c19cead9b24a46f6d708368603e267becaffe8d4e5e128f88c990c80a7f183de10fd6775f069c1a73d9e2a4ed2b85aed7baa5a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12fd5ed6e3bf081aa8028a4dbc6feb14f80a763c5ef3e9b9056af662474b5b7c4c52d679b3a5e86a42997f2c5dd4e06310c637d391a1330b8575e283d3df4e719db6b2aef9d69f07d9be5549e9dec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd32eb8742b78530c9c67436ccf5608dbc8afc17b474d22762273794c2330060f1ec4c086407f0405570f7f3b3aaec5f73018ee8970c6f32c2bdfdea19681c6ff8298745b541f67dc10f86732d57b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b72416385fd3fb6a5139081995e0ee3b8817d4f586a473eeb301cb478707cddc4345eecc594a963581600a68857066044975016a4b690bb54e459a0671d21d1a41451003c18f7d20265eac27a4e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cdbb0c030eb944344ac2eae14b340365217ac7d5c6cfb867f63ebd8eaa734db37d32c921662fc77e980c985c41c349652e10d949762e46274be9bb712e64261df223dce475228c86ca993abe73f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154d73d969f9441c45590b8a8556e32039567faa45cf8e11e616ee5a3bfe26175e865a25c2fed8310b2b12ba0daf5d88c3b4b7d1001364560b2f0de9239995391e630543e46e70842a07a531c0d01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d818185f90e7bba69bad91cfb83f3b0e8ce1a0ec63967bcac5c77d23d0f63ab992cc168e660e499da66fa172500d7010c43daeb0692d5d7c105f67fd04440b4f611b0a4c73e67ec78cb814e1f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b989043f2b7d8d38a900a93874b4e7c5c731df2d88db20249c1064d7abccc243333931ef0f1e281f20fcd88de7a1ea06a22e0e34176bf2e7a7d6aa53ab2630ad26b3c17f737972dbeea958340d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a64f86497a7e20f37f15cd1530c8b4e648678bf5bbcc653d5e86763650c31a43d25a502885385e661429e8e82cfc70072eaa33ada248b316422046fdb4b1faf28a31316df6cd90fccdcde19478f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65f79a213c98fed8a0d673b9e0fb3f0b5412dddf858b6bf7e9826a76bcee3f918fce53edbf4354f8cac9d08580f4acabe0f651302c23af31ef5247172c8b7078e83227c7a89a6c05624916e0c364;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7caa5863db4f9532c61695148ea445efd9e93141ff23e59a6957c8042d44f49ef9940dfdaf5d1f611bc60809c6e20b3edd950c1123bed11bc830edab51f5829b14d8be6c1dc1e1be028407c1887;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1707a62ab2798a7d0cb3090d060ec03c9248fdd3354aeb0cef89da186687e20064a29a12ba3ceaa25c199c188ca041ac43e3cc3a8f44d55e6624f15e98d8b035f9c785598998b446dcde01cc45233;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9be8e2ccfaf1baead6a129c996caaad502a9d68385dbf34a5e035e7bec7850d5029d6d9416b223e300740b086468c9db8246d1d4a332cc7c528efad545390abc3266562ec2f618fd2ee60a9617d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5cd7c2e17bad1c54340ead3fed3e270b47bace2f23d586a3808af0a8daa9f1a0cc71421ad2df3e7b8ac0e0a4bfd177c8e2718d6278a8523845df4b3c7ecfaf4e1199b3ada380d0290dbf89486c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d433fab964f14aae29cfe8bbd2e9649fc8dc4a55f5eba07f87bcce36fb30913c2dc85dc2b5661415a76b5b157e90cd7c37beeeeba27770ef776b460af54dffe31c166a796703113398b322d1627;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3eefc39fd953bf770da002101c239c814f109a4c4e93b9e160daa54f1339523dd427a896c0181294f80200345ed24a7df16c23815060a328a9ffe697dc11d078981fa4955c10b03f6cca47c4d5a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf11d6e2e96ef1443a89c69fc07062e14799b9ee9332c199fc34dbc1660975fc4e865afd66a881d7807cd702267a4b9420a1ea1746317f63545ff46cd3d0ef29df40d668735193330b26a344f5588;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50f5a6121aa1dee6fd17c55facd3b4c017f2941d1105d6c1289d9c457dc736ad6510be5c41bce90a53b567b0ab2f330276312a590e5aee090dde09be8789bf2799af4d284144285f36280a0297b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1122c1ce0349a459b2ce5f7a6ccf7f1f9478fdfd1a7ea619f8480131decb214ce840f16d8993ba9ddabf5f955fcf821893fdcaa98da984952e1ba7961f3f99ef207d1384317707f894a4af4c30428;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115078aa6dffb6d4b1007e75af76631b0c7d650a3ab2b3b92599cad06b7e600d7d7ed1f912c583ffbc9767f678f0d7e76efdc0990fa2de43c90fc182c129be6da3c06afea33c3895c431c614e9d8e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ebffecfa62678f3c6c0fcdef5c9276b98b92e19e5fb9916145dfa49abc837e7da7df74b77a2e702fd593af6f5bf1b36b41a60a6acee2438402f7780a641408ce756fe6fe16c90618e20aa72b01f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e7a0e0b52f5796fe247f76b652ac64d6e9b5c8697496d0c22966f15c277c62ea8caf02d206d811c2e42a18e82e0cefd8d99623e63eedf74ecfee97918456a4b4d7ccf5f7ca062b041d9660b1222;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcbc574ba326870f8060029bfff8ce507d96f30ce1dbe6a82a5d6432e97ddf4ef8bc97bfea14a690dd6f7a4c2f2d97f0ca20e237c3c0797d5183ef4b6f1bbc889522cbd769c467ef9850e436dad2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16333d268d9a0d43402a2cf16854a089dc40c45acf5aa0fbea208eee38eaf7ab18905db402adda6caf36a030799aa2ec7c747d585ab5945f41d4b528631b46454b394166626a217e409b94e69dd94;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b0c3d6aae867c4c44f4653abece6a08d9aca327c3244daaeb8b53f82ae4610d5f741616af8f12d2bf48c39dc38f5334174d59490ff2721640dc1e52ed6207bcecbb00620247eec320eb1e55e208;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e1533ec84ed20e0e9c2d08c0718d00aad33826a016f85fac7447e84ff236fdfed4b93795faa1c1c482fb3f67677f45777cc66453bda4e36936fb06e744ef38c0087ae82a799dbc596d851aee749;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha416a11e50bd81ad76236dac9c25c6671a1d9da5bcaa47a801ef318b21827aa014f306c5ebc25fe2a29cebd8339cef80795b81bf88cf5ca681092d15156acab3375a181192e164e4e0b4f931c445;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he40b9bf9f60a20cca8a53f0c230aa087848e1f1aacca9f93b21bb45ae3660c26def8fa315449e1a90a94cf0a102ea3ffbcfffb1d257a00f27dc88a004c0f9a8193e652ac09778571ede92ccca830;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c8c7b23c5802ba70461a7c611074e13153b74336867aaa507b0ed61cd0efdbc8d647bddd5c645b511b22d240e41e955d554557ef4081197cde70d3472b83470362100beb2392dd0fd774273b8a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf55b55f2d03b8630b711e84436a0950d2145b76782fa8e5da0ef931a823f860d6ad39a4655915cb57d946d37ef6b5b8d982c60e76ac69ca4025b98b2830d67b929bb112bb446037bc5f5ee510b81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b55a0f590057a3e418854cb45aa0d1803b2603569228cc28210db7aef98823f5addd93b0845d3f8871cbe91d36d508bb7b5576612ca2344e5782b98139b81bfad589fbb352d90e4fd3207703ef07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9420368dfe363ee82b8cc39a917a3ef88942596c756658c10179b9a6fcb69414b80d35511b38577e83312a138026fb6c8b6e995b942a9ebe663ad22066a229ff23ed7dcf28813d048b263dc24c30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc53f252e5d0e09c9957ad4d9a751c8be87e7a8c266b5885399aee64235260ba220c59aefcd6454c2280314a06584a9d07d78fc722d9c4e5b272409c34c245919abb1ff33386286c6b3edff1f58b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h41c0861eba6a104d4b676d110ef4369bd299e3d66f312ba970ff31b82e564794a656df7973ca38680e6316fb5d04b5f794cc0752baa5aab289e36beaf03f0dfcf2970f4e25c4e125acc7dc1585e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f449e0eda4c52afbf81ce4842551b59bb0b18c9dd7a9b9305da8c445e0e437f297b481b5cbe86ae65ca1bce9b2e32b6e5c9d5097aa10bebc05c016620c2e07517de6d957dc5c64a7ebec5edc944;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95173aa1d93ece160695ef80ac09705fe553e40dcc62db0fee6ce2cfa479296a5444589d9de718584dae7c33851aeaa9d58ba7635c0fa76d31b0811b806a9648f696c8f7186f0d18af17dbfa410a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40d2cbcf981b1a5c6d5108266a4a369e30fbddd0616cab88171bab1aaff58896ba5bf4972e66191ac3d5121bc1da69f394f98fcb1e069a802958c9dc2b626121f832bfa671d0e0af18a5dcb4f9a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15885ba5d1877bf2b8627ece997dfe076aa9f57fb9af6df7ff4aa4a77e387d2edc01f75043c260db51e9496faefbe50aa9ff671193b8467e347706978c03ba0703955e90f024dd56feb292fe583c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5d626e79be55fc43650d0c5140ee87f11d781a2fda6c84199a8fa466c2f3e427cc5c54fc00f5ca95b27a1d8f6fa874286778afcd774156d04752af6f797d169d847ca41bb7e125f890c912e3482;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117a06d60c4dc819904187dd076845deef1353c39413e113f98b4ee9afd240b03c63187dbe7ab725f1ac648f994fd1d21cd83a33ad1120c81585a59155b624a1b71987a77e4fe312ac9451032bb81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98ffaeec944444b8fda8562b842208395663d52070f3d55566d5ca9057f9dc8f5b6962492f4f791ecc985ba131c1cc3692e825b02232b209fbdd3d935a354022770f76aba5873fc67404bb29756b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccf6b85cc42f94ca6675bbab3a20d97643165cfa1f76703dc1c2d097e68845097f52114b1ba9fa7c10c4e3d2ed1d97a40f5a2e1cc571b828f9bf49ac6f8de969b49ec62f72ecb6e09ddad5c79099;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6a90b23305d599ed8f72b0ef96a18f994a30e01cf7a334577cd58ce3fcdd2facca4b6efdd9181019040cfb5acdffe17fd37c124ae7a5a93b8771dda462cd5aefd0f8dbd5b9766a6a8738e55f0a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h518c10318f5c20bd80ee8f60d3f46d9e4f5be12e97691545e6bdf5e32a22a2c03fdd2d2ef2f020b8a864057fd2b65f8a425658e4ce92745e13a086e1dd4f45f141b75d90b0b710cbd901548f05bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df12eba1a4cfedb5ec3f14729f5c85aeada88454a7bc81f7dd56d99de95185d894360af549e4b2257e77f2cbf36d9a4be11aeac1918afb099aa8923eebeb10ce5c82c9297a05ef039c7f4ce3a0a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132cf37beb220071bc194a642c22fcdec057ca773a8cdaa9c535495e26770960ba8fd678481fdfff831501da220935e8b5ceae9414bd172f20ea03d47170c03b53add1ed576cfd7a8a74de32d8fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130280258db3d43716c3d1e01d90f3f60759d35926ba106234d7809658222c9150ad2843362aed1e376fb9b98567078a7eaa17cb8f60f04fa76b109ced26a2f5eaa584c2ed7b2603d0be6d2e5d96f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f47b8a400298de63b986cd2d63a6b5f9b1850010917e3f7023a0e99a6b971ed55ad6a2f6b66beb9c618bf682c16067a22d6d061c9f70ea3d68ef19bf646f2f9c64b08f6784a6ca1afea0b9b15f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b94f9584413b8ad84e3cfda1bbcd865b437e291ed0fd01ad87659b384c3bcd63bfb65d3418843359c842c914fd06c33ac1e83d0939969840e04e14db2e91218b6be2af45d2f3e5b73090ba23cec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e50faeafa1cbb598dfcd62a35695769c3a7bb41dc0f5e81e2fe4bd578086c65df2453f1ffe93ec8b5bcbc4b21dc1100184807355cb8a74152a2f75fca638627fdf14fb52742c08120f01517c95f9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16086496b8e9949785641c0bc4c7ad48568ce2a117fab3e475c665016d58ba489ce7b1486ad1120f98595c5f7249d644fc84b36a18a100c281fcd48fec59dd4fd81af58a721f678a791f4283c0fdc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1151402c51ad369fef4dc88140ad8216cc4ccfd25ab207cc248bf367a0b70e5a926efd0884412bc7877ede5752d6c7cafae36b18580aca92da7ce98224269f7fdd6d10211c9e6e58e8bf7367f0a71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6c18ef2093746d551fed6008bc890c5e1d09eb539209d5363f000803a77b907919d88ecabf6ef553fde628fd12d59373000fe3bfc362f745be398c85328c549d441a0823a568156d816ec08606ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e395c073b22fbdaaa5284311c767ff8a576ff4d5681023a996365bc101792ff0849b758698c91ea6258f5110106e9f5c52079f586964357cf856efdde9bdea03f6670c15051dbeae6f1c5dfb5c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd41b69aff4e072a1cf871f0dbb4f2b93da1ce5d2efc8dc7eee4e636281c4fbba2294d75343ba075d9d0f94d1df7169260250cfeb879d744e79cb81602a6f5ac0bd59a38d9e811dbd094fd393572b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf62f96280f996ae700430b51b8f845da9bc91de08ed58a1a77481fd49263ef3dd5d8ff1c7b68eba1e2d04d615ee8da3c1fd97c4042ceab907b63459bda1ec5da7809de47478aafc19cc13dc37ad3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12301abda7f16607f7c0b57ea27e6c9afc64c7daac836d5c64a813fd274d5aacca92f9ade0149df50a44dd987a26f70ca5caf0544926a893526e9c1c1261a8ec07f9e93500db41445826d40af30a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a8ce3110d75f816a0a2e15786f9001e80738e7ea44f92ed998c0df7042dd1d6a7011ef017e296250a31dff2f1179c7102c697fd8c05ecd013f4d04dc98f7a89caf82d4508c3185d961da39ff5b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4a413bcafa34caf4ba72145dedb017052d3fd1abce78ad7c03e6cd66528deb59dbfd520a11aa77a994ddd80298b0d8d57c679b16b40c47b4f4c53292d508e75deb96e7d6dc9a619dacb3467998b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1220c9d1ca82d6d3f82a22630af4adfd872bd6cd2e89508d16baed1d3e817d4351dc1f9a3aa057f25993543b8904f273c4224c45532aabc58137c24049b21e5e6b3b5bc9d46751179343113d0628c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab1d8fdbb274e7850fabcf06bd691a99155297081fb2727e3c8e6c91ef4afc536cb9be964ac8331e78db324fa09e9843b3f52043f77a2c4857e55d3b72e37a4b352d8433bcae8473bad418b3ec0e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eae28e330cb12ede59d8c23474b8107f2bb20e87121bc58a228dab84725954d8a7ccaf831814b8f022c3bd7ef784b0ee7e1ecc6d1e31019802ce6723c00c89de492f802bfc548020e67ccecdc2e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4358545a7ee8b22a0095ad454e13c574c73828485e73a32cb35cff11a5018dfd7e0ec2d4d12ba279d0386c2fe46c9cfebaea18fce7db9fe381db3acedb01441354b70ea4bcef4b820e7793b679e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a7edcf782cf35d86005a2191039a68d589884205b08ae4350d0e81182bcdc389c42429d8a67783010ea7dd9579034b862d5460ab915217f985ac3ae05504cb6d3bc1f5500daf10c01792fa3b09ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf360d512bbee4ae8a0f11309940be6ea3fc60ce31d050524ec848478ffba30bfbb802074434e19942501df1941f76ef0fa7f5e0211ef7c35199202685393ae45550513a7f8ba3e4c1dd663056504;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a896be6dabac67a7dba5effa0188402f64eda1c006d8709c3c1e5be0be8ec904d49debe6bc8bdaeb1e6f03b1a435a61351727d347543c89f6a65d8cee0628b09dd394a0c4e289467caa9da17f3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a3d631b90aac3f6a2b1b93bbfaf6fd5d1105072121c41cbe80f344dfd541c62cc72a871beddbaa6226a43f1295b27d89e351119a4a493833ede209cf483c8fbbc3860a2af6d5aa50a95fb2afbb2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f4b38c678d0d91a8928cbb7a67fd36724bae0ce70d43cdcee885768334bd6dacec5a4815edfd50b1c524c70d2a2b9d162433cfbb3ce43a2992ca09b5e45a2f792a6fad120ea94657819af2ece8f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bdb4c0798196dc49d8caa31e4ff2b2e17576aa565dadeafc4d75816ba17003a3a548516f900e60f74c6b9f3f16ce8d6632ff1c3ac00ab474fb51fdbc9d0e3b82b729784bb7ebf3a0986d707663a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h499f789cdcef7664290499ae3489c7fbd1e8eada7d77a0f4d7c39cbb895e717cf0c9873a2b8e5fb2d86db51825ff0eb01942d21977ee33f8f8c6bf6b0ab52d6f8a9aae882633b6297064460e4929;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148cb8ba1e08f2a37ef80019cb5464838fda65239766541bde746f02778ef895fdd0d43e7637336d83161c71ce1fb8b51b36bd08dad8444b5bf8d2659421a433246831b60ea4d5d0ca91abcd6e06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113008130983918a5f4f39ff01f65661cba68673e71c03b008dcdabfde48ec6b089d4bc1c17bfa6f89c2f119a7be638a63eeb4e137cb3ad62316abe0ef69375ec89d5e430beea0e20ac495e534814;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cc8f084a754a7fda05cf83a873c6312d238811e5e002b73414938aa6f4086a58fad8d9bd89dca5ac2b52a7c57166b2d98977b3ba22afc7b47cf67aabf6b8db394620425854e5fcf36dd8be390d1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1929b6adf538ac3e2055df5fa6227d6ae49a577943b6d619155fe3166e3af007c8c89b706ec2b43b3f6f19ed44beeb89018e47e3725d5819e05a1a6b72e0293cc603a57e835c01f8e13c575afaa76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65524107bc169edcfa8307ccf745344e48a47279a180a3cb968b23e7cbe32dadd01547692e32f541b6c8c8b6c69f5eb0274e9677f585b21fce4f4ce35851739b604892842b15f9622eba7dbcd3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1773f8402974823998f5dc006c2ecc2da17e350e0b03a04d65540b8b3637134b8a3fe4c4f9a6b0644a22156f45c2989ba644f8b0966c6902c32346472b125a1d76b3584ef1decace765835eb58065;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf49d7f59f39c4cf814a4cd157dddc24289862d8d2e3309826e0112a4de8829f0d244b8e386b80a3a03fed8dbfba635c0e3ec0265a933f1d3991cffc2ca1a9e68fef2e91134935fcd1e460e7aab6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19796f934fb22515e69c195bf3c1390856dbb89ce33a6d292af4174708f33384f652c7374e1fe056026cc78ec9fc5a8fa2837748b28c15378aa9e13992cdc3a6cd0513ae3647bb384cc8e87998572;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fc3a3feb1d3a5e8f8c46669c5b1b90bdb94b4a4c08a874dacdc91805df5a378909adac28d03ff601fa416aa824a60f50dad2afeda89cea913247196d5cf8493908025b1fbb78e6eff455726bcf8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h338fbf5be85f55a04d7c0ec4e6e2fa459a11fc3af9f6a139468eb5e2b2a00c75b74b8b4a6f553a631c81a8c5b3fcdaaac59e62f0ec2cb4e67005fa7cd189b4d88ec4eb5e190842cca9d7d312e20a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98076069a13abd5acd2bbab96e3593caa69207b80be317f2ada11c8e34d972304a57af8e37fdec8a19618ab2f8a2685a6e74a7ec2f5d2de6ca529d46ca8419849106fa6fc9ee33747d2a1bbf90cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6efc9a5a81b2a1cf0e86a6a142a74ef266c856073a3685f637cf9d1165363840e57a1569eb60af95ef550c80aa4bcaf74a076f25ebd3865333d49fc69c9672b0ea90328f8494797f406ae4389d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132c104d0dfc7876804e9c72ad2d341407fb303b1934a75c80115d88638d017634a67d3b7d8582b3833a2d7e82769228dfeaeb2dc4059dcc57509a43792c335c3a42915ff10ebe823f53a91ba90a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h132a8fb56b1b67c52421d22ef9f4371cdb6507cb56cd31c5cddacd33e1dfedc71bd2afbe83b41b034b7efa3bc55ee9d914b3a9657858e57d3c1603bd9b3881940ede3db26f65d44173ad4c41517b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e8a670bead780a63bb5998ff6433b618a5d4864610ddfcd6cda6b0a372b4e9d7454b6108840f5edfb83de971723b8f50150f8beb3cee47fa1b17fbce66e3aca84bcd18c11af37dd01b4755cc287;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4decf80da73c927ac76bcbd60dbdedb201a3be705c31bbf75d048729c61fb909cb461682e2d05d5be5ba361f5e6c6ee0d1db51d48437e6f0b00794602960262caf54fc32cbc35b6076ecf83f925;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19599de1248a5a53b13dea375c82b47651b0f78347f2ee61b49361b2d1345776bb0dd896774c37519d1276eb32447772e82c1226286c57ecb4c77e7d7d0290b47e4118a91fa2e9f9479d975c5226a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f320a7de81b6778797490246c758b87f5941c6c61a5565d59ff074bff1e0167aefca210f18fa16bed61320ebcb6f006c914919f012c081e448ced908f4e78986001830f9eaf7fa3450435548a1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c14561159ae74bfab473b0c55847fb993fd50fe28948761cb2a2c49fb2e7c8c246c6566ff2aa80744057672949160facb927e1f089e9841238902d6936f5545dae58c049aa1029fbf38becde64a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h436d0f73ab5eb10d3226db58c1447e79907108c6d2d50ed4ce32e16e7a69ae1cc7f113d1c443d4713e8c404f737e213bd2a197ade0681928631d22ad019f073bf393d63b5e978d13bfec3ed46bc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bba0c836ba9f2fd4572144f1203604f88e1b4f9834da09f999b48081ca904968d078d8a91c7926d413a694f5ce5d8b010025f1042f03b5724c8487e38b1ada82b6d6cff81eb5e8706bfebfb2d2d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe3a1c2fa285a3ba4bbe2330422b9f0de29f25c8d996446a3347607a2d05e81c7ff1d0543ddc23f1a091de5c06a322749b4b7c6392a56d646f6da2b1338ca69d743b5367112b54c7c30dabd023b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2a5c5381d75c20478d5be2ce5e0ef06387be84cedea3cea09a171a50ff4f08e086884def22e9a968f8db585fee943c93957f9e698ef5a9aff2d818b0ab41e4a7ed6a2aa921c85882ce231ba02e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187ceb81a94d024bd88c6ead5c52b1a62b90d4545277d3cb7ce8717297012175c067ccb70e50709987fca3464961b4b8ad383f013555d2091a63ac46ceaacc2956ed6ebe350edf71933a403cc60c6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169f9a83709ff67a4c955218534ddcf45d2038165dbd46873f240db6f4d9621d86a3e53bf8d7c8363c374a65455b1b5070547f4ecbf028c2b8dd94418a3e2de80ece292592fdf0ad14790935a4a43;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha14e8cf12f83c769c4ce982d26b8f8781ca96ba0bdaf943d989148e727ee356e3caad2f476fefd8244babc4b4eff265440b27c28505d217c6f0790a406ad2362877cc7f730dd740f3550adb3c50a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f070753d6b5dc004690bb79d2277dd5421f21aebb7e99181afbe8f23494844c697150466a2b114b856596adeb56c9dee758b14bda06bb63982357420d9c7923d9fa91c35d048ac5f691367550c5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6177526c0c20c960b9fdcd7adc05caa699074fb4d885be75e3b9bfdd195a7bf822a347a3e33df70cfee6a9fa0128711e6a036d52371c8687ab77f16a92c6fd3944f1c458f1d2167f9cf8758e57f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2ee93ad64f39f23eecc2fa4c871d9ddb65ac5b22e1f577170c057c035b3ea494136b9a4ba997f6342e1f1e6119eb86c1cbbb7c396ea2067b9308f4bfbd44b6d62ea819ad9b4fc79eb9ca3edf442;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb33ec5795de71b0fa02119422b869921926f5c0e668e4b7ec5c37f966371c31679b6a16d8b3a51a66b6053151462c25762b1893f1c7cc633175ec69e3f862a99c3659c3f06ea4e71e1e966bfce5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c769d44f99b5d9e4d9f74c1421da2feeefb62a349f1d4d3c2e62b7d5f6e9debbc96fa03e4c46a0d0f30531d19b9ef1545c96b391d21adade9eb3b5fb5fb42d51f8ecfa3ee92679910d94adf49cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9aa978137b355150fe3237fa05222bae69775b5e153c38f2c2f3589e30aefcdd6e864bd27cbd3fc4779585ad9f0c98cf520e6ca0b78fab04ca89b12759956f4cbb61122a4f06ea03e996218ed4a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h557700b6d5e4e9b3e645358b3067699b0adaa4174bf43f88f98370c939d7a1095f680fd8e333a6af8b4d4a13805a4db7047a1a51b23eb4c58085a84f647cb9ac3a2b0a8555308a6d857a19370820;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7e068eb6294143220be0b3e4344e5b9d74fe0870f8f7f8eb0370152b570f38da3064e80113dd07f00221ab99df1e360a9f0744d72325c55f1646ff8ea89864ed6071af2b92445491b3270ca1780;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd66b8c19c4d309048d44b2df07653e187c91ccf7c74b14e0f12362f808a0bcade8042b5330f6ab010e9c59229c2886b6786f6284a49b600a35125fac4bbb462c6ec3e715ecd56f481e5492809fbf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bfaa411d2017d057c4c4bc0e466c33d503f90c68dec6b82251bf0b11bf7a06199cba848cc6705fb57ba2ebaeb3d3d39ab51f1c7e5cb96f311a43a1f02cacaea20643e05c5d9ff1b25503edf11f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d3d2fb43aafe9f1fe05fee65d8717675f1b2a150363670f02cf2a5f9729a74ec08cfb1a0dbf053dfc85c5314e574b1ba512e036b3cc5c1cf75a2f390055499951454464d447eb0c4cd2a1595d31;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19128b286af4f1d2cedc94899db88b2250305ef1e99124aa0566291d8487684e4d6de0630be63e0b94e3f201b588105072af3e3746c865d0b37f14fdf7a58d86b3d160f32590c2ede26b8f377a37c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1576a9488c494e9f5a37033ffb2178853504ed8466c96f270353ffad850b55042f7c3a134f437fc2910b2242e22c8fc4cd71200505b55f2ee288d960df67ef2f755bdb0259c6548aa4ab306ab8ebf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c21f1380619dec755b448c6062df3d0c31fa2c9e6ebf4e4e42a871176bba9f82c98d41fa25e6491a3daf06b119edba607fb70133328b8185679be04ed715788ad076c805b572a56e74a7b2414597;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113d28809f28c1e349c8a56bf862a8f91e86c51fe2cf67c8df4e5709e70be2773fd99447e102a7feedfcef0520481213f9d00fcb9ef7805681743a1342925cf3fdfe29f612db4243e4c158e8ec9da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff1cd7320d4399f09bea17dfb00841d587ba183a52f20decd39ef556710e9afe1c7075875e26fd40abe3c6b650717aae437f05c1471cd24caf4e0f4bdb21ac51739949fad715bfb73089c86e7609;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9646d36ad006e46a24eafc81e6a9176ce05546b8085556afee428d43ccf14bccf6b12054abf8745d9c1cdd50743bc2f8996e597556005f90dd61ea8eab7f683f8582f336a4a787daf2041d9817;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78a0ff4b69e565beecd8e13eb73d25b88853a2ec2862d4774bddc27a9f82befbe23649b87de01da1ea9b4f74ab581b3ee8760350998626d7c9cce847d82e8893a9678d865c531fb3a80bc5ac4c36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11eedf8f50d7d6aa4f51f6f988b7fc1a15faf7e888ef3c83d3f426225fc370f7afb8c296e715126457b94d8998e635484a8a5c2f6cf5b421ef09d8110bdfbf41aeb6ceeaed0b631041a15824da624;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1223c9114968622e890e21c14891f7bed9e913d2773ae3609c208dcf7d04bf3dadbc194fadeb7c0c4d5f6e14deed41879fd516e677471ffeff7512b5ea98fb08fe05fee79901edaaef8eb7a245c7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h872cacaed36834314576520d9e20f766f41e9302c6ae7148eae46d6d818b737be1b5be155dad20e82cbd13e9c3d08162a174c3613514ea3c12456779f254c3f2e61415060d46b3adc853fa9ceec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h484038a0f55b6721703b8d9889f21e694eaf29201da17e682c8f92712eb74b1f369486e95fbcfd0be56ec9d793f5493ed0eb131761079da80d4504e6cdd0e2bcf12d3f44b5022de83baccf911e8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h273209941b97f8273593864660d7a36d5f798f5ad4245700d83123f78fa2fff2e61e286e1b14e5f4b6680f044006c6434503d375b1cb70392ce833847bb6133f532ce02cedeaa7985a3b6da14b98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd363659181d4f27bd5459fca50f4767e8256b957814751ab45d39a11eac5760cb8a202d420e9eabe50b3702a4b614eb35cfd5c7b85681f585f74ed46a29fb7b1d2835f1e013ccc843a7451ebde0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba3340a45261a02c5423d82c6122bf74a0a45b8d754a2dcafc0c4cb893c4cd227d51beeb0c1cd085796ddb0eca1cbdfc8d755f15d43401b99240ae4352fe1c221715514ebddba2304373a1645a28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c09f37755c2ce316a9c548b2794f00d959e1c74752ecc4c794215b3226b63ddf7ed4f08fb910cd595e749d9ba4eae9c7a26b4832a899cf3167f702500e1adcf55bdbe805e260d907a95774d7968;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h602203382344e9c01c96cb1ed97a6a84eff401cb757a473abdabda08403999aa46839142b3a1b7c60a0c0be1fc493b8f401fdf9750c202df75a4bc05c4b24b2a48fbdf7efcecc73d46b9d9da954f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17009a100bd340cfd4ccb6ee278cca97d0e5a33f941e22f2ac8b82270c0b4baf1ea9ae451676662916c9bcfc1bb652b85a2197ca87f5eab40aa15dea7d04e62847562fc6cfd773e011b46202a446;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17753c656d1ca997d41f7aeffe660ece0fa1c8dc788f274d191827afd5fa8de00e2b8f2d79f6c82ae5c772d43a34f30a9f394ed3fb17d60aa976ce16c66ae891eb782a27e8ec614c08c533c3f8d2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1263540c13b11e4b3183aea486560d938678fb1909aee710b8dcc093b79c50a7db1169389870c897ed5d4c9eaf827e304a07869f54ac8b271b17064637bb5e9c198c027563ae401074ddcb592b3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h745fadda07551dc515df2daa3fbba88ca58eda1326cb141802e18dddfcfbb4ea3c8d9e08848cdbada7c46b989472dabc13bea55710524f22a4b229fa62a7a37151d53210d7b75b53a1b89b7a403f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1622bcc1b94b460790d3e6046970cc3beeec1e243bd375205a39d7f27a0efeefbfc1b4448147f888e934c0d24ea9f2e207b778097c266f6749db37439ab27eac1aeea5a3506abb2aed3c051dee686;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35b7e60fab5741f96f22bcba96cc08f29d76a9f9f398e352970fa8d06ea898bd0db09db36693f5f394f569d4d9da348d35f8f16ffc2e58cc3e50de112801487de3d99584a73abe67ad045ad28c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e49ff937cc8d16acb8a4551ba6c770eeeee9a2464a12e57acb8e8cf99ef2683f379f1d81940d8a89d7331c1199278715263d81b13c90a253b76640f3c1e54620d654b0823ed3e1166026a539ab2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h81f55fd1205b0af541e64e9196f51104aa6a2d580d508c2000449e3e61216fff70d7620ab8fcbeb354b65bd7ae50b79fe8d2b06f6af844d4573a5ff82b2cbb2ea8fa80ead8bb8cc377680f006b09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a7205f6e2b3ba6550a070ac5c49259b6e80b2b263423c62cfd3d2f6055c11865f904088427e4fc82d5f07641497cfec7d6e2bcc579907bf2ef52635258326577adcb7886da3abe24e62b81736c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f4910e60cb2da05d17c7ca1cfbdb38dc1546723e2f8bb5b8d3a50e0962d877ae50adf7adbd6602c68db384c2d9dee047f4925e5e9dfaeaaec912d03bc09eaee7c958c3da88b57ae8ca58f108e83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h477fcf792807ee8b3377659c028632522b60cee89179db0acbda60e5f7e7db1e2f4eca46dc7f5aba1b2ef4e2c218fff8fe4846b90ada1c59150b773237e6e66b0616ffc6dddc6d9581c84d21e6f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195791f2fe9e1a06b4fb17e7e55cd37602d7ebd84a74c453973ca732dd712c092911c8f0665c68ba459e46d6177a6184c418e77dc5044cd20f91f6498ec6a3bc48502c8ec4d483b1a3ee09a47b0b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e1b116516e803ea4ad6594ae37f20da61fcf4490194f0fcf4d3e4a209219fa84c27d2d1b3770d56a8936fc283fafafdafae1b1f5a1b8649d68bbe19bab18873acbc772b1df68faefe3fe28cdbc13;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56d46a025fa79ff7fd74abfbbe2ae6f36123fbdce9d6d848f5db77e334960ab4d6222cffb6e8f3812fd8ecce05ca323402473c9d1db8f0a6f6a67c667c5f288da5fa0dc4d4b9ee84d538870dcf51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1252895d880074fe742a67d5028121ccef7137992623eb85c8d2a0e8a10827cf78368b4683a67eddef12878d047e69d32273b19e6141fd0678fbcd19cc2cd91d4caf0752cf88d551a2264f9b3fe7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1096a3bcc2b9691da550bc915bfcf0108a7c3bfb0d6234429763bbbf9c7c69c5bac3aa93f1bb78e9219a15ceba3d28409d2b4f720b75a1004bfdeb6bfb7be2d839ab865140e975de8991e1ddd73e2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb441bf8df3a93bd2c36b8bb0f5d078f67b5d2ca6546df1f89f7cb7e7a00e64f08b270fd92efda3080703e0911732a62e0d678912f69f55559a870bf17298928df650b9a808486333e5dcc244578c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fa00a77e4486ae3b67f77fd37c445c52033d4964eb1598113d77a87c8fe1a312abeeeeee57ced7dcf5d20ee4b36731a08563eb45d7ef3a0cf7c2931626a2e7281444fe826d0791261cfe73d1880;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2e8e22b5813b038dd79e3d191fe132d12188ef4187b2c9a6e5fe48d0f712092fb11b326f86dfac11c5ae772d2e08882df46f026e657167a16f9ff1bc4ed5483a77d8bb499ff489d3c07eb219bea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5aa91fe87ca8779fe26545c6a991136a7eea4ca8bce80604c0dbc1f72714a7c838d7df5ab7da37a1c1200a8b36880db97392eef41720c12849e5021c0790d869c05b94d19fd814b23167564f1824;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde48d16e3b0b34b0dc5581e4697225b46c1bb233b2141cf805a6019ebef698bd2723925828cedb23c90a6af1f3184746df6f3d49610df83f54429c3bd23db734c16dfe96042e4775e326de7ec61a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1489476d8fefbf7c54f70092f943e1f8f060a2ff0d9319fb89c70fa1dc9128f78c30199033005d25ce8fe16bb71ea6e64d5acdd86e82d6942e9930b7165c01a29006a7cd283db0a743e2412db67a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hce27b044039a59175f626cf14fed953f3fc7604967be46d3782408464d8a3149fb9385b1ea565a18e7e88ede984bf200da8c2c24d0dedfb733e349414ccfb4d0152916ecd7f2e9833f8de5e016cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1af1f1b472efe9bdb5365e3de6b366f88ae6baae98242faf6eda0e4bdc3bca0a85eb3c26b526ef763807e8e52c161c8e8285a86537190af09b7dcebea06f00a0193c4cf9495c061224977eb114d3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d851643877fe65204e8e94b0a942ffe2d44c57dc989f581c7725583843e5a774fbd84e9cbf752f81dff472912a288052d203da135a718d9f5adb73bf31a976aa687f6a2ecf0d93b21ff9935db630;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8c26bf13461a99ac22cb6b96948dc550297ecba0e10d24f331e9ab21c0f6a5f0aa13785ae0dda0dbc21e5c2a569c1bf7b0558e8dcab3c11b9b31c57c8f8dc9ac240382e95b2770beb4b3ad323f7b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17495d885aa35bb6aa74ba5d69497c959622085a2f207a5eb2b6cf9643ede7d8cbd316129da5b9c8f8196e520c94793c0084757a543214727ababacc43b59db715948f01279314a1a99ddf94ab5d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h655ddeb0119aeed23a9b06c0d74639e70e7f43ac8860e9aca585048c2ff23ee53c4b3577f3872944b4367406210ff12baee166e51b73c7788904656d1d8cc052ad7b09caf85636b452024e1ff399;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5555b291d6562efcd73b24e9e971ad30a92d0c93ae625c8dc83466e7ef82d7481012928a91dd0f43311ccef53c4a513e020936c3f9938e72e062ea7b600c80d2c41f1999eec27770e0c1afcdce49;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189a85f579f8915ad8d0e331ffc45debd530ad37db57ec6a4da653661bb28e4296bba18cab9faa01ff54227a1bd62c86dbbeb1f013d5d535ff0a39c0100f3640d3648c2a112719a7127aa4bb7b471;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ab20bdd02c6cdb0414adb7d063ec684c6cd4436e9b73ac9037b12b5042377b1a57c37b792faa149d425c8f9712b0eee12f5042294aac5462b77c3645462a3dac9a0c859a68102c67f408b053463;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63bfbe6982de209df1a42d4580ece211e8f9749d07c32dfddf8fb75b3be9bbae93664d16ce6ec38a8002cdeee6a596dc19d0549b301984151023a65e9daaa04fc8d92ddc30708ea61fad97a7bfb9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb286824bcbde626e14ec6a76589cefb8f82011d78903334bb3eda633caedcee7c90c3ccfaee1585768c3361c4126f2968254702698db8e36371d1961d181c22eaecc2128aa2e5e493502958b5e1d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h168b88382f65204225f3b90cc93157c33372ff1eb724fa1a746aca33f8daa0de226f6dbecf8a9a83af23f84c02f96f78777fb05223b148acc57098aea702f449c71f822cdd7fb499dfb6fb5072dd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a0364fd6de6c60c0fe00ef23193a569d58805a60aa4ffcd89aa03ac2e3d818579658a6d954b7bfefc32fcddc80eab37ccc6ba39177802f825733d3c6d51491d3efc2131848763dfcfece4232d36;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1515da5c8b7c481e7dd3c8f14982307db5ef5e308d480aad4542bd905afac7d02ee206463f6710d1014025da6cb413ac84423eafa0b2d1910e3e9458fec32ba29731cabbbb3483e253162da6caa19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f79ee740d07b2062c494345a585288e9e0451814f43d8564542432e9ce758866fdb07887266f94ded9fc595a1374d821411219375f7e11503c5b33eaead66440490c8187259ff92d6dbcf22f344;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125d999693400daa6437d0ec7965565074ae62cca1efe3d3e39b1b030f54ca5f6e8a0caa0488f8d0c21b1277686a9ecde16cdc768411b33726b9c3cc5eaba98ad85543329d6586222d91312708f05;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h345895e442b910eab3defac166dfe7d5282c727ed4316cc743cc7af24c7214518ba75b84c81e045f10bf08eb3ff7d12df6db08de0b8604b6189fa47f113b7409c16f4c164b790865f1145b63380c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h766c310be45fc928e2acb96c8e7b07ac7d78e71c3b9f763a453b0d3999fe9204191b4c582f02f0e49d0226f5316b108416df3549da142c023e4682285437920e63789cc89d8ea11b845a5babd83a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d6ab76f704ac7a4b68b682871ed4fadc90406bedfd396ce73e0de2fef52cd5bc14a887efdf020dee13d60a56749fa54940bf4f01340f8c9100e25e22605fe177a31ff8ec8ed04d9447b43c9f11d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1844edfca43980150572d71c39e06281db2a0c59395b6fb26240d678727519a1d24aa2b584bf237e5e67a68f1a10cb2a7f1aeff8facacbaad47f90507d22a856ead7305be52fefcc8f590dcb47e6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10896345206d86f00cbb909dc91b532ceb5927f7887dd42fe516bb479371f5b0471dfc02682a9a577649b1e191f018c4fbca12d8b37430600536855c462281358ba374686e2e51366bba276e1a5b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98de49963f1b921ab398948f7785238c712e1127681095330f878924691fefe58795b23b1927fa38b4e73069a3395391a3f48525e4e961300c9065504179e18a697fa68a506751c0b1a6f45a3bc9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h155ec7bcf7a6d354a2c6e920e8d681e2db0fb951358ec89d336e5a4fe1d8a47fb6abc87ce48606507be652f6f495ae145c4cbbba9efc2593f43751bce08687b99c9eea9c1533805615c7e5eb8b0d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12716adc4bd4817321931e05a94f8277c5bc09e6ca88bf67ac4a391f9871edaa1410d0e0b81f5558219ae59b2518a399aae3a914d93b1d05882f94ffce7d5a84b47ef16bf6aa126533ebca09ab4a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5dba81ff685f4c7823c3d068070e32a1d9425fd6bd7e06567b6f02483836f5c9e7a5500c9814ad0a5b2fdc0842f5a292018f53cc79db083ca590d5ed3f0e111bbf31114160dada4502709aaf126;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaa19e9976ef3be4d9e2f5a074f6a7abd28cce3718a75b5781ebd8498d255cba889093db8b13a8b2aca140c82f39a0c6ada70ba8bd4d60d62d45778e77bc3d58c6023fd66461a609573d10f9f504;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c2a3af6a86bc27576be6f53c4a90852ab15025a4f71051a319e028f9d252eb5ee1e154a8173048c47c81fa4ff00868d82ae7bded3523a55929acd9e50df069e54080b2a75930dbd4f13ce3f34c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da6f3c22a11c726d0fd52bc46b39916648b4ff33802b6da07a117abddf9bce1a3ad624309f87d237b5cd4634c75044f804fe08d3fc4a72a09c6beeac724e058af4d81804e60de5abf98d127e3b9b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16aa4f963e254b20fc3faa32661e90f3dec1000e0cf9bffe3f974eeacf6a1e3db6023a7effaabefbe85ecc7ebb4f288855513f447442d6db6ea2bc6ba7e85b0128d751193790b5b9573cec2ccb07c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111491b0c255339f73d586941031dc8e9cf19337a4f80e22660f9abee3790e594e0213843605224edf823d9b84c824f89295a897f7d6caf1e99612ac1092f4ec5a1f9e8a150cfcf7c7af2c41b8da0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfdf318950a13872a14fc3b588428bd7c75710671b08e3a5a9c6813d94557dfcde699e8984fed8b7d3de841e2570348784b5a57bc0064664d1799108393154089e39808fae7e7b173c2004ea5c67;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130c425a651d6023a6ccf63b562362b063f0d3d56f616374ff2377c142d0b0a8d84a7e4c357514ec3abe059bd83fa33edfe39dbff0d9004e72297e9b3dfb0d440ba47f996869bbdb091e37dba3f93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d4e97415ea567bbc40faefd5ae36117fc1b3b8e38b6ecc8fc4f94fdc53c87fc300b5c3332bed2c667efaa22a6bd112ad463359d1f9a7d99626936f9a53c0d516148bd720105a47129f9bf259306;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171a52b62c1ac0feede9f3f75707893031d9dd692e6bfb0c5e87a15ebf3cdf47832ae3ac11789ae3e99e61b5167a18dc546b040ef1a0a53e217b576a23603de043d397703b2291a124777319809d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa1254398f0390e77917630240aa686183ac12670ac0971e70fda57a7a489f1c60bc92f5a1863977fd6eb166c1f88b61e51b4cb2ea049b89b337c439a2be51863f10517eddade7fe247fa7a5d30d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d06217f78e85e3e81ef29f454238307cd9948c2ff0ca6a253d2a37ccc6046b23cb18823138c0288a80a74fdebd422dc05f839020b7e561064a6a8c23e96a61a87111c1d1843f3f20160581315812;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc57a320df3388d2b1483721695e830b2b43a48bc919291d2b36c1294c2894c60c3fd8ec45716ea2cc4926a246d63de56ba32d4dbbc8f789fea3dcb03b727225bfa800aec127d652f1fa6c3161dbd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h661e8239f1b786e3c1dfe9b346dcf1d7e3caa386309371b311e45197eeea4402add3496ccb66aed737434b4c50054dbd1169e698d9c93fc31e71a88393b554d4f34faa02347099cb2138e6c6e740;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a06882ef2ff76329a1773e606b838ef6213b5f8a42618acf4977f3444c1389d48b55e9a0325b18a1cfbdac7a6f4de13037241fd4442330f942b0514a7b0c30502222ed585d4ffd0868b751cc1fff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d944cbc8dbb5d6b20c6241fb20cdb0dbbdd731bf25f6c5d3758c10a0345c0c1faec004c16c0e5fc55018e58048c9fb4082cd48fb6b695c5358b743737df4952560e22ca6cffd0dab180d7ea057c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ec8bd52a0436da95fb8a36fea64c9f9d28040989f9cad7c718516858ec266bfbc7d3fa35ba8b13b3a27a1190c6b449f870ea3eb6d03cc70d9219e332e8f084d06d510c4b2df5de8d139e8181503f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17adc018e1a224c19305c2e47b800fc34de0ecd8c7c70740cef3ec276d3b5ef0ac4f7bfe39e5a48d02a74784c0c4155e1af14888103527a6c59cb879631473f49455936da1ae5c4b1133ec3e926d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d4fd42eb57add2dd590774e35a619ec50241e60d0a86fff799258fc66f495aa460bd50422048ae8854e14779f93950b9b928d02cf4cfa47bdeb02224c881ab540eca78171169ccf43fdda6ec507;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9cc670b906d5ad8cc26b9e2a6626293996d6f73caff8cd7224be5280b2ff520569eea9d26249fe82315066ce28478656289c26737700302d449faa2c1093efa09e6795ac8d68774df6102d775e9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d74366d4054831dfecb6bd65c78c0ae1a7ae6edc2da32c79cb2a75d44d3db9a8966bf79b51191ccde6d1096e0290fb4cf310d7a0bf8d4e36943d06758f6f117397f1fdfa541eb3cda536c7f4dbc5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d92587d62d3fad58bf71133449c66d4988271d9a5f5bcc9a5feb5e94a5faa51910c05998205f805cad61e7eb3ef7a56f8655f143ebd993d31cc0c8ed8dc886090403588577e464099ff952c6185;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1926e1ada02034b178e9f45924c733651fe5cb274a4507f3018ad1c73c11a223fd0a3e7f46b3edd96c2cf803601a0544da63712c52020887eca30a23383e47822233e7dc39f5ac3a9df78556e17b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab4501f49876f849b9e0ada2724cb7546838f3b3be8cfdd24fe46e3203594c6fd661d0f35b02fd27f56604ed1598cfc4c4dedb7a96386f9bf973624e528400dc42ee72286949cc58f1950d2702dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9f98514a7bb7a48c5430aa9f9bd1cdd4b6d568fed1ba403cc0d4a5202d81e8ad6907421ee2a12fd82d0b9b02cf67cae8a66334aa30f914cd24beafb52909335b0fef09cabdf80fbfa6cc1d91755;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c36bbdfd1c42d0ec5ef1d119fe08390d5c8ed6c559aeabd0d4d721f929e7cdf0c72210ba6a298197e064d7d9d95a1b1a8383ae147c188d8e3cf3eadc43d3240a05221687fb3a556e9c19dedc1080;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7d02cc255dda54481915943cd84628355adb46963b9473ca3f40f060f3dd650742bb8d9c6912f34f8536bfbec933b3627737e510c392ca63063367bff7b8ce1ddb4b5ef3e3fc52f334bbb0b58f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10134a3a63b8dccba703ceebb150b775ae5edeab9f66a4f0b5ed81d9cc9412f8c274903491863c8a49edeaf59ca1fcbf3947225f49c20a1723ba51daeed8b70d0f0accb0e3afff23910c8c44f23e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa4e24fa78227493e83dfa8880c4688b0ca1b02ffb3881982bff2fbfd01dc72be95b4b4e5914b1951fb731b2e15d59ab73e40179bd4206e53a7727c497a15c971db03d3cb49d3a75106c5ee3e9d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c48081e3d5c4cd734e1191d2bf52a25e4163ee0a1fe755a9173cbfbe78a69e4a987f0701a609002c464b193e1e6e529a6c4106b72c96eac6ba013b8d877c0f551fb38090fbbcf899282a47810cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h184744f6e88173c55dce0ceb88e62a0d0c5a4d55bf4f054f9c93a43f8f6649b696452f4bf6b3a857aa7000878e476ac474dc5c42667919cb7cec1ebd07f876bea33ec9b441d58c7ee90d9f31e07a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d098deff0b6a3a96377882c2b360013398b1aed97c22d72db9db2c81a119f98059763910a660debd12fbe581a0f36b325d41ba00b5d40d94f90ab15937ef90ebe79cafc3249db2b433f346a2904;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h712004c3ff167e7ce44cfe51d40c95566ba8f2dbeb6c126f908524153517528fede69cd33f5e57dd15ad7823e76e78f05c158d82830f02d208f9618ca9a525b3aadd49d79e6d64909cd0b0ed25c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15da8e0d03cb381eae970b9446d4e50d72aa974d2e8f6daf22a566bcd64f617c4a9e65843b47fa82dcf55e52006b73ddc25b2b9047cf4584c5a47f8f8c17d23f460e5363751a69dd50ed475f16c08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8809ddf949ff879f820167d0d4d33ae688e2c5bdecad44cbe93eba7936b03494cbaf0aeb1f0d3e0c5f669beefe67086b1380430bda071a9f7f11228b89f9c91f3fdff9fce148f7ec83bf1b958267;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha714984bcefbf4d939d107819ba85cd80cc9366c97a807e1e15e344e18434a5895e2dd957794fed96689864529e17f55b3438cdf6aa27e803e04a25d357a05e239a6e4399bf79760b1424ff6c2e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d58686eeba7a284c59efa94e6927bf63e12b4cfcefdd3ce3cd6118afc18637801abc70166271cea7af1a3917315518b0300a934e8cbbf9d334b437e70645044d36b2bb894f132cd4900806e55ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ad79b0c232ae4400fb3d4dd1f54fbeaef4fc7485216494dc9b37a84b387106e4318a5c769e269fe7a8e800df52bbc4d19e8d060c967cb7387e2448f893d3d733174eacdcffcc2ad8dd344b2a860;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a80ee3eb23c2b911d33146b614c81f84044843a1965ee604c59f3d5d6f31f03373e20435cc3dc16879d8f359b5d5496304a9db6b00cf8e384fad67cc73a775eb2a03b25bcffcd54884328e7265d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha1720034d1cf4bc50ac487dbf35d9259973d289782fd07cea122db14783df7039a403ded2686e8cd93b86ef428376f19e90c85449fa3c0059c86b552b85e9746fc89b7f0361466fa03a1d9efb9d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hec054081cd089d307c05993f2cacf1270b3586c7b642a81e8e8c4d61057df19ee1608e21610a24c8e5070cef28e2d3979d567e2b9f2df34e2588c970681f61859680d8292c95512016dcc5dac1b7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1029569f14a2c592a6ce358470c98640993235c478c494c0fd71de178f4aa373512f11d96e47ae4c840d29703987bdcb9cd1ec0c7b0d2c49525854d740473a869d7befdea417e300aa2277b50096b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119e57cf4b14da9c42ea5c176814c584faaf5e37f5ccd3c5434d95588c90714eb47db2095a2e7f3d0502824db20856c681115fa0f32ea36d6670232a3bbb771b9896a9a9f20faff1360ad2c3f7ae3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17213242d59b3b57084808731421b2e921428a85ea88d6723f0ec5e46966ab1baab6b01730232a31023f2c2eacd113bf718e0d0b8c42cc2e0fd8ae8b741370a4f461896adc21a2ce763c0d84c3344;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112fcd35ec179c30ea00c7cc1394e843a384983f4321fd20078ee5e7c5856b1bc44f55502c5c797efd21abaa83997f91c3a9cb3272b0712a317a1690f0ed526202aeeec7cfb631b89a7e54264a951;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e0013e73c03d785905df541feab60dcc77f0e16ddca53654f4dde254a1b70778d72aaae79485dbc138b258b6acbce0d9b79304f9c1267dc524f7291a4b63cc31132eeb4999aa416d7757b47233f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120779ead4fbc034773609082e5756ac6be8c63673731d1af10482d12c8aba9c3f49750aebbf8f0099af342e8ef25486a6f5f6559e2b2056d0f565e39d94b187104efb1f37c304616789fc7489959;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b2b0027d38af081aad37431632404353f600a54bf34e007182a2875f6965fd3e47d222d6eef20d18e0e48bfce320f6eafa404b17801a387351da504a033e7be728ac02a29f1210a1e16611184b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48794c33ceb90566cda4027ad05dbc71533ced05e38ef8bdef46e175759adec604676f72a0cf6fa2e800d3ca356077932a00c8bbe4b563dea0d2c57d62a8b831cf1cd1a37db35871c3dae1dd912c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167f1c0802b0e8be44c79bc375859b72fc81512fe784e12d3d0496c59bfe18fb80c6640410906e5a3914c29e6fadf598d036657a052e4773662027fa8ea228ff8d27f69077692765f2781b193e3dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6eba0ddfb78379d30fa8bb94b831847310e8707a9802757a5796cb5b043ce43ebd13bdfa77eb0da507192f091a9e94cc537750011f153e54502a03c13955e6f1b7717985fc9c752e02ba995bbd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h721912a81c9c705c5d3a6068b7333cf4112fa5c9700bafdae3461b381085b3b655b8184bcafeb4e0c7c6af807350d50970f09637eea1a4d8cd6e65c25e674e122b2eafdac3234471c1bb0495dbbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h245db9b2042f44390100719dd8664c92a138df95b9513336587ff379c6aeace398a4382f20ff092722581d35db3cea2954ddb6028637c94df4cbf75b620ec24ee15cae2b81c1bc9e044dd4e5edd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150fcca70dfca51eb7599799ef2495d9c7a0b764ed39f3efbe9603390d45ca1d0c7e57f85bd6f7297ecb6f1d69a1ced4290d66fb1daf6d04c9792d42c863725157b0b2f730a7c0921f54d0ef8f6db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150ca6c86cc73171b26ec524f9c12857c187627634986c90761d19cf1cc2d445d2c19795a38edc8e2c6c05b578b819d1add97c7b63396bb5dcd60d0d8869962285b1f7d18c61e44c516258b734364;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2fb1702f7e5ea359273f34d63b5d19ba434fa601d2975a5d382bef3cf7f96104e0afb770067e07709ed646d5edf41f444cb34b41e41a0c28c864829d4b6ed4c3b6c54a3fd41f8aa09e34d04f0d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5e205260122e44166aeb61939e8f51e613475e3f2839ebc6408018e5622fb44a33ebc6374852d8363696f2d2a0e6ad03e28459556c7766f83f5b2aa14462e01deac2d371c2909c797bb98eb8f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfcc0615e3cb554806664bb01af9fb02acb732f88a45bc3c238e6516a07fdee7408a188457f9670c57ba37f46b2f8507ce1256bce784fd9a4279eb1d7d2095d14bfc9c12c1e314d0a6cc14e510724;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a8cb0c411ba7521ac2d6d4254a7c9924663584cd62a551be47a2f21fa1b3f55ad0ada7d4e7199f13a634cdcda3d75c8007598a15afacf3d030a65667f8dc7c26cef17aff04033533e880b04001d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e68cdd9e09833a3ee74bcdc56a23402eb33e33b0447480600a0cf38c00e52d7c28e82915dd509f70f37fd405995303e7968fb88b4e226c3140a03bd69be2ea4173f6958e8fdcf39b661d68ec1bf4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8cf925763f46ab43aab3f979f803b901443ca608ecca881ac87404a7a6130ab2644c27e66224bd02af0e2306552e26bc12526716fa5a0c54f064f3e8681a479eee5da507508bba61b34c98d5368d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bee01c7a06e8e5cb79125c75486fb9d5b4a0db57c2b3db088650c0cca5ca7a0d0d7e9af25e4b6fc1e00f56c62680562b82c1e23afecd7ea12e2375336b8de1c54f2238dbfdd051a74e614bd31d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ddeaaf5a19949169abaa97497ed864748d82804fe56da5d27e87abb55529aa9e3c0a90c93f8ee9c0de7cd4b9313229a52fde4815df98edb5ce258ae04005ca02b337965afdaf2c9d80924ef10ce9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1866a9d0125ea61ba60326fe0f2835823511599d06dd2f9194d0c762510052fa540d292708ff4b48f1c3b7a928525c5c25d08dab5edfa874c2e17cc024db020ac9f41165de4318f5844fbde8e1979;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b5e3932db906290286cd804fc61ebf39ec9a3ef65c0bd3c9d9ee1cb434f0a4bc0e029e56bfd201052cb3e3b54fb9973758fcbc1399df29751688850535c4807d61cde25fc1559fa75b23e73adb0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78168eb0d3c0a4b63728ea10a16ec8fe8f1b9c1326243030b6f63f8019d89180bae9247cd70308a5777a47410aed8efd8b991c21f276e8d413ecc2caca6c3e53649aac242661d448833f50a5388f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h568c11683d69005ce7c32e4496a4b27ef1dbace8cb7cf705fd8258cf1c5d9e6dadc07de5204477da7ab6b96477c210a830a4bb0a9b39d830ae12b0c1ef0db8e5f3eb88b65121ed9790f0aa8bec65;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f30f82ae91119d09856a56da835cfb1591c5f5f0e3c260b92db47ce54310cc1ef38b4d07404f1afc73bb6fda69d1cae3486c5f34be28ca16ba5b6cafbb212efd1616b110cd3111e3ef5de6b8ddd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f9b49f2ccc5bb52a21192d31436dff301695d6366e406b7d50a24700d4a1a84f789c7076c796d1015f8fca85fde38ba463d5f06372ae323325370b1d8291839b7540339a78bd91185df573e8483;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ce6f535f5f4d082ac645a3d7131e47197f104b5661dd7a33c82e58f685c3da03983942b16c0893b89b8e621343aab2ea541f80683e8d25f4b62bb406605d80c14bb25636b5ebf3830f79f3b3b6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b357ea047a9d60760511b48c21a243058987b7f41734b9af2a2c12028893dda4accace1d42700cc9c65e642c51e727341853aef4bdc0f46202eb11e7682706438f2a95a2aba7badb7a96069d945d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92a55a7a101be0f77346d5d0a63f0d9dd323a367d67cdb7d3dfece045701d1387686032b37a8e4c48e92251bf56b175275b79e943903557d29eb3865828435a301ffc2b959d7d4971c0b448bbfe3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34675fbc82efe409e2abf251d4d6bd1adad763a1f9247210e3c59c7493721624ff0f4c246317ee1b4f31bd872a2984894bcf6d2cb01cbf409b266a6e1e8965cfef56e9befc5a1fe8d2a649e55b66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120272d64efff3c0a9ed4256db0dd4629f8d34369efed18fb69ec4c90a25b857ae5656739454b0b1f98d15158d5d6d6efa35b4cc500570eac291365ad5862481759e8bf942bdae69dbf3609a54383;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e55ccee95f0bb6aef938b3d9abe3a08d86028d9c67d0edd52c1eb231a2bc71cd951e260ee7c17e1c82e588c5d74992e815f7cce83dbf679cbac7dc4af0697e8639f283863fb2f46d2411a16f1cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f57d9b766d8a5fc142116a0139563613cad27d79ee196d8cf89d0de78d025bd56c06bbd17d496a96a5b0575db940a841633b2fc42e763bd25fa8f58732679fe0750f33e5ca18626c5fdbb578023;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17713ec33af3bc9cf1e09393a1b08c420e6eae6bb631806214c7a92487862b5f2c6b4bba8c875947aab917ca7d74c9c1d968bd73033db4335c8bc511ff574b0c41922ece84817ba95e583e33961d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a1155b844b23d34e82a2b49012a5d7068eb82dffa7143d139658eea88feb3f445050bcf577a1cbe0bc63c4676f946f91262b823e88770a738e8ff0baa39e4cea5494f44116d7e306f8765fdee34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heab7074ce347e737e271f058f919c4a6bba83d4e49cc98e8c46370fd2bce7203f85bb0e38dd6a6cbeb9958204ad84d01e606b4a04f8bfab319b992baa66053711db9c3e17cdde178b443d32a026b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h113770ffc71aff225801b81634ffeab75af689ac083b22a02a3ff75374d30569d22defa5fa7e9d5ba2a5caba459ddbccc312eddc5d1cc987057af62d4d4b0019d96429ba12b7a19770ca57023ed10;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfdcc7aea6e726b6e73b8b51856368029054bce0de801cc773440d6ae46e5069887da60db872e996dc030890fdd3dd4d7452b720592a6380ac2f5d48bbe5275ff4d3ce0343f010bd48d8bbec12274;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb0df32badd3e7c51e2b14b778c8f7d0ce8c50153a47dcd19e6f1f1d89c281895f19c97eff19c6d212361db8bd7aecf2423d680cfc2ec4362492853234cfecc734aeeb469c59ca89881dfd7726d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b4a03666dbcf46648f3d73a35dd25dbe42d0bf089993478b4e64f4e6e61cd4b3a614d9665c7f70964d9c77b05d5e41ddb3d5f1a5778df17ec0c78c74a3ec881ab8a499013ca9ad1abca4b4cdf56b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1abd27289a4568e95e8129747cc5a934cb85a918608bcc84281b843fa6b92a2c87166091f2b7b36dd2ad0d229dc0fa4a5f72d5604b4a16851c0e1632c6459534193875cdc72fe9e1832c595607bd9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce737873c4b2778dbebd47fb03ea2ef6d40da071f22283c33a45d7d51e189b0f396da5ca17a4afbfae276163271ffcaccd3c60d54795a030f3abf2d0ead210fd45a5f59e21bdc844550f4a750caf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9917f4c115e259abd3ff9ec371e5410b2e33d8091c7d125e36187912676b290cdb5fe5903d47d06b1b97081bd3482844db802c33f8a64db1f5cad7488851202348cfee91ddf03c931ff6a2707552;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2af6a37b04fc0ef403c256074ac7e0f333aa00303b73a7f63336e030cf87c59a33908b7f253259e750e34b0e4cfb0648b1766f0cf17ba1afe0d9487d9b64c5f127b20025e336867f4e936f36e02f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112cae07c6d1f6fdcf10a5ee09c78992da1c815397641652c24203d88b57dac8476a28492d709ce5bdafd16ae4231dd39a60660ad164f6cbe258f094b524495719e6181258a8ea043e682c735f7b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bfdf30f170c2a2c2a1dfc1bc8e966f7f59ab2ee6f0a1dc4999cc53b20c67632f0a3590865fb8514a60bf7e3aa9b5721dd7406a16b2511f9fe7658ab4502a53de310d87c7840b173a89f70aac911;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h61c7ca0070755dfdf1f53bba2fa9d2eb8022915653a3e38715a9a37cf398d9261c40337879aa70cf1e1d27aff60835e441b6ef48f195ed9a38d9a7dd3feb71e4fc7bd8bc623f8ee80ff8e79eb4a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eddbdd6582f94502c5f8f9edf345ecd7e5b7261c93cc5dd260d4689a1cc3d03394452d45a8d5f69796f2ef3ea71d4151866963124601443d672f6b5e002758d5343192d7f652a1410b35622687d5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac34aef83ecfdcac9b1c09ba0b9c2013f8a7d277fba62fa2426d407704837272519d8ab3e3dc89f8bb9fccdc4f109f3fa81d44b99a975275db547fdba96c08f98f0663428e00092b23296e343621;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75e0387a183d13cc250330c2959be1f839e1b1bf3438988d00c9f6f6fd95c65db271a30f899f0351fd92b98512a8ad2901f82a0515a258c4ad7f70580a82c19dd8dbc892d8455926ac56db3c3196;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h805d6c3c23a4a242008cbec75e34b6d51ec6a2d854ff22be3d5435411c45b857b956a923d15f6cdcb8fe59dc282eb6006be3402fea32c0b66f217f6f363cad6c145ef4a50212a36dfc28cda3cf30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119d89c12ab9d3de393ca3a65aba8cb21f638724b8f142026bb8bf36b970cc49ac39a790428f7d68308349dab3b4205a5e06f6ba625f6da54705b371348fa5ea45746d256e7af887ce4a7130762bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1eb6d03648587e49080d41f75867722f1fbe7f2053d5f3ef38abf13f7a9db0bb7c45100614c5c2234845fc50853c3d2b8bca69ea5b9a2b1ca9b361f1335b3d99e8e7f9c4965c89edaea978b0359;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dc6bd471171ac97536feb9b00512880450f72c58ce854ce51bdb40dea60003603681ddd2331cf1147b8d7f5449e80c437f04a9a6be8df07a9499013985c200d2becdd9004dce80c2ff87e61b1d60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6176c69215d89500c2847b5754371a101d915eb339a0eb824a996bab484f44416809aabf625076ec452b0d4284956d8ca25ff8fb0a33277c5b6b511a8a0897c111f348918dba7e2a4fb7f17b3cf0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1743bb9d510139f12f7e357851a1c30fc7269a2fd40f36adda12ebf2cf7618c0e07588356b4b5dcb506a3674c80710a9b4e9abcda40f500cd553f0a6648961ce2f6e687cc954f69457fd1d4d3b917;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131506c4d2e4fdfdc427ca3eec8edc34aba8879659adfa4429ae311b39d670fefdf95ff71c555b923b4bde4ab4baf409b0417976c9f1d0506c1ea1a6d75902aa50b8d8922f8497960a49684a72e50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9d1eb583608bd1ac364a047d208f182c01a7a00e9c96becb107608eb67827575294383cb4d90ae90dfaec6aaee88e825549503bf5f5b1668dfbb6f3fa8ec7cbcce83718d6078157c9db58cf33ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ce75c0af7ca0b9de610735adb04379d976c323f96ccc2235bcea7aae6c07cc4a1975f7620a6a7d740e28b1e0c2aed95b879c1e0cd2fb9e902fc5be2c4b3e8635c0d764b8e4d2699aa35b4a6daf1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha11f215ad23704ece13b49bd87310908d0d0cb3fa67df6fcf62aa5e2ad4a28ee2d520868cfd849dfc9f5e82c65acb79d33482bf244af3104c86df15f5154a8748b4da8a80609ba35fa805346981c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191a7905d46a82dd61f3aa16c422052f8998194f4e6f6929d0be51f9a78132aa6bd6ad88a464d6b3e1552adc4f73217293c1531d4111c847a4c74bda43e2b28064592c808cd03d93a6de263cacf01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1944b9a061166b31d7b29199b3547faffcd163e753ccf596b45235f2374b1489f9229c7af44462c874b8ce4e3a46f3bf84e4e5af332d340bafba698bc4020fc3e70f572c6362a894ca4824037067a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1847485be84628372dc71243715a02b2056102b8b494f130d57cb2357f4a9bd698a10c44afbafb140763bc07f958e27b37735c349982293073f958be251d27ad3c8c37fcdea31984e1736dd27ded1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h60eea5b4496d25d998a1ab2279b6e2ed18cab0434613de543714ceb39c53aef060b2223bdc028ab9da4b2c1e70c17341170ac31f70a2b4c45a788c81de524dd3a468e7f31f451335cfbedf5a4fef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b27f43feaf77e2a8c5c412a7b0348e2e25091b1a94a5617e76e1afad62263e5b7605b3504f40265706fea1d592ee37f4bdff9635bb0a53fb6ef5547cc9ebb7b96da7af5a335f59d15f419b1fe3f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114d83444455c0956d2c423a7899282fccf32224b4400612b53901b34530aed832855cd5e1f38e42e23fb2fc8bac05e251b02cedb3c822ded71ecd2791bbfe68ea827124a94a39ef5aa7aca6acbaa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b82e42f3338d4a0de7c1faf389672313e2835f9e96256b6dcba546c10ef8289094336d6047143494abea61472c12ed73f2cfbb13b28d030bc61473e664344104d83422aea9d3ca65f48d0c4579a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e61c87cc49f54ee9fbe7f252d91ceae0f65a84d17e0f8e22c7afcffbee2fea8cfc61385723b34bc0f3833eb7d328a8ba4bee657de87b7fccbf55f7a87cfc822670580c37ab1d1a85eac9cdf7dafa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12323c2ea496e1016056e787172658eb16c84f3b0df37b2575f8321fa428964b5f9ff34b67a726b627412de0ea3b7e6da8960a04ed52f6f93ef86376b058d3582eaf9f0e93337b16e96826af1f285;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a44e44e03bb448cf431ec9ac45000252e7be61ca888a30dedd0edea41fe45e1c439c9d604629cda3f238d63404199c65cf8d1b756d0dc1348e7cace127e1eb03c50d05e6676c952696b282e3d624;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1182b2d7a02a1fe8ee4886f54361058c5c66a01afae52ddf33b4563b5fdaa2edb3266562b9f04183e42e03ef9812ca42223be20f51e6477d2b756feacc2a230d061963e006aaed83db3a454a3eee6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e430135e3ad9788d415fe7b8e7639736af0deee9a97be9d119744e6ec719a7723546db3fdf5521bce7177a30f3a638b9e80447a3da70c2befabaebf50b29165d88ace9c82b2c0473e96cc9f62bb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da8b3dd7b923d4528e997b5cffaf0fa78175cbdafcc3a39b9e40821d762efc28012e26513b9297bec9d39e5520ec6cba7727f459ff4c4bbfc550d9477d12700572c39ffafa48c9e0fb907892d996;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbee6bf96b65a931495e316e090aa20448d0d4a455f053b3eb58b7388cd8da9f4196237f2757d45bb75c4856c0b141f2d5df964f744273e02be909562bdd7949749eebf925b1f47fb3334dc278848;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fdde50ca47d6704889ed707d5cb4b646145e02b85ac5609971914e425ef2393babbc78c501a9a84bf29c0fd982cc03e927e9ddb7c62437ee2f915218508609ab613e656eb824247c1f3cf40d586;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1243bc272777b3170ff71779d197b2cee02aa3517c298442b82771c592680d646f5c6dabedc1df2a984b054fa0375db0aeb46df860c6ee9c2b21d0fb7b7daa3cd51f2637436626ee93848fcff01c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ab16463ea2da7d07e7883fc17d51803ae551025e9d3a04746730f927e3d0d124442e2289e772e8c90d550b81eeb37370c3446b0e2e4ad3782ac608f75962a4b5f5de3ba54d2ed442dcb73353872;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d962637f96ed8f42b4f0c53f97eee794a543387ee53d4b7136420629d4221d85631b43052a59a2ac240586e5a72532200557620f76e966f6c108029e3de014943b6378ecb0bd32d434d660ac3873;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82836e503015d0596e9017127698370c6614948a8f50e37686fe7da36a5bbac16a2138a3a5577b5055aeb3b277547d4acba3c0dee05e806c8a60c0ced2828a780553b44e3f827ef274df290aa6e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16700704242149eac7d6d980f43e2846774ac15d446be29b8f7df15bd004946e420ddb5c70aff84ec736be1d067c86d8e2bad58206182f20cb7649acea8693cd864e791a57e91f67e3cd39d6afd22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74de2ddf488e79ac5bd94c0ba056612e63cc360c55389b6c5d9725fc41396078d693688a83febfe2af921d75bbc83f66d294c34bea1b3d02adb447e01a0b17f1bd2a71f1704cfa8cdaee1cc64996;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd4fde19deac38716d798a8cf80aa1f2a4877a0b1454d31ac560761dd776c198b8b4ccd1ce06a07abfb70c32a7e848079b726ae1c7a766924105d3fc93281ce8628e110cd3616ecdb50fa76f2b864;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7be27f15316723fa80bb06c65256efeb77c35d812361ca5681ac39c53d5eb91f7f24cb9ef5f6ab853f8f3e4d9e7e6c3e8c735c456c55088fae291d2dc7ddbbc4d6c6b921c6ff4961077267b269a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d121a0552f6a100ed04918db9c75ac73ffb4dfbd0a6595caa9aa35b67eaaa22a8e8d9198127901b17dcb6c2ae66f107d8e43aca1e40792b4e640361b900b7f97440bf7c2c4e634e2b5b89694fc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c25282bd46c6e9c52d935a0ccc420a731f3fcd791a51380fa7cced41524e02d01994a4216b1e91b93e77702db48dbacc3a80eaa28daf1142e10c1cc7a07abf9a8f8e9e535b26d8e01972515f1a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5c39e9331dc9fc0eb4bea7c865482e340529f7db70ad359922b7369333ca27b7d4d77abdd1b3856262c1dcb47e7da224b9ec1d374b09b338db69d64e468f676964ec424effd917610b113b4eee6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5fd81ee46fa385c5240f66086b5786b60fe6a7ca0772a88f7c53db7b916a567da74d15ce2c34cd8f4af0360f4d3ee32f3666f2dd01cbba6501e836d068b8cead0bbf230bd43f80449f2958d44d8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7303d2ce54d7134b5cd05e0e257739733ca5e3b66ccaefbb0d60a6702bc12e1334eed713dbb774eed568486ba12f594c663603a0f5035895013e4b472b9487dfc0b7f81ff3a542ad993bca8185c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0cf26b76ab9cb2f9f8b0012202f64d9aa99e53904e81919ecfda2fc04217adf09c7c0b9f0edb75259cc6ca6bef574bdb9d38b424bd64354f1512403ee6b7fc33cbcefa0eee6681835e58efc8c00;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb38d0f08198c0b632ec824a1877bd11294c0d910eae6746c26d5ef8b325b40784fd970ee997b93aeae514cb653d5c10830a2161c148262e9a49449247eb859712e55e0544375bdafb3dee48a24e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h623cad36a45d91fb0a0ccd4d24b42a637bf2f14301ec348f029a05eee31f83a0c4b8ecf96db1a658b0cc9cee88419b4fd60a07b1b146813c2e352d2514493c0802aba10641321724077cfbd606ae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c5d369588127f0a0734eeaefe134def8c83cd241edb0209927db6fc33dc6b78c07102ae9be6619553802a3670acb525eb5cc8498335dbdb16d407059cd0ec77add5219887db36e0238ace498433;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187bd1796cbca63c3e9b517ff769b8a401502c2860a12ddd54729a20b9497c1fd80fe1877b1fb4047395bfe36b35ccfdcc5488aa53cdcee0dfb1db88872da304828157dabdcf0eefbc0c969abba21;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146eca0dc94bb9c845f30942213d14cbecd83e95b2e0acb290353931ed11f5439f3376c4359476373e9c1261f0e69badd72e433d57c34aeca35deeada902b0b46640aef1403f56b4972ee33575ae6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cd71c101697ca18f5f10200494020f529c8ae131ce4d6763f679d22dec1ad176c0ea6c1d38cdaf177721675dbefd57eec92b1ce15c2da26d685a88730984dfc21f174a6b1f44b9a600f16f79da41;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b85f4ef389453fd734c1226c7eba89c176efe503f07a526feff5b68a7863d32e9a59c288788dda0cfbc1818c47a771e16cb8b4eb46a7179b5b087ed4973495b3500e65b36f1928b0f5e5acf442a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbee48077879160ae8bdc093059dbc1eda5e529f4467b63420d8f838a82e686a350f5e6194d94af3543715815cf6f855cb2a9a001074ba84eaef3bf78862124df2ede29347b3ce23b3694126a6ff3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b24e71892370e6dea2549e322f718f43fec0669536bd178911fa2ed6974635327d54bd9feb86ab860b406eeec6d2237157d89fe09db371daec980229bd7862e2838ee77bd4caa33d8c491880be46;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e13b5e5c35dcedc4ece836435c25f9558a37a60045c6da7c1004df5abb08694a87007a06914c301c35af412e9d5529cc7509f4b859d46ba50db67a16f53cac79d7fbca18d80683adcd7607959994;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46ff7e771f4fb692ac98a72f3499f887199134e9b2427eef1c8f77519a307ae63d66a64bc33ab8237a7b08ca348d346b4ca7ba5a66712efabf56b40ff5c07f417e8c77a3d5320c6de0a0b4b1e6c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7666156c363cf5d09694420c4d190489b89b81db916ab2cb718a41460c5fa64f3f085afabe5ed2401674c9f236328729ebecea7b2f482ab1a87534c760f5a47206d5d27acc94b1dfd4c10ae1b453;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109e93425d8e61a81028cccb24c346622f9d1f005826565a6f78c77342fef2fb26ff36adbd27799df975b1e1c9ab267312dea661c7aa3351ece78e3733de6b60a69168544b31b3d920089f2579e2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125856ec1149c1cc58e7b1331b467c220d55fd3609f0bd26dcae927b73ff0e8a6b3fc900f0c4166fbd295ccdbf7db5e664d034846b5ff87b8ef24db8a5f724c9a45f3ddc08e13185bae3ccbc1c159;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c7a0aeb17db0900dd1bbfe269316118a6e9a9ff8fbc1471e6a1372e769f61bd2f568093e0543798b91d2a2bc55f48ec01565deac8f0ad66fcf7159d7cb3bccc766a50086fbc95c4e2e8515ccba2a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b13076c6d1be28df2b8966589722370fbe58e4d2f21ba4229a1fcca13b6ee0e4d0158f3083723dba527b799a4a16a556246c037e572436236afcda378c38256e3582f6e46697510d8af7acaef8a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bec479341290b45e0564cf8ed56986ef9f08c8ee310969fa49af2a503bea5ae6b910dcd631ae63fbcecb839c08ef30bda277c7f08f57d6cdad8c9210a6a794084dbf733b8d0accd251bc6f13f3e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1369b8dea79eadf7df03e5cbad1650e6cc7ace6432840ad3d145d47532979ce95e93f59af42c271f22c210e1df4bfc9ac1712266484e44445bd5b32e9627fc3bbde38fae721662231139fe4877c51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haf90c644c12ddd3c5a23f8631fe394d18cf1e6079a81846d4da444dd48db9fa5d3f5a57288e59be02e5307cfd129f0b9d31edcc1c887585a0776afc56ae472238d0b738215f17076e8f8711df830;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c4550165e19e2b8d864d9d0b5295fb3bfdc71f0bc5ff1f72849ab581a12ce1f5f97daf287f080d537cc2aad1924784497aa7b7d8fd5bbccfa1b2b23984968b39bd081e96c0bd78ad03a98e4359f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6d7bd4a337e996f0ad33b8a555d301647bca5cbabd82bc10809056a4f22a9a90dc99c6def76c58959b5d49bdf026c7a61180b9cbd2c77d78e3ad9553b420d133e4a3cbfeefee32566719e2fcbbad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h401b3e67a46f2bbfb1f2a94efdb2fd9e56c120919570ee35955c83360003d7a92486a688ce3348a3b38fce34903cb0e9e50ab054793ceebcbb8a5fd7e713d551f2adb379e52a244fd5a53f386ea2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185bb70fc87e8c2d6359c76b55a497daa0aefdd5699edb774b027ca0642802e5fa7c5ce3ee90360aaae318861990562c9ccc7fa37047fef82f0bd731e03ae911e30d4393f144035904a2ceca8ce93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83d1da4bbaeff50eff9c2e50225c67b1da3f599c8754280607c4d887a8b552124c30dc5edc41c05cbe00e03ed702f13126116fd504fc951c7257804bc7632e907bcf54fc84e9b08973847af7e5ac;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f5a2e155fa22c27022d15d2652279a8024d41f83a21a300744baa2ebe3f3bdb7ba20329458a94aaf98642e28fe9658b5a8a031334c52244c9809d53d95d1658855b30676b80ff89393d70d7b211;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6f4cec418a92dc1861c9bf9bcc35e5976bf10e7c68d0eb6e178a399938e78eb7c49efe4db1660f71f69b014ef8a27f94c9e84c8d976893d06c6def3632722b6271095670ddcbd8868ec111a2cb93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169f89cdcfb6ba121ab583506f68905060fb8ced197b47d42eaf1e448fb6eebc7c9d2483baf28c5125b1114644fb48f67dfad095a3a3caf36bc81e17051d9d22165823d6c0c0ec338b7a72e0fa77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e35c8830eb9d5ee0ef958a8317cc12e4fa2507bad9354522fa6159cd05bc6b72de77d549d6aa5aebfffe62749e2d0415e14015db58c7c50435a125e1d60a93f0a7e59118d7fab5fb88403561111a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc194f5b04144722dcf5d518280261d505362d1ef6b5da50d5fc42d1f618eff438bb42f82504e7ba4f8297de3091bb7cf3cf07404babe0d4a9f8b672ce9e79ed469490d50f4c05386708c972062d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha43210ee424436d9e1d8b803ffdc18fb435615e5b08689576247e8e0bb1df4b8135b2074f4df127cf58ed885208fade04cf114fb539535dbc641f9ff0d6eff94be6612b1b29387b5a5bcfd95207b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b0552b4e20e3198d6860032e9d24ce5d546bbf37516c1c6f3a7c974dda4a23da162ed252f143a0c5f0d7f011afff903dc546a9e24ce5e809074707ca7e8ad62cefa552fac3452d905286807a3d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a70126f6d83580ae5406bf3aa141a8ba67cdd5e5afcfeeabe2c0da01fa8abda676addf537623422c787e278afaaae1b3e61570153a28bedd5c1192b3fb68023fa24112ded5a9d455ee41764f62c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6eb4b3c9c1e5b3b46547dc1bc30d9082395ac097b14419a0af800c43e084c4e3b7a75f3c134f50db0fe7312a414c6bacc6cb6692a7bac63d55703f2a2ef346f875fedd32c671ea9980622f417444;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93564354fe675252a04d759a809566c1619fda531932207b2d0e3bd0b6bf461e79482ef520921f772e092327d63cc794d372fe1a5dad70fda04ccbb6d9d4e653f368ae2246c941fcf355783c676d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa1c8419600fcbea408203aa523141ae966497f23ab7507180780a9e0ad23cc20cafae0dc64b842f60acddc917b54186c9e9a4f6779d995082326e29f2e9ceab41d823a20b0853e0155db457cc42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef1db5023da930fc691b2a852b679a71377a626c0491ac10b9e84315c7e9ceb4703ecdb29037bdd49bdcee9dde860d0ccd939131b9f9b07a2b4f31b2317341eae017740a159cdb648bb14eab75d9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b4e981ac9625835c89a204b59758583bd44c9797d7a8083ae0a8ab6f1ff821807262022dd33dbf9a3d059cd516bfe8fd7f90ab6a493bbaa16a0fc0fce6e26e62a16d15aa7162279716142e0ff39;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d3021a60e770057ae1ffe59122d226452a469dacd38f19d36434ed34e0a1bb352977d62120e3ec0475850237d53c179b45f844cc98ac87ece3b5bdf7e8285cd9041c315b9e83c55e3f81347068a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h669e2b4aaa109efdfc5a112b11a1cc16c4b1f712bec98deda81b0161b45a054463db6063a0ede9e776878748decbf6a1e6c4a9f73490fe1537a916b622e206ae477adf1330534f6766592d19e004;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd974df92ea02ddd0ed4b0948a96ddbfb0241693af983b4c26f30ba3b257f040afcfd56dc6725544d42dffc6eb3b91eb5f1372332c3a436eaddc6889baddf7351a45e943dc66585106523c013b2ea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc87f9b9237173dc7ce70331d4070508cac33a0cf5086d4da283e1ba35853f80da509d01b20435a0d16147715cdf584f1a873bccc3f40af526aef092327fb23304fd257b52baef2672189e76ab22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14465ad55f7f9b9929b67290b6142489f0224fd9ea0f6b44195178ed398d8d8b751005c83af4c153e54f53d21408ed6ea49823d17b708ad1f5fcdd79dd3e3e0262d5d6539010cf6658afda43c5db1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a2e957d2025000ba481e2e38bd5154c67335c950eb65cfc2fb7cd8e0b94b82af10a020f33324e3d59993605c5e6dc4a13784172a67a0e5ff8752b6ede404eb75e71ecc2d118eaff9cc4a17009e81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4e7da9b4cae2ae88f7d7ba6eedfd9edfdabe0dee1804dec0d6b0b6111d8d92cf0208e0f2614aafb450490e1bf029c87e93bc6cdfb9f0232f350eb29a5be2d3ca29072048456f0a32a246d06d95e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aaa5e4f2c3710b21c5fa0c48aedb8138449f61043eaf472b4765a8e712e2323e754aa36ca667c6611ca02cbb1fed5d1d663032b7f43b3bff092512483fdd885087399e35f5a9dc3c373977bef8cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h167efd6dbf38537c4ac7e1374bd72cc0b6322c955846c6ef6281f81d50c4b4100866c9a4d43393cad16c9f2eb59a3bb7ff54fc549145833825fc4ea9bba0229bb89a725eacace3bdc275371785ce5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1566a1eb7b0d2519f42c6dd17bad758f8c48e9b82338a9513b02766347e08a33c533a7606731b491cbf044e925bafd99e04b301cbb7efc36ec1d25a887aa848d8309355f2e11c460eacdee1d39192;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ef221d62031c02c9635ef1a3d126c9a219193822425d569b6bb5eafbe6773750d8cf8051d62bdb90ce6d6f7a624b483f6a92c2950a116ae4ffcb23d34ca298220ed330ace4a639a6a3d43c0d0a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb78bfe53211389ad4f2898d3f21a90da964b7563b12deec23b4008c2775948a50c0d0f3050076364691d646d078b05e00c1dceeba5c90624ffd7ef5510440031c42126332570f5f2a69eb7f25ff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h552690259c6f16a19ebd33c83c016add5d74875c02c636757b3a94ed9a84899d80e8f12c7f11c8a2507e8090c52630ce12fb68f916d21826cc5041483479396cb006953c394c8396333a21a099a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bdf8c9978b5654c01bcb104c94ae5dea298bd6dc7f0252e1fa8d50dc644b035a58dcc6c5a217cfb3f9dd74aaf97d59a48b7da29f9826a0feae901b60188cf4ac3a9e89611acbea1f5de5871f4900;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183973628c60f0faa3150918ed4e6b9b1584ca0f84c74a24ce960e27e486d2ef79508f8938a1d735e13c5d3f6deffd2fbb1b2aa8acaa937855b75f6e39ed42f1c47d1073fbf29f7b6cb1393a36ac9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f933cde3d0b5cca92fd888537cc27d6931d1aed84680543660f1f346b1c07d0691c8bf3e4ad021ec2021bb732feff9dc186b0a397d716d10b1c532b2d4353579bf1c525d7156ede6484590a0ae2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6b7df31f884b0d2e405326c3086f351c42ef221eb80657d6520ae2efabed5c4ea3c1e530e499f211682fc8d9dbac191ec9713887367968fac523179ebfaf6691168cd9d5af24179cd3864b01e81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e92f3aa77d29f391406981cbffd1680015c14f8e43ff7ccf70dedbb3a8e77013bf8e9e52bdb447de75327f91e0cfc26492a70358f7b0e7c77563bfd03e2d0c0aa2c6f657f1d3579e989a78f096c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h100b133209dc0fc55667c0e975bbb6675845290069f963cd9a7cc1881e68baeb096ca04e4a4011554d75efc6cfce9258f3219ceeee7df424102b5596fc344fb158a27e84c758eb2d3584c0dbe2a6a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103beff7711cfad94d365b3e0cb686df3be1ea4601b241d8b70013c9a6d15292fc73693ff49f8a3ab99bc75d82d17b89cdea6634b38478489ef5f9508345ebf8199c83aff06607d3b16ca7d288af7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18130ce43c13ada8c10397c9123efa40917f997b60e88b5227bd504b6be8f1812eeb0d78e362f0de850279f71d0f37392a79ca113a941848929eccee4f8210def36ba25dada4a39e83433d65258ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11941ea5f820a60ff53b8573ab84b0263623795c81895c2bc6fb368bb9626fc5606d84a484eb6d2a3538502bd013c544be21d546f163793bc7dcefd9b3c06d2639e34e0608b295169e06773d7dee7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa7b99b1696b292545433440693e882358e60a528d08fc528f76e913c8c1c154ced9d06afc7f323502dbb420d363b47f43dee010ae3e9b2bbe1e3a7e1326598e99ef1e3294526edf3e15a1cf527f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e17053d156ed39a191fb42a2d954f0ed9813e3bcb7e50cfea6f55f54eb3b21adefc66d767ae77c7ed13564112b67982b01cb4d7664b5237cf49edb892ec435b1ecac96364d934b97e14d89b70f26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14777266fd1bd97341cc287f302052f7dbb54dc04d16c4741c64b4ea6e683f1c301d172d283764819cb59e22d418603182cccb6faa874ba8dcb61866789d97403785b681f5c07d0668aac52a2e2cd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8695f6f247cbc952e2babcd12d8f077b487285009598e1f024e62d964d50c26e3c3d49c5fc0aa5c6524bea21991db74023949ebaea6424034300b538c1c22482b78dec3418a8500013c7e146f4c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he10cd52cf48e97c4318340a2b9d84720b1b406acf6ed49bc10aa51f8cc9467b133cbdaf33d5110ee061a982a84ce744b0a8cdf88437f5775741bd00b2727e41fb080b560a7adc6059da0ab98c2ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfdb1095596b423c214b60db76dcf523ddbfc3a4a3479132686126ed3121815141fe144642d125409e21842e90cf89b2dd37c148365e18bc076fa2c6b24a2d3f62db84b147b9bc36a0b95fedbc3a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0499a98183f0f8bb43a12d1d2f8b4c1a44a02670016b4c108a9ccfa1fa4d2480e70c2698b0224d09734fe471efa8615cdcac45d7c05365bedab115b5b7dd294dabd537b9b0f91c48c6b4439fcd9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3101c08255839139efe0ea50c573876325cff17d1c0d7f5fe21d19f36e01a50adba5b93f6e1e3005fdafd4fa87dd14e8b298599d7c10b54b0432c891978671d99996595117e331e5a5b295965969;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71c5ae45be977da4d8c12943f2d02c77036a14a9d4c0cc6a542749bfea28ef267e95ed5a85633cdebb6632a2b049cec86d03cfb74f25c0717c23c2ed8b38fe9cb1bf6299f39c704ff692f9d4ba84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13728cffd7d0472948eaaa30d2324aad9bfc01a2714c4227cbb1017e29273a8f4e720183cf190d0a86d9af514a4f727b75090f4f1af789fd52c1f2376c0c96ae868df99f3f2215947ae6aca284da9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h51cac4d69a527f737d5a67e4261f6d76480a1285763a3725282005e228d141b9f065ac3b81fc43fbd55bd5f4ff912cde7b96ddaf3c79f334854551c3a38ee8ef50f265747057b579f4bc4e68db07;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7eebfc89af250a0d287f64b0207df3a6d9f38efcbdf9f4198985fbf3fecd1793a02a989b79123312442b73c21bc21c26f376d45d504cb25d3d1b47aaceda55e79044343f8d33484e57c946d57f7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf1996de9572aa9247ab0cb25ebdd7c683409dea39b453b62cbb6663111688eba9e417206d13185bb3cbb1f55897dd0301c9774e51bde82c3b66351a39e7ebbcaf6c75a66761402ac5bf1dabf6884;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1efeb7418405b968996832ddc063885ed330455c98fd0b77a4c1633cfc7a278c765bdd686dced201fe54bf9f5c19421e122db98ecb4deddab12460130cabe6b6e6343adecdcf2d8579eef2a330aa9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf03a37727bf8cdf359498734c221faa1e82740057109589d8f1ece2ca73e1229ac42f8f457f77a64425d4d631cff1ffebe29460a31d97f4047cfccbf249028ffde7558625e7c4187a07ea4b0353a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h815fb424b06a98409932b9a1069f169a723dde5ba188428f04819fdfeef2d2f718cbfe62523adb5f14847c85b7cbf79afabe8ea994a2dc5f2117b214b830312ca4e5d382da3c4f0e477d59e7f7bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125bb04a04806777b0723f44c703da29a6cde98b5bbb5ced2a2ccbcab451e0c7524ed2d3544ae31735112bb7fd7f69c7c21076b652a96f74b4c1b51c8c98571d7f80b91f1b12361258d9dd7e9c992;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd77d8d0cd2d1a67ab278341f8a8c7e6dbd3566b38a861bece95859f94eee2a6b3c84d19ac4ccbe0f11a733e1da32233668275c0a51d1786b878b5d43a0b25de1979ccbbe86f3812604f57f002934;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ca71d8ac890fd76dfc4f5284dcc6536dae2a8d1e2d5d4e8b60008f5eb17fa997f7233b6f8c847e1f7615a257d10bcec0f5b096a8561122f73b329b7c90f3ede67ab178cdde0def7e5f4d09f39ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12badd96fba18a6a25af4f56741d3626f67f2ae6e93fb6ba2330a415e5d55d0c0a23f5ca17c292a6980c64be24e91aad18a529eb82ae1b0a2995bb5a13d75cf3b6aa197d01ccd813d260b592b90b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f2841589c593a2dc410aa577cb11b0fe03fe6e6e730ad5d8067f2439b79eee13c48ac5e6d01aebf027d37f670e3f48c3a0e454d1f7e7bdbb4326f059749fb0376a357ce34bc61a0db8313bff6ef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49bd53e7739b93a20bc6ffad5a57389308ff9e74f7976366cf16a87b1ba3fcbd7c181390f16c873f350610008db53e314241d99a48c236f25cc00ec39d68df8390816d595f71798fec2f19247ee9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a31dc607a3b6e09100f7890c7614f9cc58f34c7c392e1508ebacf5f8857b66e184cf795ff60f81d88ff6e6c18080cb143150699c3f415d5822ad60059e92ed34f26ac60d3f3caf275e178893ad4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35ee5a7839e834646641878d906316e467b2138df6270b1f0364b5800336488b9f39edc9f9f50da4b0565a8086907166e3dd08f54381ebebde6dbf40e73a3a49253ce70a3e2c5dc19d4c25fb11b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a1d9cd4f981751b224b09a954b28d259a1de8940e9b5e09a5f754a592c1f4d5e85984a09dba64b0ebe3c671d360856e386ac83e6576d4af146b183a9289cb9e68d063aeb41abfe8731970e5990d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3ddc096fecd8dc924c0c416f8eae06080a6be1c6e270267fc5e002d479f267e816bc8680e8b7181399118960e89830d65ab1d285c502de55afc049b1f2c567c39b3095b9156518c1e2b7104019f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf80c1b79623bf29c5224dfe3794fc84bab5f598e5d2aa35d751226cc9ab6be8e86e9fe1e42e1f757bb0135f220c74f3ab9c3773c29e3aae90625aabfb5700a2477f5b63bbf29e8c2d769f4fe8816;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha51d54e8f84db4449b83e3cfb1fdc1ed0a7f6f82f8a9f6caa2b3625d7878ee57790ee8b48e6c8f88f309e4d8265bc50d055c44d7c942166d7210272771ace4259b287901d5ae6ce6754820d8d41e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cdca1d4ac0956b2d59e9b659be37fc73903bcf2aa671ed60f84b1c92bb00cb52b34a5dee797eb1a5ba57220ce2e32310ef9e1dc929c8bbfcb1d39084ae123e559e3611972db0f513a0638bce80c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bab98afcc76cd74c7daf0e35f36f630a93c0eee23862f1fe0b3379664fe7e963c412edb58256cc5788d6de38ab7329465ef9d9fd67b22f4c756596d2f37a092ce90193fdfcb24dd5b53c7f63a7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e37106cae7a02f7a7e9c63f41d1d1a2861ff8daacbcf27ae0ffe8dcbe9e752a65380def6ee009da35033ed00d1efeeafd94ccbecce231366155ed9982a82470cc77bb2ec759c5c51f57a62e1311;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c28e08aeb1b9d13d7a12c6e4eb50c594c4df5fe0278090850134ba3050414d54ed3bcb6c3d40780db27d55cb2256b71ed5560cb3db8ae6ff8e8003cd99269c1c62b9d7588c2852bdd0fcac3157a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6e730579b630352d77e550552608ea76341e8347ff8754b03065883c598263dd7cd2e81ac99d5d80e365c48c7a6e14dbe413a766f54f5134cc37ad973a7add004af38784f5a611051533e8ccb0a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b494bf9a0bfa9c2e5912e61205a9cd6519a522df43e3512e504f70a7c6d5fb88394b3491092aa505553f05dec19d047f7a829c54c119bdfd5c2001d780f01154ad8dbde0dd9531ae7d1504fd9e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176ea02ee4ceaeae3ef37016b1a62d943255b29aceafcc33f16e99bb5566b300eec2a9c6dedb513d9cfefb93f8783278b7a542877739fa46f6c1d8325066827c4761a932139d857c35e15a921e19f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h403fa98b7015cd51322f6e63a7d3648eedcfbc72503bd49cd5cd9657b6b14988819e59791116e3fe837b965d9ee0fe6d371466d203d2f1b56c05801a0fcb82b003de08c55faf1c7b33d320056244;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffd26adc114465a1b6cbcb4a893a46e33c62d96a5fb3277a7ed9a087c58f25de14de157b3e936a7eec46d55e90af2cddb98450f94cfbf13c735ad5f20a52168631349be34fd70f29e1818ae3e11b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31bbc78160853155a152c5e1771993d54546f3f1b662f66178985da7972cdcf3eb3e3ae15eacbd408c3db187d1560ba644fb83bc265397c66a39c6eb571f43b3ad5dd7bd08ed6fed20bf35af475a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1041fbedf708ff925709ab5a025beab0ffed2ffd38b420646cd45d05ba92dd10bdc3e584c26e8cda1ef9b6e8f72df89e1478000dfb4d6270cc97d46eeae029f68e10797567c1755d66d1a4df9dfe0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de61d00b8ab27a32f833bf0cf0559af084bb4abe4310439bc55193dce76924606738cb15e36438f59744a340360aed5f2b17b44c1ae2667fae33adad78d6d7d8c53cc2e675efb4433c1743537b5f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63594df88063d4d4100a6220b166489dd362a1c6c1a512ac9d2bf2ea4b89abe09c198e07057f4819fabf6354e55f9023e1abd757f5344d9bc592a73eb0c0bacf7fc3e956be402699d76be897593b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h180e3b77bc2126d4ef583f6703c8f9248092c2ecec9fce72456e058ca5079ae57d1505015ed0ed98445950657d4eb5c9effece4f2063b94256874ae88a0460db9398bbf14546c1e497c1d388f39ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9c28788e8d4a3365979dcc62fd0fdab5e3b08d4e8db73bb2eb7b61bb3dae4cdd663c41537896f9b73cf5f0389d92ee93a5e178df326c3238a809f0a2cf590937a00275f834c662e2647c21d453b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9cbe983807a6a6dadce8f7cc5239a13bbd9461d79ce37fbfdd4954765ff21d28c22e3a5ad545ff545d40432f3731403c11acbe53e2cacd1b3eeaec06566b801c1d09dd50cb0e95adc27b2551fc22;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142d8b000a61cf1e67890851ae194fe393b4c875c73fe2cbc2d8fb120eea374737773ae4dfdbbad660af4f17e84081927e1dbf02d740602c82275b65815186d5aa2d4552ccaae77e52dcf6af85631;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8f3bd9a24442d2455569dd2f719ebf59a7c6863498afaa5363bf960bfc5a8e2802eba2f14c9f08f867a03657fdb8f6823dbb99fb3c0d5849553d621c09582f90cfe2c022de24985b5b9c065dddb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16492335e509619f73daf743408d73b0ec097188c8a7ccc83fda50d6465cf3cad4872821ccfcf132d33de080602f81da8b760026b555c9f6f45d54aae99000beeb3e08da53fbb992c45a74c4c9f9f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1471073dbc7e716faa0022d5905ffd90b1daffb9addba5d1a5e23aa1cbc11f2057d21f98f55454768a9b13dd068bda71e2712e3d79fc035c8fb88d9bbe1198d30d4ae51919959152c2fcbf0cfa0a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144299f22c2e7d01ce11abc76787d3712c0d8090eb5773e5a7ecdb318fed6419624743aa5fdcce69944ec66db95309a2588f3dc9c6235edfdcfa418531aa104479800c7a486e8228264d543be6100;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd09cc395987c6f69d6fbc7ebe104f9978510280da313b49804a6359cd35888833eb4b64ec33deee8a022f69102d46ae41f01d3a9e18bd48ab0612515bd50ec9a3ef86932d12a5aa142ab31a72ffd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ebbb9ca76f7eb873b21428e91a2640c1f444c2920977f1cf7348870599fd24972403494712036ea7e7478834037686e5d4ad37f7638a12efc8fa6f685a073cd859f75ed73055282e34607fd0431;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h846daf0aa8e833c6af52c1308b720d52f7896717734a91c775e255956327995cbb3f68eda2ab456ac7b7789418593442da8fad4fd32ef8f10739e2dbdd586254e696dc2995a513e6f489a8da1394;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3fd415c9688c2d15814f034cd4f64a545f592b34e69655f533b8f9fb76bbccf0bd570e82d0e53d72f15b57d26ee65b6eb26b9f130989b7c70ad92f6152ceb6bfa383ba1711a9fcc0207bd3a6847;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b94f0bbac43f1fe07b0bedfa699aa9f510c8e5ff585e1bc839ccd3fa68fab9feb9c9124205f1f976699d0a4b3fa1a9b4fed1f08b0e1a6391f5339b95d5a165a9a074dd29decd52f88bb3cfa9cb3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb90b80446f178bf408fe2dfb715e02d7be9ce9dd3f34025cf7fd859e81a7f975bc91f3fd7a438ed78111df2af513194ffad39e4f2ba8a55759c5e0ae0f2fc6da399916f29cec384e587fb86ba3c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c3803ed2edc5c53611129f26e421af1a7fcacb1dd5baf8c6a9839563118fee8996fb32b7b800890e17aca0f39d1100692b403774dd43adefbc751c6855c8a00785ea91badc61ec4e056c7541aba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdadf3d2a205a4f99175845a2ea018497dab71e8095ad4e499774baecfd90661c39c5f1936b897ed4bfcdc9d6c696cd475122d9c91f08f8aaf5e0363235f3bdcb51573f427dbaa4a53c7fd112b21f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8927199a2df4d2439921c0ea017dc8eec6dc6406fee7f049382c46248ffdffe32f454bd18c77f985804a61231285f60a4a4d2f7c2d2ee3a0f81c6d97bebef6fcd56060936cd7f39e40f2bc50645;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce8a48effd8c75af84fbcc33883dad6ef0cd5de896861ee638ae05ee4b48b6625075bd00e70aee994904fee31a05e950415c99660ea5bc12d022dd33fd10541ff4b13300fd044767727a0d14b6d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b59b8a4f7eab4164136b826d424ad2d7a6e9b2d672d402693c22c741f4d56ac3b49089d5635128d8b750331f38f5ebe034ad1c2dd6c5adc29788e4f093c4c1866088dad4cb09f4ec06511d41809;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb57a8c0116471d5eafdd930967075a401246b3e67d1a715575bef433f72a7dc1c5ad9a260799b576b88d42602d0155683a089e8b3680556855e5e8a7407822d98da00997e08e3332bdd6fd5e858c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he964da4102ae2871ad9a67bf32d88a5d1a2a5ee65d4ae5d7ea2575cc4b06f323d4314eb6966890979a289fc45cbb2a5cf689263da28362b11171279dc9e65ce56ecfe8a563cba0d87bc43ce5db7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdde5f31d51dafaef961c5172b3a90c650cd98932dbed70bdbd912c7e85f69cc147f61fa4443021f2bedccac2fea026acd29703eb0f6c959bf4726347b12dd27928b501c77b172302532a218bb37f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fb606042aaf549e438c22c43456110b12b18537abfb2a2e661073065bb8c0c26fc6887d7aea42214483cec150817eed6547f84a3ec8be9916e4ffe6cf61fb5f57b0fa8936e01fc5c1552a1b8c66;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ab8f40745a57ddd1a7445b5c3069bc9d388e6ce12303a2c7e9f03e316b2b2d319e985b3e09a2393ab7a24c1360a25b6f67d7c522267cbff72fe6165402776e9e986a875e367e2f0f385e7d05aca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h122ef02b8a89724aef5e9c5907bdfa4712b20472bc4f2bf173e7aff807b9d95b752977497346494537e10a794fae2cc6e6a577ff6ad6d3bba4731c850e3a3be953b2e53dc26ae5c780eba1d3b3296;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h737d3bad42733240d9d3aa9ca1ee7f399a443181feee23c962f62ff398a11be66ec931b979abe10fc5f60b503e9c9adfb4c7e6323901f559ceefa446cecb23cc950c4bd0ac78886185acdcc27e02;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b19b674de04bb6313346f8247ca8c734a45da0bce52f48be48540e438c16cf22007383fa04028adc89d2a992f7d48fb63d966b39d9323a83b2788aa24124ac72ebdcfaaaec8ef60d80fb5ca2118;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf01e7c145f3f495e110b7e53b2acbf9ffa8f6bf40a583600243d49a7e56f1c1969775c453bb56b6d22a23ac8f1b000f383a482fc12be4914da3e518a125152d482c65f25f8a00a8d8060803662c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h252c03316b0e58e8cc37decafbaa41fb793d432547361b854ac80153461d1c08f16d5f4a1fa33d31f94042f7be533c6400f8834b72981cbfc1ff0baec1982455d3024c3c8e6f758aad9f509b13be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ed7c6cabe34971956d7afe6a1709239aea70f0ef04bce87586aa383c9e6c9ec2c5f0507fdb903a7d02f269a8ae40e5201ec93c8e9454af3889a4ecf02b8e60a0cff2ff3b08330189dd8faf7ba9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h671068b54c4e6a405ad8db5c7ce9cee2ea491984f53a6d06eaf273f0b64f0220cad737ea034ae6ae752c17b1228cfeab77c869c20c1fec0d9e56760ba2e199d4285550d37ca970e6248b92b92100;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb92f04e67d92afd9520979dcf2e73ef1f895e5f384fd7128b24e444850c0ad2990b813328a01498e9d61406cf988560ec0269033edfb1e3d89b7212692691683ff65cb02e1b2d10d634d7442aa40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f7dcb5760b37c3f451e4cfdb2cbd5c0d4ee11051efbe5b7b2c2a6346b1ce1043713628d95675a491a55c89ca266070699cb23469353cdbaec6188e612583e0ed3ee3684c8c725ac64b1cda6d9972;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc51cef2e9f001a706ac40b4bcc048c9564517be651ff96e36c90e98e7a11ab14262c15248f733303058875096465625e87e61a8d9a8624249d4265564f70918fa730a48e8d0d0db91318870e3448;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfc24897c6e30cd6ea9d05a59f731d42f68ae665b79b62a53f4f04d6b4b5ad798a25b8ab01ea92a98ec809fa1f097a3065a31a8babb248419aa738ae6eb19ad889d4514bba32f045e5b0b22357cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca0b9d8daefe174311f321d93f7459021fb72b4b8f980bc17e7d8634e427c5a3fdbb76cc7df99a22a91a748195969d88ff0f2ab025d30ba028c2c403215fa9c0c851a527914f83a4a4d8ea39ab34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24aa77bc1bd1bbca52e5e2755306f0aa6d787af92e10b99075525728685bd7e1cca5afb91844c56721cfcf70c5bf8f1ec294111a1d0a11f9ea2001899cbf3b7eedb746d385a610f24ef6f13866a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha350d14a720c4645a1a441cbeee8c1ab5499455f9b0c52527192f574122fc49460b09530177e1690788ec98689f5a490015488d75288799d447cc953c12a4e50bb1e999b9ef22e99ce7b23b5e808;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74c5940093321b108e75870f709a9deac47a89736d854d4e313773a84edaee0b1d16abe820d1b85df14aeacbbd2b884a5af1cfa57ac24647ff9ee34ebd2086d4b38e255a6e90c3cbf2d3ec3a188d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7e3e4289b6b7aea568ae0560e00dc7d68e9e421dc561d4b991a35eb16c57d4fb3f3591a7b8ec1ab93b87d1b4f11331929c5e7b9c6db2c5a778ce1237c52a2358c52b0cf61dc15cc14398d59d660;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfeb3450b669efb4ce1e1ae41c3f6fa6f7164f54c78badeed3e10b3ef7aaaa5602723db6814b7cd363e07ee53a5f9aa4446164ad6d2a7ffa83e4663684001c1e5ea579b0b521a48159323c6a2d34c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5572477939fad3dd8cff491597a39118269ab612e15d0ad05d3cea4475f4d5e268f9912189f85c8ef6a39255460f2f6d7899cea3449f1adc137e5f6c2ee919ceeaed2bead7ef10e5f5f4dacb381;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a928dc1cf88c53aca8c6666795514ab0e7cf92e7b0c8af6dd167c7de8d325a9539ad76de2c98ee88d3e700f1e6fb2e9794bce628e10cfe17e33c6540ba6e555d2b79b67e3dbef8197715b5cc1df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd4c9702d46e97190373412242da3cdd996c0e04b41d47e3b653156dff578b33ecc5fb41e0ca4c4277376aa6954d11c14d94f54bf46ed2019a742d169556f959ba8330a6a8b36340c0bb3a056708;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118e286c24d4ed596f1d057da13a303edd50b7680dbe0f0b2fd1c187058f237356fec94f41f60bc1a3deb54b2d2ef13ab92dbfc2ec1fe4d9aabd45559a3e8f079a699a4d429bf72db5d244b491b50;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa5245ea563f5be221514ad6c54f359a3e5586dd41271171013acf10fa1dd92ab558bc86d451a1bb0dcbedf3a0343a1709eb421785734d9801971d7aa935385c115187dcf277aec08fe7f9b4358a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ad173cf90bd04c3e7cb2f8e54a7d3cc8c0e4fb3daccdf63cd851eb5840c972d0bafbe22fef03d557007ce765659a067c49d44c9555999d60906fcae2eba29af3373f108582fcf8261d9ce29a4e8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1351c1a76e9191581ee141a411268cc42ec828ccc2863401b726b5bf51884522ac04f8c0d01bd0b98882865a8c505b572e4cccbe52bf6fc6e64ed8bc8abb24016763f7a98de6720d4b9916d64b61c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca404c68fff445d159f865a96660f4b76a54543a8870153ce06aac13d8ff031dcb9e931cd63e2bd505c48f84e430c2e2232fba3aeef8a3f05581bfaba78ba7bad7b011ecbed36743dbc00ac7c3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16827983cc2a2899c10c5be5089cb8cba0c26e2280894797b31b1e90bfc9d76fdafeb0ecbd15199d5bf41fd3a9461fdaa5484fe7a062529dc15f9894e81705fe69e1849ad1b67000ef32cdd8f1762;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h196479de0e07f260ff8422cc30da74148bcd0e76d458a85108ffbc73e64fd4be9c5bd0c46f1e55c58365d662c3b629a231df58044e90c2a271d213a76bf3099b62680f8bf6c8ddead6dde4d27a8e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13eaaa252eba2414688216eff1c6ebc76fdf11f583d613b0fab0ff4ca2447dbb068a31a5a2c85e74d72ee26a90d912f3f57dc84c480a8db529e2f91783a9ef4150bb9f425f27d4d2be6a6b3d2600a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ebda0d863f97c1a5fbab20d8f16fb50a8c0b2d63d692acd3c1ea42250685617beb9066b515d03a083d096c64b7fcd7f7aed1292a7b538e5864c17d296cd200d12982af17013168a22d52583087d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171f2634bd6286621060ff1f671c25307f2c6c7fa618d095dfe054c9dedf3a09fc63ccce71676bbce1d135b638c0477a56912048108dd5a6a4960d2eb1544b35826f2d1cba8bbe63e95d694d5d5c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2ecca3705e6a137734c4645b76e4ded5c975de8ee46feec857fb8d65a130d8e3b50ba87f31ff29021c2e41f727c102d697ea94bdf7f2345eeb1882202faaa2470b8f1911c5a28640597bfbb2314;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h102f79e3b92e84bae67278bda64e6c3285bfa75085db5b455524a034a6f7c1391ef6596ad8b42c75eaa01f652013ffac2b83c69673d9c77a3893e0b61f4cf9e7c6b2de1516788cb659523ec8379c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10bae03f24c641525b9c7e9ce25aa9df4f3ab6ed1ba9e3b5a6bd89a595367ba1f71f3bdd36290779135cc8c5bff7aa8ee7fdddd37a87f00f52c71feecc7233d31d79b8215782a6e9b978147901613;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c4665b533b476497bc35e9187dbbe5b6d20348d1c2427bfb5ee6034cfabaabb1e449c468aec295eeb3b456787e6da9a2d264327d501fa58fa089df9fb9e815c220ed07217124635ac9cc28bcb83;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3ae83f4ed0442c1a099c037fddc8d3830d1b37c27d911bf0b43a4dea8e3a47727193fd6c86205165e2f1a83cbd7c4a9d7016eeecea26099e84493c003b323e1411aca280f4eccd693921731d0973;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1486f2a0e38a0a058c59ac51d70c45ca2990f518250acc773ccba4be85717371cc75014078bb35f56e915906f571711740a6eb50dc710615550a6a68a09d9c987257638553e41bb9a79c58a3ddd56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h665ad045eb2878ac3031137458dce07d530723e47b20a8d3d247c66db79303dba2258786da3cb0fae5c9335b0d12a9dce10cbfb08bd970e8df9d103332b50c16a5135db6871a947e4f45eb25c355;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a6fef6e1ca98ab7eac6163c8981e190c3b3aaa2ba82a12f0ef5a62334b4e06c90e667cefbbf4bff74e53ada68378340008285ccc82ddc2520a7e8bea5673a0c9974e2291eda413f2d6d6b4d3e0d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194ee3d91ce2380c36f205797cf829e7d152d1239075e9eacb66984cb8216f048e6589e846a1153f1acd29f83164a2e84495c2e5d9bf1152ea5eda01cac567a6da987ef902b509f145d6964677a95;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb5852a83a566bdc64928d22d7e6a84411cabcf2f2b06180e44744abd6a77ee0b659173cade6a004b9650645f768a9194c0b41cbc6c16111a7d99e32b49a4afb08ca131336342388a212108817f4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1033427fd9a63420b4d3106568a0187ec850f8c49fc459d5d2edacc903c2ab520f2156b02e68ce63e164c36a8ef7b940f14e21130bd5e86be88d8f51e3795aec5f636cbd5cdb44bb8ef009e22b4c2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b650d0ea3280964be07e838e6fc1d86b8807c616053ba43fac7d7d3b57083390a40c9f811742e43b9f3c24ea9e4912f969168af2e2c8b08611c9301846cc33f913c7df10a36e57d94bcd99889b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b073a08af159a01ef3a6e2d442bc364e0e3819cb9c5bdda184058da918fb9d8f711f8b014e992c44d3e2cf0693b25da91b1156bdec3f7100ce2cfe8e21e933a3bfa825c02733eccb8b60edb3beec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14a20975511be0cb9f4da55f785379bdc3d0235575409d72b0fec73ff2b7ecefb6fb176ff916511e42d56d7be74220dc8871edea329f0e859eff9d137220232664cc1e74f0539f43934917483a1c4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1227b26005107e0d5680a8faf55f226dbceb3f840658e8d7797c3abeb0bc6f27a8498645be27db84b6ebb5016d5a7dd386d9307e2d388962c12364ec61ec449fcfb7867fc8a9d5f98bf35de52851e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1adeaf738bd7fe77d5f3f2466da46cbf90ea52f2ed3a5ccd9544852aa0725ecc7eef067568b4efbbd3e07c3ae0ecdf6c6e1ef25122d53561cea81dfe0b66bc4fb941531429bb379f064ab8500a24c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114a34cdcb91b28d0af2e45631aea769df3537eee1f8b3746b44ede6f8053170428a203b6711cb84511f058d57edc370242f12d77f6a9a3d6986a2c13fd3fdd7901aaf47e4550073d48b8185a1f81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha5edfc92b7f57c4860ed5baca705f94919d1f58ce63faecd94cbef7bb09f3d5ea8bd87e5c9dc9a8e2b9fe788c5eac09850aaadb1fc5630b916c3ef38cf790e7a8d651aa759283b3996226cd591b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4ad40138b2b033bb508c6ddddd8dedb7eb6226cf24756c94a99d33ecd0797f04379ddc87feec59ae8693434fef332162f00721c6e158dcee1f62d26b8b76140a2d20320de7c5d5bcedc272963694;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193c0c879ec74eb0c335f4fa1dc9630041842ef3e7ee99e02e606cb6c95f439badbaed9cc79006428e7064f89dd0db1158807cfd1cc36bbcb21314433d5cba59862be28fc8874b0ce6a934da88492;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h185ddb94bbf89d634b515665da50c23a5d703d0d3e4a0a8b25cb7dd94815d9e1946a8f272bc26b9ca00b7186fc14c95d18340f91906165d8b19830bbfc550948740ac6a1ef60f20abbaf6408daea5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1922cd6fd1404031d7272e14ed9cdb0ffc71819019eb80600c99ab6e99ee22fc1f5365f2f71b2e9b77d0913612552b81b6903a3fc0a23d12297ac8ec8ad8e575ad45d5b7ec7964d4676441ee458;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c55eb42fa76d131717947a813f6cfa6bca504199590065092d2e332fae1875697c1dba5e40a711b04c2096cb1f6eb8e28a6b3f62c170fcd29793f2b2f773e7903d9ecfac880935cde6a3202bafc4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a7eeeb21f4d79fdb741d4815c28b14b26766d636d1b23ade7eaa1190da4d71e6375a3767339d5ee1607d7805c54574329963ca491a597be7fd02a71bbd04bf1c988985a1f82440a8b422dff6e15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b5d98bdfa6c9498e1dd9137c00ab11ebd27a889a30436c3fdd7dd95553c43dcd4030f8cad5d777b965286da079b6bab0a2cfc143e34c1a8ecc9190decd97532de82abcfc8e676db13632bf857e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133a7893d3653134a8ed238884cccd6e7a5ba14febad97d935c1c4704064ec125e1abd4235e4683fda9700a4fa4e801cdb7c05ce3f18323b27041d2f68d6bca1d5e5557ef87b54577c9d42a3052a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc9fc7315eb7fe1bc41a1f04588ec862d418f4eb58b6ecc70c12bdbe97d9fe4850eeafed0a877a77e4666729209eb9634bd2804ed249001ccb7511ab838546a4b4178a52ca222bb0f006e1c89dd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df61b439d015da96688820c635c215a633742eb819c36ce457fdb0aef4352a5278fb431aae414efc3095d07caff96c31762e571d1e9315f301f51a1503178e3706658516bd9d50216c704ad5814e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbf2463242d5ad70b454fd9a937c5c451e6c373579c60e31537b543b6d6872c8265376183fccd61e32fd986851dfe0dc795f047c5f70c8b78d18f9f13056e875169e1f02b8288da53ca51bcaf451;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c890877e0c514a14d4d9eb8a3b1aa6a025b74b5e46e28bbe2bdf105da1a875459c0cc139ad164323c12d57235e30f1453fc7d7a963288c99bbf2cda8461acde72049805e66d0511c47a145d7e00;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80339cec1f67848ba65ab193dc1fda1fcf7416e43aaa66371a959b50b762ac62df57a40b280e7816948f16a9538424f26c748e8d047e7fb86fc65efeda586bb6c67953b7426751d4d65441470266;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h183dd2f7e58d6de7d2c11959aaca8b387e521473fa40703974f03ecd475e9f5b0ebf68b94c1ba92e85859186a3cf253ef2a4cbf6a4e170203640f6732d5066c8598faa3c0f442e600e21c7d438380;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1588ad66745041e552e266e55efa47d90c28bb3fe9008aaf720e6fddb71ef2be471543ad2d72ffee9f087d05adc5df4f32bd9afad0c9831e3ecfd458521b51202526c16f0f71863ea2a0cd41676a8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3835d792808c78b3aa029dabf1f0222c0894c7a8a0bd425b05dd46db068bcd701c2b7e2e90b34b6427b286cfe574b8a6732b068997381df44d96194fb0fa58094c75cce340e2e2de31501939a63;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182101bfe37bc0a7cac864a3f4e2c970b0193882c1c22a837fae153a617ddc63cbd3a1308af108c2203b7d4cfa8664f69a4f676dfc5b043a3eec46acbf71e3d40d1ca338eea6acdde358599664dc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c42c1f0dd28a305e454e8341f3a001a74dfb6e1e95467c43cf4f1c0f1379a8f90fea359fe345f13fd98f3ba2c605b1022d40d8050961b2504976d39446ab22fab54ed3cfc24e66146448d96aa447;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h762cc77cfa104fdff35f5a66e6040193e4473c6d7f62c3484e61b3149d256aef2b82c5a60f6b5813c1cebb971e7d7745a3a51feb782ac286dcece1f942a085035602fdcc5efcd53103077675356d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8dd63e9f03ada5c761077e4527c14bf8f98e59549fdc2f43e48fc89b3a1f72b989b7f9ee87f57378ed062bc9bbbefff732473bdbedb43d30151c2b554436fbda5301decaa2062c15cddd118469f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6da009f3e8dc70318b609930bd81afa9539bc0f8b2819341a8855ec853c6dbbabae2133b2316413d593647e86ad2c5efc46a1f32e1fe594b58e17918a928aa6df79881496958461881d88ed1553;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h296a170de1c6f6cfa9621cd68e128db74468d994492279da4931416e8064aa47b466ea658c7f7051230b360d21532b8e6fd502f2903e923a016dda0e2d60df7e890b10aff68dba8f184af8bf1596;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1445966c2ee0f0aa350d2d5156db8ce31e4ffe007fc74bc2289c0930e5db1476278d66a68c3d55fb98b0cf9fa0c574c900c666e30d539f273c316cf45a036592aa0f8ca802863968a0d63ef9db5b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba5218de3332271d0ab59d7d92728287f4298973b37ae372c5baea8c566d4d9c9e5571f2170ae695292c7eed6d573afd38ae384e7e53ef642c765fd983e4278bbb0cc7bcdcb05607a3466d6e881f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1385cebeecdaea61b461c3fe85c63b475479cdec89acea650cb3477bd3e356b4bc30d22c65a622242db6a06b8220d3d731201be8ecf4c3f61d190f090069d8d2cd2be9ff4aeceb43e672551d5e9b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hded7907ae90b63a405f1766a05e6ea41b87a424754a97850101a94e5c5dc404f8da071c7e3d11ef5dbd445e18ceaaa5144abfc178ff524b6e8442b6fb5bd4b69967ee0d69a9dbfe4113c7f17533b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18612daec6510307bd39a4848a279b8f146d6c003f52b15271b0cec4a906ae594050707a15e7e4f438b7943f7a5e76fca23b90619b0b85b40c762397cde4a39f5d318eda9817d6c8d1aec624c8dcc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11f57bcf9b84e047aecda13a82071fd9f7e24ea76ee57c48f5604e86337e84bfd74c2a4528c13c180e90b55decf4cc361821f8729a0cf9267163eaad01a6a085d07dde5033a1039ed1ab9ae35515f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1c3bca089d520d599a37a4b75b9c256d4358dd4adad0de08274039575f834ec99040768b60aef6a2c0ede3ac532e9646cdb98126daa5cc7f7718ca2b853d69f8a583637b7332fb3b0e856caf3cf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19da711625f9f83e17fbaf4d53389d1491726b8b6d98b232a8563c03530ba2f6b6596b97bf8d67102ad3371afe2234804166971035b1e38f49c915ecd224106550e64724df94ff3e52e667f2243b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1040f231da9b854932dc99a5a246528e473210f8a6ac39986571d262336f93c9e4f2faae578ee5a76bfd8410b5bb60412295b0d93a01a15d15e7dba7f54b3b5e8e1c9a6136c9a166fbff1edb74ff7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d546b41c1002a522ad8a786afa688c9b0b71c0078b1dea6b7f37c8e463298fa2ac0c41b68862d531d845672900de116d5031f6b92d6179ad00dd4475512ad9336e5e39243709a3494fd601ae281b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152dc3ee57cc720d5826abaa3a65732fc290f9724297cce2a8ef83053ec96dc77bc212d12ef479cfeeb04fb7caa839f8dbed3889c559956201090fbf0811b9dff7fa3f2eab31f7eca3a6b42cafd96;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h49744ca6a9e13e24e2e4e8e5aa574eab7998c3193bc6ff9bd22b5f7b89497d13c3a46e5125a967f3482f129de57c60f9c6187568517c1c59034b3338479c943886cf2ca42e04654ec5ae0236d702;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8bdc3aad1a58ad33b64fef5ede5b5c7fa9678b40348e996b04db516a8c010a73dc51fe10fea85545d458b7fa9cf016ed9157681b96da955e3a96fb8bf7a24de8977e34c15368c2cc78c3fab50e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a074c1efa80f3103b22a1029aa25f62c26c251b4e0fed64fb6f1bf8226189c4fd25a27d559824ea6def847384ad274e3a75f6752db90590267d99b0a8e1f7efdf8496449fbaf1a7a388806e75ab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed650910316d21e96d79fc7b9264cd5d34394f9ca5ebf141be470a25441f94383181d7eabe96e3086556d592ac515ec629b4827a0ef8af278323c96902bf11bc064b0bb75d571fee0053825d4058;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b36b16c78245e88db40501a81115592fe1502124fe717f7f8c025762347d767ebe30069620f31dc575b35e9700fb1cbfc595557e0c6d2d361a9ff4eb8c3a7be8d92e9fe8bb2b0e0454410dfc6790;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b95d09740634d51c3ce7ef73f893c0552444ea60272e73f9e2f4aff5e0963d45a07ab3c3b0d04908cb649bc1e8dc969410eb634538100843486c1c6c6bdcacc39368d578cc0078e97f82869365d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d6797b32a099bd1ef5278cc7ca3026008017af305c48d415bf1bfe7921f578ea250ad9f10d6d61df97dee950f793cd73ad94a190f3ee7aa3fa7d413c8aabc393ee69133f30ad6701b370d547a30b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1004aed76dd335d2b55f34d4e7a928adca113f9206f15bab4d71d57abe8dc010e6d0430daade18fce05bc804ddb79de421d7f5ff31cc771481ca6a2bc9928f70109a47b90dfaf3fa7202180df6bb8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbddef490fd7d28ba237330a84fcc7656bfc35d79fba8f34b74cda0f28721f4e733c2f5856056f1647b1b9ce32f8747795faec6b0d2fd55de9a2adc8168b074b105107f7ff57892e6b7110639db60;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h71ebd23095034ea1937a2a200e4ce4af903a91b4a347747adb98c5ca8ce5725575614d0d3fc0d02902074e64eb151ea4a333c102c4694d0d07d48642deaac17dd914ec1b89d0d4e509b215a61866;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190f986f3dbafefe045b29dc5ebd1da14286754a80468f3c1ef890e15d643d763cf9ca24016e8b58124ae91e877e3d66f1c3e61efbb44ed9484b5f4f0327a90898c2f4dc0e0dfdc2b74368425aed0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c515ede7bb92790abbf07b0b966bbffa889af2dab48eca36da87184fc556621478e26256f0b105d881041dd13c416a56d85dc2842c02caca60ee79032a8796dcbd215db2ca3c44b553496856d243;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1461df433bf1dd3f07341ffca3c019097136516ef9ff4cb64d71abf630d56afcb7f193bea1ebf81940425a8d0f2e71705c92a1d813834ee11d80d92645f6dc56f494b23a88e0641f34f9952081e29;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f5aa3f0638b1a504e26b6e560706a4cf87332bdbaf7babdcf450fcde30aec428c9b0e0e9f242c81e6c503137abb3549f22cbfbe0c4216374351292824b42bb9537b36aad9e0ed5afe5b9f34f053;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10074fc3d3ed403658541c5be4650ed7ce011480842f7fb14094eebd1ddebe8c04a8329a4852b3208980b6e2ceff4ea9d9ad3cfb6cffe5f7d68bcbfc93c25fe6a80bfca6ec2c6afe82fb0a05b913;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18290f77d92cf46b6015d0b7f7b422712b8ba3f3b7f4ca598a7f0c76c2842768d5ef008c87df2194a7552fa470fe2e1466f6407c2d57c6d7964d95c0972703580b9d0a99766103044257a7ac1b77f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c021a0cf07845c263a24b15a8647632eb2b54eb5e629e06a00f6e69953b7f73712084517a57c6e9ff28bdbf0f17cea546c185b4993e9eb3678f9d38cd8d11141302d2d469abb5d08baad40b0eef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b2fe00034b71a47fe7ce619cb1b31abfdd4595d02ef95245efd3f5074e8d011a4eee5db47736255ea56138cf1e9360b61b4182246f8002f548700d00d40ba07c826a10e6aae05802b2a1eb779e8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5175846431b87d5768e3ea43410fbdc88f82b92ec687cafafb60106aa6e509b61be39f96d83b347e2ec06c044a4766eaeee0461dd3ad7c62d041304dda22eed288d21b0af54c031be59a220fef7f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf6070de0f0a41b5007f9f1bb5490884a4ca0313ebc8277211d148a1f95763ff7122dc37c77900428aad058317d56534706d6c53d0229b467cb4651c3c8a5eee8c1bff9438221ebc1fa5501dc7c32;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h842369abd2438e0d3adbf29592293ce57f1b94661dc8fa5519fdee83bec30783d43d59cf9c02b269859f3c34cb6ad354bccb99c79b29643f92904f01d54e7ef9bb8e5bd868ea8f2658881f6bebee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17a110dee65785c385883f2619527d532518b0906f65f2f6a082dc94d20c3acbd15208708684c87b09370b195762a4aa18e438dd6e4d8e9f6393dab710951f19babfbd9cb57cfe6c358f506dff1f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d1b69067b00afb337fd61e213596e556924bb70b4eb5733e293d34c122f2971c74414fa26fce833048b7e9f4650ea2e4aab7cbfe27b7b5ff0e7b1353b1182331d13a6557d214d05b3f63fa457fd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8035f7aa6c0dbe63197be799fb534b873c4622b701bd7cd20886ba578836594cd57692a34eeec428d41e8fb8f7326617813e691d4dd8fa12f1d17b971979ab87bae9a5f871f34ba09045d2441c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccafdb0d9fbd58b6774905d18c327ce6a929b6a8d2b23532b5fb8566f543ef12268832de2a6e7abdd1f64a202f70a280f02fed8dbb518603051b5b721e2c90f8eea90455a9e1e1a300c9fb2032e0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa5b67fce4f062cd1a650535b890d08196156510d6391bf86bc43101a5382c5568aed7339d4bfe607d9039b74856377cf8e88600787f73d72a05b131ca85862fad726ebeeeb80d18d9e14d83b3c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h370fd143813529f22e5a74908ae55ed04a0a0f457ea324e79a6d328b9c162c59859b56aca013d7fb7643f3950581cd17e04b0099331428687eeff56a011cf88d0a2c59bdc82b74806f0a53eb71dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19fe74d5d8d6cdd8cd718929e5947d679be4a3638b147c59077d7dd0daf407545917a51802315fab2b45b0b3da04594c15f3f4b68e1e94be879f630e0b321590568155f08617272f09a6d95d12aff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1790a5e6491720236fd2cd3f096c12ab7d9472f9f87bc6c110a28d065ac6ae911e6b16ce4279892b0cf27d5744c718b2c468604dd43e5abb84c9bb32297221c163bff668650f7aa5e6a86a0d1da4d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ceb9c2a57b06c29b2d9937dad912d966563ee93b5cafdbee860514a0f956a387cabcad2a3c1ccb73c521c679df724ce51725005e518b4a1f622b695a32c7ce94fca5308039fa0dcde1a2c34a9ded;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf68b34dfab03376961ce22120e2051265e743d394cf1b919382c9c1b954e274e97f5e17b2c06dff4f8d53559c5ee5ff694bde3e9ff8c0037c2d2eaf391b363273dd0512dfd8c4b7ee960899cd1e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121daee5ffbe6920576fa2484e8ad6479d579ca2f118f3515671893f5d54d40902bc68535bf293e7d3e06916892a3fd4fdc098c9b29742f3e1d6f3c1ae3411d1a2ba7ad5aa29c6d830a60a8238c4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6528ad5fef8dd69280151d1456d990785384f76ccf55cd5cbdfd71ad24a238a97da9d260bd0b4850267afffb33421d3ded6ca71e4b3aaaea52a2355704848def02d3f64fd13f0fa0cb7320e9b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha82b3cef1b55c22b160db8fce22717f5ccceccd0853415eb4aaf40082c029b982728e34db0e9eb2953ca682dc0a07ff63ba813cfa66cf163925ce6228a79ddef77350104658bde1780fd6bbeeab5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f087b005d4d2902742b4de6652e2308b20c23cd16bb4f7c6e000bc6425921c6059132bdb8c0df733cf7d1bd4a3b94f668de142233e38e113640ad3b8ddbc2accc14fde51a66612e61d55524eb139;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5feb11f40114f4096fa855bab21f16ef03a088562b34ae05f220c3fffb0aba52aa0a48fe79c05154e97ea25151663b65f174f177f240e512c22fd90e21e9df70c83cd8a556e488f6ba293f73c4f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f70cfc72b9f03d7706d9704334aa996cf12a7bbd9f9bf2b670a9ef9d569213153e2163651b5ab16dd8781c5ef28f2a04ae376bf932ae2a089e8fd3317196cb684e0343cc3f083d9b9b077974c55;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8811271691e4ed1b78fe6928ed286cb4f38bc919e749e1ff51ca92db3e9b8e5310d582882595e108f81ff5e6c6941fd11c1b6689c7cfe92117f804f54c3877f5672ab1444a37e5160e66adf1958;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1994d3fbd42867d61267d0f86c2f91ad75494e2fe2cf401e8930f2ef73bf079f6eed897445669e476a713acbaa4062900e6c998e629de0b93dc584ea583ac9cf370ec1561e1eaf3eb4de2f4e7918f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15260ec97374d20eff09a64f5a7418979ec33d059ec189b4f519fb902fb4e28f1871383bdbaea3e161202375e436a69867d46da4839c7b26a12a8cff5edcb1b54a1bb769131b258ad8440dda2a491;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c557ebb5915d6748298bd345e7a0eb4de06207aec7c5e1c2f3a598a1f69b4e41a5cbdb2db287cfd97a679b4730bd2e06fea36b87efe767fdda087d7ed2d02ff40df93af160a75b08465a986a3a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1f93d735ab0923439be645ed9db73e614975fdd9a43a0c6028e60e6a8c256b899da965c44b067735add38bdff9aab98601cb45c7ae8700998979d7c200a7205be78457868413022ec087b9a6571;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h23c57a67c6bd6be2267ea7b0d589421b09d898c2b8a4e75e6072121dc3f92315dae9d394f4f2971d6083bdc46413bb9a1a86a0f6a6f63daeb5b534f787b3daec91e85a6b66b1cdeb0169324d45b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191f8c120e8bc67124303932750eedb170678f1d612c1fd363b890f187970862750878180ae7bf17a78c28ec30154b2719fdc55cc8b3832c011035469ec4b0d16c446f4ab78e3a70af21bcb1b08e7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a596db75bfff39d4781f8f59f2308c1940ab11dac3ce5fb5459edc4d201f23196cedd305eb6b831c9bb884c7ac3085a92d2662f610a057aa8f223dd04e4084884f3a1c45e3baad5d65fcc3991422;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee406f86deb7e5499d90ab6fa260051dafc22849455d30b9967dc39a92e1d9a8b720a59b40f7094398a86206ef1bcc94c6e7864af5289b6653a400cd499ffd3f3b719f1930d784111e99d45030a6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163b9db960873c99f6d1391dfc9119f04fc51ab1160b18ee00ec3dacc857b8e77f47a881f3020e52d46646489c43414859cedbd77f738ff3488818d8aeba2853871246a0a9c4aace9179a4c2254c1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1455cc28e2f30374b047560ad05cd3d1f68a2aac044049d22b382201ce514120a68c9244c257f8035f62b33856ea63b44ebb3287de320155f2dc7ef4457544a3f11f4ee517c9c98ccfb0f5f8ecc01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd95eb8691ef50a2076c4d8475fd917cada045517d2ccaffea7cedab2c6a7797cf625eba04b8722385de7869e81f5fd56e69b49e647430d2126ce4e5c3ebb0988fb2e8854e67c126d7263dad789d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187d457f1666457afad68a4fc75058d2aff246e8bd1959a21551f285ff07f6060e6c5196ab04bf0b2efce666e58a31ec2b0c16e0d91b0df3a5bcb5f6a87ced8746f26846f23ff6b543ff95f72863d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1427923514b3cbfa963d0a85f1dc622a299ba90ff8a73cf407f25865ce63ae5b4122bdb7cd28ebba7f3edee950b5e4fa3d9024317ef93fbe31ebaea3c3d2c3cad8b35d79bf8da0d8c4530325c0fd7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f8e2aa36a7bae0944387327bd9155d09d45b79c6373b3fd6585113ff93e2a34a426e211279c28b8585ecff78a17036220d41776bc304522f0d82c77a105c86fa4320b61f1f64ccb73e36b2e6b2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b6bc8a3ee72a344cf09fe0957d0719720b644be40c3208a1405af777f69c9164b3591590702a4ac3ffc2103e1df91cd24793cbe76fae5706ce3ca0015193e4ab9cf0235e853507acbc4698fa012;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93d778fbfbbfd18e789babe04020a697860a4efe1b40dbf899886e9bc2b39196a579e3c9f4427492a1cbd88e95a05ad58041cbcd89dcfbb9917d8c7bbb8f2297d00642ae061a0e5d35912a3c3b93;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1b870af8928efb4f466bf25e8b991f3a3aba68100054e202f253902342c59cf51a8b8e3ae7a8131cae047860d472c2b7d0d14ddd5b2de40fbf14c8d5923ce82697838a121e7ef3769f3b6b93dd3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135f610bfd65b069d57aee7a42521cc7f4f8956651829807ea056a8a3501dc45ea5fec43645a45359b678b35a7195c76b1a588e172ce76d6d074c79e921affcb3b905bb22eed65c410150af6c056f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1a8dc3c929b0e46f10ebb11435b60878accdbf66cef5293410b965d5e4d206f881df9fa274d21c55cfc88305144caa3a1d311c29d8b2dc10e5a23186040390a2c2f6b14e06ca21d7ae5058df854;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d71090a8fcdced73244c80897e8815ba69fb085ca7508901a659fdc38f9f4e5da270b53a865d8d5a6eed3e69c1213cee7101b7d420c2facf6eef27e59e2196ace0bb0fe360b1fc17c174f0891ac7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ee2caa2b7b8bab9a4ca9e981da73c9eb5845544513fd97c8b37d2edb645bebb81d9607cd88142b20ff9a15b31965caf180d70d23e22aee258184e79bd9f0756c15ddc7b7407c2fe5c54fabf65b48;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff108988d45d29ed366bf4acf369aac5f04ab1bb60c8e95d26d72e7a6f04685dd0fb923ac39c05a603f92c1cec95d8105e8c5b1076e859c8f8f2e059473e91a1c7303b1d594de832c96e5dce314f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4d15d444ff789ae39c5b2feefc0bac17483c76db442b1de14eab581014c7beb45646a75b2939da690a888c535fbf5406fe70f8c1dd802b3d39d263863daeff71f072d90104dba5a46183c69092f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e2922c3916d6fc8aeeaec1b59206525a0b98b74e9120e694974a61eb8aba723c33fde7b44e82bbd341783f422f8f789a1e9f7e9f67c95f60ebfd4c4f7b7557d75536053ebfcbba3c2c94c62b97d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0f3e1605f4cfbe8cd4cecd9a401f4c2a35fae5c2e477e0e60caa175d80179c21bb0ff946dd6a59f80042883b6c3ab8b1915b12f0e9683b0c819c625684729f878ef1ea699628ab3ca95f48b9170;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1253053463dafb74e489309fd84bae28094c682d64816a3d4515ef51d096f9106a2ef1390e126c487564d673843df9d16be25dbd6637da4fa4845fa2221b1b7a8a618b854c568940d619359c28ac9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc850d192a04ff2eb6bb422c432f360de23d68b08f8ec1cdabfa07d0928f60d4f3e6fea2e13d70f28b796ed713413b057c51f29a605938c3e20b6299f9be1b4b0331750d0488ecbae3f65edf5562c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2735230de88909de281450f65e7e999db7e2b131f69af72548953eae321be5389df18e93e30c7f0fdd06ef9bd35a35db23557ba4c28d1eaa8528f461a574dd01efd97c067f5d6162235f774754db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1948081b0ba3b09597c4fd39940906cdd3706a1439fff6e95398958de5ea4495ae93be6f12f2fd2ebd4572c26f7547b02b5c0bd031b05ec493dda50fa86a64b17cf9090034a87236f99b124d71c7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e2740a5e5500f1a1524067319537c565d94c9946e58c67164196974c8c29c71edf2ec2ecc9b4867b45d529f4371b3c1742219be41ab79515c701c1e4b29c58130252bdcef29258b68b0f57ef3ddd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1850e160afbcfede8001843f0d22f24afe5c562ed467259acb3e225e63311c1412999096404784415c45d28b11feb964b531cb4ba69f6b4a3f95377faa6d099d2dc629a4ff8396c6c312f59a86ecf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111039b5050b642b6204ed1b38a0b2d938de1de31db08b5db3d9d9823b74ffe10bf0316cfedf2f0d2019035a346a62c46ae48e24229d1a3bd0689d7be1f6576eec6f03cdf33489af67efe76550807;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62e25a9c24ebf53c4f317e64650f9d9aa8d0f07a092a24a9f60e490aa76400a7637fd9dc6fb0bb1246022ee5251bb9e2588a9eb15b1013283276a601cee8f7205300635466327772a03b7bbbbc04;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h458257c6906efa80f2db8bc95efe7eb12af3b0c5b02ab4668d3d6f362ee8ed96f426606c727bfa1b3a03eb12e3ef8f0aee22662a7ea6b5a9de4eac98a5dafc20157c7ced47b0acccad88420e5520;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1979db6ddbf510be55ff03df30c432e9f2bc58e0c3899009a53460b957cfc6c5196a5171dc3c75997c927a9d9fa0e82fc55a0201cfbde8279abae8ffbb3d775c8c39673fbaae637614e0d24b486f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30422eb5c6bc76d44f8284e08352127da1e77e96f540cde7bf0bc65131dbdff5b333c6ee0b05c8bea661a2d78cb0996dc642271149385c6d15ded0ca10c2532976ca6cba300ca3f627cf5e9379a5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ec48a93b04f44e2c72cf1192f89e0340062ee58445b6f5050613cd8c98ba7d40c9dd70a4f4e51c553807a03216ea1857d1f7ba458d458297e64c65f2045db4643e1fd7dc0ff0533f0410d48c417;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115e6d38f828ced4288ca874291baafd183b391ff00f0718b3436f9f2b685d0944f9cca6505cae639e046410626f807543874f27746456f87822895ee503a5092656d728e1f6b1744b373ea515fb8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h39978249a8b12990f62390590c5ccb3bb25f84fee39c7776e392accf28fcbc1c8e474cea6c11d517c72e73e8a0ef296836649004265feb38230183e56c1dbffbd743389f652c397076505dfa7613;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2046876fff4e447d95ca0836228f06c4b2a07744df96edbd2535a033a4658d51bc1b247f9750170de4c6755128e800b321cf60997a6f5635a9a09498bde82eb076980283547e106745e22564266;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1512058de947d0703b4ad810de1bb249a03d2fa55d12c72ac3aab0b487b79f0a96d2f6d8d4ed2cc3c11ac47fb1dde28c8cd43db86e30e08fe70ed3aaaf11bb6c915eacf9552d3205f872d58240397;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd99c72f2444e647f1e0982d564bfb4c1fecb84b55f24be9223c991f672b317716e1eda8274263f5cd391458768152a919da9e86495e2192cb3f4bdc7d0cf0c0237fed2893efaf9603418a74d5d19;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101acc27b24368d925369df7a7600f9972855bfcdc7ed7bf43ee56dfcbec9565a2bb9fa2e8f0b100179e3ee583e5041b8180e4a959e81f5fecc5ed12aa722236d14f9785024b8cbcfa8fedaa1eff0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d88ef680be14de0cb1f1f2b269d27f30348d0b67e2a8fa278084ff97a6ce54f852c4de8fc8aacc9341d886e7539bad2e45bed6fdeb2d3efbaf45565846f4f91cf55b79de7b9bbe40a05757f6c2fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eec9bcfdbce1c3a4baa7937594dd83ce1115b971fd0896f9a213ee3df8630409e7a38b64ebd8b31d6b44f968acb3c573afc53736cdbfa423064e282013827b6adb247ca3e768af8d7df6a76cd183;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd0578b2a2beb33a21b8f17b10fe337e5e80d12dcbd24c1f47cb75e983c394565d96b727bb322de6d3263bd04968ea604c6a5c12e065fce1d316106ab13debd1c8314990c995bc92ea29b0a268958;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had161c0520783cd16c1298d9cb41337fb6252895e25624de72094a0788f40a27cbf2bb9b2d9aec80f489c62c830a2e022e484356530b04c141229fd1c9d715a49868bdd847fad712d25bdc6f35a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1702737e35c1ca909574084517109a51af6a960b09840d840b4db32883a1ffcacc4c0e605138f9c0557cf5d8dadb1ef1635719df73ae90d3ea286398476e0c7c620003e72c01f238b19de9803b85e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he945fc9bce7bc264296c84f01f4035297ed7d4a3247e9d29205e3b0252232d570da06b4f86964adb6a7b5456c2576075315909a5099f2293c1df429e4b02ca2badf108cbe4644661fea8028e007c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h508756012825bf3d14095cfe23b3366ca194c868a3841674caaaf59e564efc2587fe667ca02864e15d4d4849c7c426bd7df67e5bfac95a05b4b8f9b547af530eecf8c7e054e775722f34fe0b01b5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h145e66c7cabc13fcb5ef5487588effd8fe819e361190f496a1699f1a3f3ad3517552b83ac61af44b59b7635a3e83542298be899e04d28c0df6d4309013831c18e27d31e5f8bd6a8a5e9edc3a53e7a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h282d7e1ac937fb0b7f0d41858371cf12d751218462662d53ce8da3753bb987c3a87a9b816c0bb05a7e19387803709ce40c32b3f7e6997baf27a4ac2f01d6c5bf91430f5ce7f4b93cf182ffab7999;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h616ca82e78cb70d7b0a38dfd8b2779d47a88831842655d8e344894127502a500a00caec7bd576b0c1384f2019374b215cd5a5515a6177ee94a0cab106b09adcc13e847e7733018ebca74fd9dad75;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b8cc7e1d298969dd98b4e366711d58e635353d8961f625695dc94f05cf01d8e7df6f210c5302aefa8db3a5fafea4a8d7373b93385161f1623dd10cf20c0cf84446b63ddeba094a365e6f2faf1fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d3b3e7b33e7416654d76f30fa8d94a19945fe49677f2f4420283370c4ff2ec53a73017217183926342185fbbd79fb6379fbfcaa00b8576d020d5d30185b2b27cc973bc7245a67e3ce38f2dc51f6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h962cb1dfacfa66481bb916bf52dab3978d2614776dcfada928ad257bb2f64fcae420ed46dc92c6f26794e2e10739b057f4f32d5aad88fd686c81ffa67bd2752003de77213fde9c4a06ee16c31ecb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h281aeeb403b71afcd8bf156fb076e7b9c65442649bd3cad78c6f57023717e7c23772cd685b658f23a4b4987ef2c4dc1e7e82af805329e4b91854aadaa2e96b89c29f5ad0f6cf182cc63e9d0d5f06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1261e9eb95989acbd133132bbf942786f8f327879b5df49c4d67ce336d446cc0de4d3e82b9cd4bc5705539290c69bd0753626168d2c2422f8597f3508654a6384eff65c3a12ec3f61ebbf74070a80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75648d2df46fb8cef1bf4ec930c129d73e11e9a0b6ae512932f8a5f4dfef35c2eff945f0ed772fc60d22501750e8a937ab44dcaad6cd795e080fe22d4a0ba09561ce61a435f5716c3f12f0e75c81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9b359fb591f85f4e8ec9dae30e9d58f9e50bc216ea2ac6c5760f6b255c96b0a87a083d18f7ce228d3d252e7809b4ff43bbe3d2dad4cb65cb0d00d6854b6cdd6aba5dc0b914f25fe3bdcebc96a2b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3cdc4328f34a25227d97e29e64e6c4f02529da788d3559f45625267fdb34e6ec4e2388923a794d51194e30b82b83d0cf638981b7802dede1a12d30161cdcb3c82b22ea6a9665f8e79187ec158dd;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0684fd3077f28b27d8b33e0bfb6ef3c86dfa0628763bf1ede892136efeb8e022da43edb93fc2428261e671dd2e84914273b0627c71a7820759ae325cb8d7b7721334000df8ee09b681f72a0c5b1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e5e2db58f47b1c31cca71737967966fe10ed13bb125429e58bf0b5bde41a45881c02c1b000a678fd379bc7cae8f0d9abe9760286423abc687afd7b71a17bf65f52f3fbbbfa845d9e98e12173bba;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9b741c077c9f6be07844dbe0dcde34241389985b87e61a7cc66d24eb8c32a71a8e3fb87cd9408b16a2881e73c51be6b6f384c922f1d0c8fea54b3f4f7cd08fb49218f211170d251a9079953d842;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1bce5cdc1c042011e4a34eac833936846da974152d688f4dba0cf59b409e49846bbc53d2e0364bbbf7bdf51d15906f3ba9a1a546adb0e817f2c411b521fc1be1e6ffae711a21009c696403a2803;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10425d100b07c2152de431033e360afa4e3040c927218cbc3adf751fd2b7328f05a5d5ac338b595889f6173bcd69b6b38e3dbd97a8ea71eedeaa88410a309f09cfd0786c22bc9c244fad6dbabfe81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h118ce93dd7e614f619342134c9d5d337929cd99233ead4d62f0c3bea4d62f8f1cef6091652725bcd936dcedce02ef1c1ecbd7d90bb055cb88f09c28650e79c43c164c088dd461405964e48c28e508;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1680e427232c299cd80a6e00c8024c75f4d622f4a4419f176f60c14f11a16eda63fd9b28467045c59434169062fb68cd306b67c78aab7186016b9d85b6b52fe5b7e996eec0cfda89af1b3bfb8281c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c4b2e1fd4ce9a0bbc6e0470e40fd98773207566ecde410b4faa0061f837eba9f125b9d8adab755d320603da6f8bfe33e6ccc7fd39eb64430f310a484549fd491c2e0671d51cb450b55031acd45a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158d02c9f36f7c8be3ead948efb1835eded851a629e72b3a66275c2c9208c958e7bb63c911f3d649d132f0dac8ad0092939ae67f98f8d404c8fcce2df17c7cd6a6a0e02f3d8aa514f914257500083;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2280c2a702c3387c3877ab1a347431146ac4f21afd1a5448d8f822788f398e12cc2e1191b1b25f93040192d29e2950019bc980b666c5e1e1120d8425dae92501d4da3d7652533dc44a41e00841c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f8a5cda6efe2dc69e291051e21c35757b3ce0abd6c34082aa126330b2864fec85029b74e780e5cb4840c588a4b7bbb5f809714b403c00b3cc50e8c0a10d52572c207fddbcee16a9a2a6f2fc71bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bf50f0aaaa6beec976e7a81ee59793d1eb73666b5a09e3f31a17392a3097f149d5b1bfc74d515b149f089e7b36606161c06e2c8b1584e0d478e8ebcdd18cde9dbfb4aa23a87a627b0a87aad2fc2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a906a17a788e5c41dc0772a11b0fd2c03892831d7763c81f4def7f1a71ca4a6fb8c07f6999f26384d9f01f300609da76bed6b387ae97b1cb23aae67e5270b44046923801efeda9b02b7b79b3f206;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdbc8244a7e867bd52586d3c2250c682bfd275f4088271948c2f5d58fb8ce4e6aa38f94563a645caaf30e80a8b9f0888e723af22ad6318912a36ad62640a002bc6bb33505e3814858193cb878dbb4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aef6c22e1d085b8d1c448cca6aa80eb33fb6f7e0cad2fdfece3a726eeeb6d21e50404e0f368930f449e05f15c0dae83e50ec9462f261bdde8b58fac914a428b6bbdb778385b5f473f8d5cb7d4ff9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc935ebd99e4c6486b7402f8d8f9493f25aa2d65157d2fb52737536ba001fd3e28b0d9f83c8a4d1c3813d74adb9086cd9bd48c7e032c6d31e8e42bbf2f4af586d59afdc3632c49b86ad5c148526c7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f1fb531c1c7503b7235360701f7c11aad9ce84120ab4b7dd9af178a9f537e3ba2af05e747a7a08fcd7a95260c8b6a10625a713143a2f1cd93d0b953388533d20ea6286a7fa5aca6973e907f9026;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13e04875e40ef905de8e70e63c48f7e1de5a4dc2b452224b5825ae30dfc86113ecdd01dda988e235fe5a2f535f662ecdbc820d8ac617fd04f71c2c73d5a9d72ffa15369918bb51a1eba9e43c2fe28;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dfd08efc1f0bee8bf1e15fab731f1baa0d0b9386f41ae9aa03b0682a632cd35f50d4d3acfc8e6298bbfb8bfa16e0e48fbf51035040036bbe0db5e4ab3009fa167de09cb89dd78ec582e4a8a62f3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5de4beef171078b0c94f684d27f10cfe0f99a67448e5bfb7e2da1effeeb604fa34cbb38ce21d4442c84900faed55293fbf8f1deb51ac72450035a693519cd97a066bba74cf8e74dce3dcc1854a4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb504fa928c5187626ff9533773069fc39db3aa7520f2840602742cd34671a74de550ad6e3bcfdffa271518de6924f957e1e86bd2a4dee5a9e526dda75d3dca558090703d29c9fa47dfc9eb6dcbc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1efbc859d46ccace4ac694f29f0fe04c4a4965aeb7e37a8fdb3fe5a792468f6ef10e4211249245ef8ec2ea692a7f1b8bc08c24b0c142f5cb3551415d05372453b48cc675b26e7fa5e31d3e71c4c15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68876b70482926c11c94c3f5a29760ba1d083deea7e9aea4e66107e447d92995250b126e958b8dbd1b52bbab369ea4af65727b8c0882852abaeba80b90dbe6fdf4b6202df803de0daf902e5878dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb067aecded4b727c89de8feb9d79835f3d0fe13e63ffd4e5cfeda080a98bde6047c208d3029d8bd60a3715ab80e5da3e9d2719d8b748268bcb76e6849c1eadb1c86589b2c5d56f6bf15191a13ce;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1200cba4a7ac801a78b8e70b390c5c3f025e45e84e39a2914443aefa1f849337eecd0c6e071765ad2b58a6bf3dce9829271d1ab6a85ba6117912cb04d4c5495b7b94fac8b872c1795db0e790461aa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15ac689dd13a1159b8611d51db1e51177e678de16714a6c7d36e271cec75238ffcb7f33b1bda7f265d7f8cebdac883a6c9b90a3a98fbc6bf3c35f42684230cad3d22f535d8f3473a49697f4f957e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75b196cf3084b5a26ddda78bb6a29b3b84e971729ec4237e7a382589fceba6d59a446b0291126c833f8594c5650b595726fca7ac5d57d40c339ce2b3b79835c2fc256f59905ede581731a1f76185;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1adf22f909598368d60dc858bccf4ceb5ab35c2c35c581b1589e18c8292f0ca9941ccb9f91c9253632bbc7499791298827bdc6bbf05024fd2f40c9916f0ea824a9c17a7574122271017715aeeed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a47ae63c85d317638036d1003302ad9f1c3ad6011dcd77efa7b36db5d91a67b9ef6b370a756484cf5e3b6aadca0e51741436c525dcd722f7d8b016bd0a6973d88af4e60a1e4b4f7e8d4f79563d01;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c98c12ba9299f01da5ba3eb7d0d3821fd7a25326ae95d423a85f978f2f3702468ea639a2f96eadf9da70957f43d6b2f001d13d10309f6bf9e0f020a9efd02eb563a7c175ac31e0b847f731d0d986;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb18f4be722cd1e22dda5c4a017a3ac845002ebc1d49e9d5e26397db2729c688bdfa92ad6ce1bdb95104712e83cb5cf8e3ecd4f532952ddac0c2d05bcfb54fb6e31b59063ec561499d336c938fcc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a7da37d311228cab36d0a12c93037e92b12d40a586eded50a9d42863a8ef201e32db3d3b9509e736bb51fd762e288338fbacb129e622390257264093d86d675cd5dc9a8d377369e15a25d560e98;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14775ae49190cffbb5b33a138323103dc40841e95158ed5cd335af10137d210e329613023eaaeccedfd1e0ce1eba9e7b64428fa9d05022ed619e7c533151f543ae21d62ad0ff84b7a222f28ea66c5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hffa9a1865f23ab0b3c9eccd83d508b13d7b5b1bb82d4ab7892a743d27c99c702a76375c0cf18818b586569090798381a0afc638a3c920a1db0c0fe111c302e0b6fff07f87f20d7130205d424dfc7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h218586dd02e3828fe9117eead8c93a95d82bc6abc5871dc10c5bef68b5649b44a54091dfdb37b1497531e472846d1009133671c57fb774fc92c1d1775005092831a322343ef0cb91ac257f974628;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h790471d18a21413887acceabb96539fb816861263165f5323b1cf92121e24a83fb0a9c35babf59ad7fd5e272a0364522038064b0930e4ecbb455921e840433f5a64314060b0571ecbf7cd46cf54;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101e10e7c0551d265bc5102bbef2a9c07dfabe2df6cddb3363afe8afd6da2ec828213bf9175ac87416a111a95752699be22d701ee5dff61f7f7d51a9297d6d0c4b72e6b8cb89556299dc39be717ca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1062c669d8d199f6517fda42b73c7e5a2a226412da6830b1e77a0ac59b7de0acc624499ac4cc705e9065e7d1ed79b654a1cfa1d59fa0407fa73251e264c301ce4eeeed895cb562d5a18023e4acc94;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e92e49322073155130a0ae51b53761f765705c59a048534f770f04cd065fc1e1964005b44aa0364a4a32de069396ac9e2208c187246b475c887f0148091ffd72cf5d2460c7005188d59c7231a3b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107e1612f9dab96543b0b070467e0f06162094725ce59aee11c6d4e248049dbf1c3622db479f5ad6b4aca0edf78b91b4075aceb6a76a8c36882386bed2e46ea730a75617a600e9a999506fadb3294;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4cdc978035faa1e6958f23ab6516a5c48f7bf9077731239074a0ee6b212aa14ec89bd0909f9835d1948f1d670309ece396963e2eb92bc7bff6f8536eaea4e082c8af870ca63f69f9c7ee30a05076;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1098fb97cca7e910fed14f9e6783d085897768b06f4d63e8e3e981c627abeb992c3118d7246ef6b5624d25a677c4f0f41b89e37718cbff52e94ce4041ef68bd73f95276f1894a85213dc981ea6d0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f78cac39fef2272fad3f85fce73cbefa6e1f30c542878520751caff79976e7d23dd066ccb83d5575605c82750cd1221796e3c257ee28c75cc3bd0e775cd93cbb2475f4d4a3e1fa9b45a4598c818;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b6effdc5fb665a81c8ce4287644b0a8aa093a4c76586a50ecb5521f4a9f887f3a34be0dbae06de45d9d9e62afa78559a6d97c4724cd52c49bbe08485265d5c3c83a35cb665c0eed991fe35a02a0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb63e4faac61805fe05c51e0dc0a0a349747f2fdb2027d2e4f53bc5b178e1efaae7288cad9cd258c0dfc5e39cfb40f8ecd71f2e6220ad1a32f60c95ad003cf9933527111373930f90fa38b222202c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12566c18901923bfa96e90f179fb953b988243d7a663cb4532f8f019d9cea8f053aa50f24f2dc8ea5bc7ba5f4f53934a6c8eaafbfda405f0d47d857c3db0a9b4cc9fd8990cab59bf491c00c2544cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa8def83e08fbf83213a5f8c433c084f0ff1532e4367ae4888e1ac42138365214225d260fce28ad93605fa232a5ec5859b5cd2ebea07a182ee24c9e292e7b2bddb6d8cb5dc89d37cb764f18d01bc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107163ee0abea70d4319721ca82a9b0b00f0ec3dcca7410b6142afe6ca241dcea590e6bf3c2a0970f93fac0545e36d66759f6877108d3698eed1405f4bab052c6439a18b433c784095478cde76028;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1322d56803c7de4c10143d419c868c505c001467105d9097ef9679937990b8e6f1ae78869ac388ba65872b76654fb2974a8bb83313d5c5be65481839414f8b503ffbb13438845bb91014e0fceabae;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f1c8c1dc7a930ff27045dc393bbfd89046808b24b21074ccac4127929c06b9189bdacbf724596f0f38debf3f0b6ff3326c6881b4baac8fe93d947bf5442d750e80debda0e0a38473def9345dc88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef4376546f3e763f1c9f0daeca86378d72a8b7f5b1196df738a98d23f475907656e67d9c641ae589f51108925bee071c7c1dce5ce86dc8f2f6e5b43bf651db4271103ee088c7b1a10bc53528fb1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf27223f99ad8b781abbad399a140f22f8352619ea1bdf8c50f4a49aefb663e9a6f9ca6ffe3cf27e41a1a3f7a7730fa6414a8c3e9744deb3fc51dda78e3559c87cbbdd67ac49bc4a9fd5c074ebef4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfaeac6bf7b7a4d2f1983b5b807897809187983e7a6ab22f05d6e020bcd5add3903d9622a1c107ad1f85d251c83d0f58f53320bb400b5fa3b20906aeb09df36f1744c43eff2b4621518c493624573;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e76c40b554ce1403cb6508f42e92f15f9717d5b44f91fabe4fb22cfbcc4276fa4a90dab407f5453e2e8838c262bd653d57f57ae5ef2ba819e8c1bba7bc9725f8bded9d0f12fd1e6105dbae5bb723;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h791b7d7491259c1ac0989ba0c53fd6bd882eb988c0e7e90b4f98ce1ced13e5de68b59ffc346e2ddbea384be73842fe72053496fdee9637e12dc575de6228431062e7b7fd5a4a9bd260bbcdc1185a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d747396ced94e787d83dc1c0654fa9a6457489b71d54d48957fbd420379ab7409685f5f59b4a731a46175f2990fdd47a22d315a36257af05729adffd5b1f715edc6dc9964d98ffaa0a6198e14cb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d1402fbd1467e62302eb231dec48ba54bb66e6520b3fbaf580f37206dc4c0a51bf912ee1602795ce4896bb2c0ef5dd0dabdc9864e6a43d76d4ba262e65da28fda526be63889e953cb7c99b687a1d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb704e8ff555987dc19e5ba0ff60f7663126384b644753b66884db99590975d08bdebabaa82ca8627d046804857501990af790c1bc247a1aa5202446929a8e98044f55c3e26451384b3d014c9185;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137d8ddaac404c8dbad2eb3d56b086851129918e16393cb6e9bd32bdcff636ba05c2f433ae519a62773b79c9ee7ad557cd7481f43964d92dc416a9cacfa38827c3b8ae6f2ba6feb1a8f91b07eeb56;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb5966810f388a9482a9fa2596b019f08968d32039e6de81d773e102a69cba0198e2494c6ece19fa805b924000eb9dc481b759fd8be536d9267a6f9ebb5a058498379b3d0b0ce5679c99c1290c01d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2b11f171dd2042cf959682d69ed2e580a71a259eb96daa335a87b165ff3015a1bf8525cdc83d16b464334f46c4f6570db0be9b9eed2ede142b6954da25cbf8428407042b00f386d798d38ae162f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108f0c4722a408311c00af2e0a1655ef49542c9576de103e39b490d4a957c03591623e0b00f21b74592422a6ed8c2f765234599b05ed0c2b36f87e471d2957253e15eb5cdd3c662313a440ded585c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f8a9e39285764b1b03db093a782bf7cbba0f8b02fca7318feccac585d917fb3dcfe62165d7ee68210f02dd401a0194ef342b4827eac7738eeccdd4d6a36e594faa045c62711024a8d1840cd8af5e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h42974ca095b1101513f59da9f8e46cd4e99aabb09c68db29c80652ea50aef90692d11d5ae7a37056b7636f2f040aaeb8dce7887b29263070d53e89579ed67c38f9df5f162efbb761d3fa9289eb26;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ded5919413a378886aedc2b5bffaad265871d7bf6fd5703e3c60d6bde84f6494f6d6665c817affcac18c55efd50b2fd270411075da7919c466abefe432528efd3793cd86b9a56e79ce54b1aa7ed;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14bc54bd5bf9969b5d5ffc01fd4ce09f62fc38f9cc7904e0d95b62e054aecb213c5caffc0ba9e03fa8619d4f5a33e2e10c0bc365902ea56bb6b78e405673b479d63923fa93cbb397082ef30983983;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h65b36400ba49631886db3e8de3b5799e9eb8428c936eb382fa1db421146ef77a6bc3e39796bcf8e5a91a7c89f72c480040c633a32e024c973f9c30e4e0f53d284075129d1474a04cbc3686b4f4e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb103375745c563a10788b97375b27512dadbf3fc1efec479b09ac6beeafc97b81ed92de81aa1f8d3ba53f56094f9e31e8c8c01a1330370bcb63875b2453b59f96bf0bdc6b5e4c8fcf1538400e557;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f59d54c5f268f4127eba9da0973a8a26770265b7b645de3ea476bbf383b0a5420c4ef12c3a870fdd6254f5847e1df53e6ded79758a85bbc6b0b04b3b11345190b314ead6563d60207cdea02516d2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12e4a49439cb7e9b5a3ae392744ffb24af910d9db485f1729558f11b9be4fb364e2174af36d08a57b4ac6ad922ad00a927061052e1d08d692df8248e5602114d8de5c278760b720e288515ba157da;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd4e925ada08789c1da9cc3210a58ed7c7ba7d7f0ac13f16b71e2879745a6a597aa01f4072bf65fc602efe67727f738a7027661ef1e1277a250ce5740d6ba8dbf20d3d68949fa67e3e16423cd86c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11db3a1ec08f38ed5674d008a8231c648a34d18aed1b574b398cf3b8f1f33d508aae6b684046e24815abf4e22e4b735e1c42aa5d4f59869df51c9a87eb17ced808b6c7aa6c6ee9895577aef81d428;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2b7d3814241c3d57980760c90d18b91fa72bca5790a268786b45ff3ce40c03dc3987321b143c28f705fb7628e81cbaa9b127518d3fcc4c8452fe9741b8253beb66e3311218c910f546cb1bdb83f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141e0be351e534c4ea323c1c63092336645f01ba6f4f7c9571aad8efba336a8d9046faa6e48e1a03922f0f0fd13882866c10b4b085cd631a3741608b46130fdeb852ebe1590364c0c645a7a2a13db;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1133c02294cbd8f64c8b97e5d7560a95ed283bd8548524263a6eab47915cecfc4e1d3909013e97d1bdd1dbccb613d4d0ff4bbecf3b0f89aa413e6b3e72b0b8152bda84faa66d643343f9edf06e249;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56b6d11a3d232df691723ee54228fef5fee4134c82497fc2a00522bb484b42569d0775b9908913b974ea816283de52d2456bdd0fb54ccf142420c315a13ab9cc09d19ac38b37eef8a83d7ae7c151;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h618a8eba10b4b3d46650b9ef1f355bb114fa2ed621dbb1434a9ce698ffedcfbe0af02d6c445260f84c9f8e4a0f150fafe647b9069c341512aaf0e946e897de6ecee8ebff180ef5593324cbf08af5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16921d71e648f5482accf0301f87b087c7d761aab9cb392a28a30cbe579b2ae06ad172b6acc968930cd118e1c02baae9453b7b0484b293eb84e8822791a04e400d832fb8c1b881bab1914c690b2c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2643bf7daaeeee64485f4d696be0200cb4d0cc88ffd87395f38ba87af1a8f5f0f15aae483745d7e02ff7fab1f22d916a660f2f6a2794d046c2d55a574242614dfee09e16b6067986201c637dfb5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcea0a7289c7fe0b3e36d3de878cde0ee32f1c96a06470759e412dcb9b765ffecd050130f9264c734e73e14a3188a87a11824b96c86e4db379213d81f856eaec52f60a1cd828c94b1c8fb4c3cae6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h671f532c006f50ec5a0515f959ca95ec520232a1f14a5974157f2554f4adc6973a139a9d99e804cd7f04fea8475f4bd2656e41bcbfb603012342ad4e4f85b7fc6ccdb3c99cd17ebbb3751e1c3bca;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e63bd4519c63ee9786abae3b455e9ec2a95259c62cbed910dbe223e4084df14501931958e0db0f62bf6ac66d08f8bba8283308f709088339451cf1c991577d317c43a6e35eea561b407e5a5d9766;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h854877b1e7a3b856486d8f8b070a50cb36becfb1c14cb12d89a080ef366fd978367015802cd3b83567453be2d765742d17301521c6930f3ee3062a22bcf0f326f8b9ff85232ef8706c47c4631784;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c756254c0a82af697fc45ed1741c0ae83d72aea552b6f7a7abd021eb433d9bd875ee93ad0462a7ddba42f82d736cd097e852c1c5476d40be59ccc7bbb2cbdf88aa5a16b86512e02392ac1ae7f4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13165358c3770b340f5de9f2bb9a789604f46af91b925360e6aac96aa13bf8c5c522a5dfc4036992550822459548c3c5b842df28c01ffca5bb7c65a3ab6911aa6a36a4598d4fbee35d8fc871e7a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f0bf857f4ad818ff989254d1f4759e85fc948fe150dc2ea66da377a6864231061cf5394c46dee08068bd94308b3991fbe108a7227a415b320e46f225d9e9b0c6602cf0518efd9b61927b71c00c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115370e32c5412220d7b0c88d883a16b95bc068c01c48ff96d958c2903b8f11f433841372d016ff5a9fbf05e4a0a93240e0f531abd3177384a553356a338f0b033a8fd6b2f3a1f96a847ca66f3724;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb376f759d130e848b2c7a1ef3078ef26f72f34dd433e1b1cefa50554b69de16c3d0b4d57f95c67532d561b0a97c7ed65fab55998f98c8fd2bee1655edc2d33b78e24ac9e3dea0eb90777de788e9a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf3b912db0a6b931746c18543b44ac39460503141ded90248cedde5ebec603659808eac874925058ebc78f44091519e7a5ed4e5d1b4aa2e1e29b74df5d86cc53ab0703a85967d6c76ec61ef2f470a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ee58b975cf118988b83f774a4026b020ae22ea13aafb61a0a59086a20404d83dcf09a2b880d5224cae0e3d77d6ed22facba1fe22dbb5c09a94cf80e8cef9c16145679ae9d972824ca22d8c55a7d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d48c89c9e6ff85f83cb82486eeee350106fbca0f3a5aa0f242e4712d3dd68bd22e7ba9db3008537e07596e486d69ac7d1dee0eb0d73c6dc9a4ed7d063c421b37ea9e7dbf249da99b204cb65d55a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7850016938ec86b8510d5ee998cd366bdd0f941658eede4b4d46d90a9b6262677782c732e7676b0d52f6afaadc98cd54e932096bc02e1363e6bed27a3e09e79e5f8dc61a5f81e0bda4f834b7ad80;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h22c6c397bf77c3ce0ec06db97774a006c7e328ea055be69dda8a2999fa78b2ad15cad4ae8fb36ef16a8bddd91603d1bd6dee4d0407194bdbe7c56323b52da5da845a0db4130127cff8e8d9753b9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f79ea5b99f1d3a62fc2552d56d56ea02288a33bbe24ec706004c581afb79381ad7f6754d9065fffe67272aa02a44943f7ad58f4434c03d841b76c48bb6c54c85883fdf17aa657bd4f94746c3eaef;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7b63a34ed5fba6e27effc1d7f211d9fe153837149604b2d551d735a85a8206d0384707a8b4afda2a123891be498468dfecb39e9879d9327aa6125f649fc15349048232023a8f092953678740809;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a03419db9f051446e5086a113cf6f897d201f160496c66f1bcf0d224a9384367862dc923ea3409eb751c1b2dbc3c2e774de051ec08601072b54f65eca52abf114a505fb02f7cb9301012fa8a594e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b09671bbaea638dabcc4b951e45c6f61cc563c90fcee2348775b7eabaeee8ab0366ebc1a3c8edf4718869e429e201dddf9ffd214682f7473f5278ee63c35afff87f855d3dd1c8a739e4cbd8357;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11450237d87683c12e6e19ea0ec7f7019ced88ff8c68c172d052c3ba59b36add9c7b0d27dbf1315e332e06564b7280097d4350aa283e229848def1897fdaff7243d0a2ea033dd3e960ddb3e3046d4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f5765d0ad1ed558708e978aa2a9a6ee4019eeaf0a684cedc419200bd4c3d6c6ef1c4250d10b8b949d06111bdb5f0add758018218075c2fdf8d8d3b453aa90fc842ee2f7f0bd3f87659051b8f35a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7db8bc828170df241acbb11cbe750d013e94f959b8a8df3532c22a9f712dfe5388f28e172ec6f1f928775d9c0220f470f9a6d22d75fa90b91bde0283c8fc4cbad99af604182dcdb8ee584d97e0f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16bc9aab243a2f33d5ddcc954b06a0537ca4c19347ee27df0320faad2d7e74ed970a761b2ece25bc6b7f4bba7a3b1bb217500ea7afa6b641fe69f70c18d227413d1f121f452942b8a10bf0d872f6c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha06118cf84ee9c6f3ff1ffbcf2dd90e79a812a4fca8536c59056ce99daac63f43dfd43860842a4dee8dbc4c924b07b2d122b5dc75cfa6f23284a4c42ec4c87b3812e19affa6dfb0c29646765c3df;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h894d40ec3a9b23f7aadebfb2a7c8734e490c19a9cd8bd62080e27682b66bd2d141dd1c2ca7d14974c918f70e9f9895f867c44e80aa16709f68130b8ceebe2c5fca29535118fbadb1b000a723db92;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19011c0e0e5195b8e50a4223ad6a367a1802fadca2843efbc4b060b16302861e4c0c71ef242b7a02b2b2af12a56fe4c5ac191848f6dd6e5b71a08b6063ccac5523480a35e9a7d495ad064c3d8a6b3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4e60b6f1a4ecd3e36535089f7c685ea6b5498747d2322c766ee1f653239040724cd4b6822d91fd21a8b946a272a1b441ff58d3ce5adbd389b5803681c92204940a7c115b7a4ced6c6551b054d51;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161239ea858efa384990a67866cc17f144713be2b73c5a25078dea859bdcdec0e58e55d9e89e3d83ff7e733298c98244b8117ea8b39ad05e1eae4276213d4d6ee9508ddaa7a35d40dceaff49f2ba7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e39a726ac76c4f0e35a20d507b9282c19b7dd4904fabf423a62117286d837c1ca375e422cc52cacf1c87fa1e7c81aa51428067aa6a0fba2023fe81252ea40dcaf43636d2dddff45e73f7e8e8bd63;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7bf93dfa5f53e2b180d7b06a07242acc925b419bb0b1e1531fb30798b7bf11879cdfdec47940f22ee5aefb1bc0abed66e9718f0f691964018d1e48e10430bf663bfd27327ea147571a1baadc09a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0596cbfc0f6723ba0f0760b94d761bd195bee7ed90715d420395ec03e721871b98ec4d961fa4bf3aef6612e384478c0db553da5c7fbcebe2521da1f61c5675cc32680de6b85ba83cb8927ab8fea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd138e000147095293138f2fad4c0d9e5e15743ea7a15d5e76a46a438fdbfef2d0d7aa0b980f0745e5bd365e9ceccbba8a690e2c31848b7b091129f9f4f2f567c58946abfd94f6648b59ffa877a42;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d5047bdad6cb8e156ee75c7312f19144bf032e2e1aebc4a320fecd29590837ee1a91ed34684c70bd1918b5457ef3f53ffb36317584a1b3266eb02fdf83ceea6eb848844720a619681d9b3590e1b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e26737b9669fd1f1932ad019630bd1315efa4820d1e8f670980ffe464b4832cfef68ab19b7279dc4a49d88ac6268a07368a08290bc88a775db8f27f9a85497a1b6d415c91e0a798547c50f07166;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdfebef5323d0e36b4d6e0cdb26e154bf62cca29980696cb15c2ae4e8bc78e03eaa96103ae68bf66bd5424aa5dd117c18fee09ff8add638d8450ef449fa193efb38667268781da1cadd2228aaff09;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b8d7315d6866eb9767462d74ac62e3aed823881fd914f1c8705a1c59ee43ce581cf7f3f757f6c7f5e2d01e6d305a710434fbc0e79483ba623edf40a7ea2833d047a9748bdb6620754625ec78b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1480a7a0a3d08e5a41e6d1bc56493813e1c97c6366d529bfec7e07ef8385b9975aeeab71b0dad527cb268e8ca7297eadffb83977132c1ce56c57a404391ccb0df6f11b46419b36159bc865c5237;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hca5fa65a361349c7c6de4e7458d56392c7863a04e804d8af7d4ecc3fd5f80694fef0fd750fee90b7dbbf2b3a1508fa2519d61fb97fa4c00f1f05908b4223feccafacbe7c106f28c56676670987fc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f3ed2f8e0f398bdb058dd99153a11eefc544cfe3eeae30f64421f993c33df15f21da588f04ea9a67d666892e4ff03ebc334f55a453921af514da3a82bd88b30d22f9edfcc311de50b24f7c1248f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cec711547b8b1cf757308e5e937929a0b82016fc1980dae84271a25486efa9ddf58fac0ea6754633cdcbe19c9d0a6631582a43bc68b7bd5925517c6aabc960e44a025615e5f79d5b29e37e6e9bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h157ee15a39e4ed23540002ea102169e73015e6a9ecccd494d703a9add17be2002e1ce6176b9195eaaee2b9e43e9cd5e115b138a1fab1659c0b60d77f87998dcc066c3ae6ce54bb797a995b52a0613;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3e2a3de7ddc2c86b0f05ca820fafb29cb047829525be8538136096ed72d99f7a4ae34d4280def3561f37a9814b7b3a91283004eff9044f2c0c1020c22ed941b153e13491ec14b0bccac3a40f43f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e19751d692e723e6c37c6847c130c0f9064388baa875a51a732f0d1e24405a1e1debc29bfab2cb1433757e98caef99c86715f468cf7a4416084fa85142d83f3db84cdf072ec0f19d3c8a4678d71;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9d1159f96096102e6058751c7ff7d81d0bf849c7c1afeb6996e83c3d72896c109aa3ff1b27bf22886fe157b88838b2bfb0dd53453fbc593dfdc901b7f413a2bc85940f5616af7c772bb4f80001dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c00a6cfe3817acefd593e3745b1853d38e4df2c71b76fc0b2f40cdc55bd2817e1f6e1abf8ae616ebbaef25a52ea9369ecba19c93c8295fea3c8ddacaf263c93a7ca1666ff89179e14abde021a4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba7d501425d792ed136745d19d0ba9e39ddf8bf5aab03e3a47cd8cee92db6970a9d40816a52bfe383aec87f4067f27d6df9bd2e77a9c09ac0643346d424c4daf62624643396c3d297b60d4c8930e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b50d9933cf030aedbb88059d01ce46100daf4fc6e69008b64283ae06d491c586ea02f69988d7ab964fdb49144193ea7f3dc4f584400679d09a419f2cf194a5d8a3f6c6833b034193b88f5ba49d6d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbe52fd141cab44d4f1a6c7e274bc84ff910becbde4997712d97fcf4ee7fc692afe529c87a34459209db6386e1ffa33a7a80ba15e478e892c2ed2e2f26d1f82935c5374ef787250fb076611cd9823;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3d4eb7bdba070927be5f5b1a49cbc5e9ce36d72e1ac5df454d1801c75b87bc3483daaade5c3bf92dd3a786969254e8021a0c18283542b4f35934eda4e1df9592304e2e72c0488e4d432b167566d0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf348fa846afd3f42dbb352d92ad6f35725e2de4000dff9cecd76667c2ade237fcabd3a1f44f586d7ea3b91c1e187f51d34b2f7fe4b4ce30fea3affa5a5d4cffc2495b1605b8933127710dc81103f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h39727dbe431d3c4c0e2a87e007ddd7e50dce52b84c5e777b3953779060a9f562dc34531baec344cbcd7eeb63bb872182f470e128e407c0a85e9071b0259fe8d21aec5060698261ec72dc63ccd3a7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f351e2997eb59c6090b3ff68008d3ff4cb8b3f09774582f190fee662aff95902cb5a021dbc3ca2f433c0db332974606f3140938866da39dfcbe2da7be9ee6df4e90700a7f17fcb15c045eae10252;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h378327ce0041c51fda45741ca972dd875c814f3c53bdc2cb2b57e50128fffcd2cc1371cfef0dcdd4b358e33029b17379995b1fb2b764ea92cbf4ec62446410551f4f960a0a9dfb7ec42658331e45;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h670b8f99bb33949f64e10f6383d2493e3c4b544fb05f93676856d5cea77459ec9f066c239b67b5db3206f194f126b859b65cd182bde284e92ebf8623635ad5bff2dee13a3cdff0ec42f14ad7728d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a531568ec64c44bc90773ddaa1ad8336bb8f48b15cd57b02e489ab2946add88938e64ab55e21de96fcae93c537218653364a115b6bb5d303d50d9ae802a83ec758b96afeea76ef3017ee537742c0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha53d9138a077a264ec3d24e56a2d3139898f5ffb1e0916ba4b285d75f860614656dbf6568bc95539e6d54ae2dda6eff68f42231cb27ce13aa8e2226a073b7405f198f789e2a95c2213af8a696d64;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha12b2fa6348bd20efa3ab220eb073ef9febd9702067118c105d8594a488ef6159c964c2cd25765be91d5fb46cf1b46bb6f4d234fc4c5b829c4c996f2762fca9c0354e8515f1dd01bd8b5c73ad3ee;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12b02015173edf71f8d13c276cbf9254c05cd8860e43805d24123b61f43d9626ad902ee69b0a754fbea9f27e5c35aebab7fbab91c238ea9aa2d73331add4a00401b718285e6e00d873564c85cb48b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35cfce020786eee87ce86b2bd30d6acab7eee826b2681cc97aee987dff3420368337bb9d8b716e3507d34f8b197ca55864a2c5b85fe4573fd63e7ab73b1a948927bdaaddeeb9ef6120cc397f3608;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1a05d568e2cb2a3d34a1f6abacc4bb8778e360392364b95f23dad1e6717dd19f906f292846c7e9f059525f0b41db577856e76156bd7481eddc22321356af9c375049f5263a0e768dec38f35b3a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17966b22f073b329261ea504056d8fdbc0349dbf48ad02f00716be524292832b99aa5383b6e5528c1d16847ba01caaa18d13e0a03e7b1065a96b152417c4f83de9151ba6da1b286dd2a1f75bd0273;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c6aa5f8fe53f34d937b9dbca990f605ddf19db189c50fa7f75c3abb86c64728336c0f66c89aa50aebe1e85c10e641029a700357f9f5109e18e01706f8ed12696481c8a2784b14febdc338d673d1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9828bd37ec8a50cdb2426031ae6877fef8b178462813544fd78c9cfbcb70902eda3a9b3471f7ff6813e4962560335cee4863880ca9ec4dfee76b18d1387a6a837c7addff3cc0d35f52a486aff2d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c00ea727f86af6b080aa14545d21894cad0346e418bf47af9ff59802f4b58ec57ef94fd975494c8f482b0763c494018731269d20fcfa6f4ad8590cb2211e77a30acb6aa369c8b4126e43064524d6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10724f254c6f2bb90cc026f4db929cf1b3ab0f53c6edbd1d5b6a1bbaf9eb2001723d82728ead238ce88d2b29db492f2cff998c7eb2ec351bdcb26d24e5c11699239164abd494143a9e1816847db1c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fbd8c8697a75e29f782093b67b409b515040e5a864c0107f70eedcbd383dc40e8913531cddf87f27b64ec71011128e3243926dbef7898026cee274b09df0ad570fbdab12769f39d19730adaa121;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h757d184735d063fe737c35a6f5e553c094550a664d926a81e039bd25b20bb8cbb0cb4ba122f93729ab78d6aa7f711601b443829e9b1aa92fc1e444612b1e85667cd774ce3614bd6016aaeb49a2e1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35b8000a5e863b958bb9f125f4372adb7fa79116ba640f9292950c6caf6cc3a33e7204513798d41d46550a524289dd657529bc7aafc95b017ac4a041022b110459c84b42e2d7f7c8b6e032adae7c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd078ceb1b194e494d5cccdc5f04a4c45cc3a4e0450b7c9cd9f1a9234fa8e6ec493ba9010e24815eaf1b4c95316c460217bb124fe82e084c6394527cba823f83667eef0ee3a49e6ec52360571520c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3339a4eb89029c03a2054cfe9bc387da39028d9d7c65a57e1990c2913398c1a175577e5d67ff7b86acfd545b094f52f58acedba72bc6101f9053ba95d8b3fb64587541b8aefa0544243c1d384f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1beee1b6a5d81f910e02713054c999c768ede87129196b793365482d668a56291fe23402e8bf3d9d6d720a9206f4ea953c5874a4a20e5b1f2497e0360e9ad6a89b76e5313ebfd74a27e8b9fa7b191;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b24daada3ecd5e16aad21507ccb2679b69533612ab03ac0613a4233c1af9b6e65c38e943bc51f9855b940cb10d00db0770882d8c45f7d3e84f23fc987708df047bf559d71a6d5786b077c827dcf8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d27cd0582ce0f7b595992f71d6795bb108bd9c7842bdcea5a88776a392848d5b125086a9c471de9569f5012645e2daeed1de8022e5f93c54694a173931a44f946ecc7b34867111343443d450f3de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he296558d7d1c733e92877f05ac9822ed358612b8b1a17902d86abcc8730d85c9f6e54827b92f2df5a3b732be87d8edd27fc87a1ae1fd8b10e95230f84774cd84b56097fe1b29ccc5a371646c2443;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb2f7c6693caebef0654056c178459f9936e7960fbba7a67ecb4a1fc3251217738f288218f3bce7fcde3df7cb0b58761360488276fa6f71cf197c2141ab598551a57aec3b606acb655d07780cdcb9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e64c3d5c612f5993e86d2a53ea6d926cd877d291f4fa9f84dfcf6039f72640ffc36ed45f858a2f6420e2a34e356c76db2aa38de9be4f70bdb212db6cdf4c5276d16a772e21b8d6ab97ee250898;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c4d7cb305eec9d4c86fcdd8d0bcadda275a5573a5f6062c3c321bcbcb3671ddad48889a8882f42ad666230513e9fb7aacd9846f33dffc3fc66cdd2d276aacede343e726e1f9d84f67d01b4da185;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfd1b635ce70d6b9065a22ebbae543f37b861c8c112945cbcf6b9bd41174e29a08f0f41b0eb868416158390bbc2a0f074407865ba26ad23ed7c8b37502a481f342af538921e78327d1b4f220d8205;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9eb5a18f8c2c4f7d502976f6d420e2b2874c506eada41a40ff6606dcaf422570532047f880b1bc24c46d7e955b321a1a69eb4fcbcedc427e1e44fd40da95780c4890fec24b0ca9a54d1c648ee890;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h376948262a4841639d2ae94b8fb860fed98dc9fbf7a82f36ed01f3433e1110c106675bec89fe3d9a3330a2d9fb58df59b9dcdd78843f2a7e7ff0a8ad4ae7cb6e1376bd374fd0a1d04f5ed1e950b4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa6b1495ff044df0cecf6dd8a9b7435f5f6f1ed0032d0925f698e40819150fa28adbd1d5dbe5038302c96d22010e6777eb44fcb8be0a885cfb54d2d32b74064beda136f27dabe04c06268cd20bab;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1829c7ffdbc25af49e6558ce3489071c012c66d4648b43d76d417ce259bfc61ec56e8a84065217836ccb6309f0700a631024ca6b739002fc2c890b3b8f4779ae7043117e19ec1bad1ffbaf35555a3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he03a27e92e96db30e8f14f33f056063fd857c17048f83f01b537035ca6b0b972309e61d7675daf5c6d12ccf0ea641f2b11d26ed3cd02983413a13283e70b05128a9595040d34ebccb4dde8902bb6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab5c6606ca3cf8f2523ab1c4b4a3c7846e77fe85861376d4a7424b912fe368067c5d59fe793ca45a3c0aba21af6757a67ea6c8385a6b17aee6e81be7152714c20a4685e79903856e31e2c18ab141;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcaa6bcbc4c2271ea69eb75e9b5013161d85b2e92b2d9e88de9f4e7d85b153ffc3051f8f2809bf8233c3d16d93fce09a320610945430836aeb25c69c0005ffe8eb72486fa19c03233d845868179ad;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h438461afd9123c589f18008cdf0677f0e8e860f750771eb6a3d4155e839f08f83d324b8aad8ef0b5eb09d7547f448a963c2e733a515e93676b1679231e157bb5cfdc131328a7ad74b23fc181970f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c9f1d0ad7c44d37ec1952fa96894078cbfa53ac61f5e964e6481f656c140d6a73c52c3fd601f6cbed819fc519ae622711b7f270c81bf2917912873465b6274144fc8b7fe8296587299ea6b8e676;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1c385b3667083f66c28c1cca55b1ad87810cf0dbf84604141522bf28227b4923d56cc61bc1f866aa14335b259789a300a1d5955aef458ccf491617f2fd4c5b752189ec2c17dbb2ea490b86dafd1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17392afbd41ea81ced85b09d7804675b7d8ebc593eec0eb6aa934703321ed75ca9edb2d04c3b2996bbfd0f2906f6aed6aee56e1ebcb52c9115454d84d6778667d3bac329798597fe25eb29326a406;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20678fb52a40d075a929558f23090fc8d2d26f59cc36a06de211a0219cba7f546d454ec20d12c9ed21fecf57ea0a2f50bf0b00f580126b006406e344aa537d67a6ad7222b577e7c41922fbbadf2c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1271c02092cf226a748c29935b17cc681b7b5ae41b9e1ea14ebe0ab62ddbd8e8a672633d4fbbed68ffd9995683f658d1956153fd92c122ba5d7c9e92baf34ee17e16f4a8ab2bda5050caeae8493ec;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c6acff0f362fa07241605fceb7eb0718ff72a1637873c8bdc2329a8203841b7fc639d9f13b690e1894d6eba6e35a4dc331df76092afd36a02d031f73bef6b132f921b06fe4def8bd500589a43de;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b9c6ad77a0305253fcd1d53e43ed36e37f6e637befae239b12e60c3736dc6c3d91641f8f7ea78e67aa8079499f2d52bb9df1779f9aeeb3ad2cdd8d5e8acba2748ace96b165bbb5dc3f0fa413dea;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h181045c42f465a17f18c6708e846491ca8ba6cf807e60c3485716afd2bbfa144283d9967d51515bdab98a40e6d0632ba926ab384a62fe5f413068e252d40d861a34efb5ce56a67ad8090e393e6b9e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f0a754af338e19946c77953a7a74ee86702328613b94167d6b7395ebf2b5a5c088f609b7773f1cc48c93d2b3dea0aee1dde51e2cd35be5d97006123e21623df0ef66daa53634316493e6dc1e756;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc117c4441934d15eca6a3fec02ae36dc69063a0eaf4964efcd1aa8d35811021ddf777d70592ae2b1d3d205ecac1efc3c5675a8400923d13a85e31afb3fecda8e59bbfaa71e8052d1c17b7a35afd5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d8c5a5906494f2edc187c29f51c2317eca7a130981b75bc4a6ce939a3e7d17be0e4eb6d1f23ef0cab45427c931223078225c649996acd1185ebf3083ac662aff1b9754af1ef5ee2e53e0ab8bd77a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107c497e7e97b5761d14f22f7e77ace750c84cd37392288e8dcfe407ead60840b54ac1c02560e40d16693f470eeac9c38beb02847ba337cef8d11721cb99c0bba71d4733d2cdf6ffb0238d91c940d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea46a6922a5cd3e3a8c24cd50abc0b8996cc733b33136f4042bff3630664b69289e03b2e3d1d370f8f1a196251c89e05f6fbee423b311ecde384517096c6ae05c19181516ed11a166f9b72e24cff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7f02bfb78955efee890df188d946950233fc6889dc6bbfeaffe9d902339cbaf1fe93799737ef57c177f497301c5d719317248d113d6e6f0d669771899432c183fb393ac177e736b0a140cd653d3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h186b96dfbec39301c2adcfaa0119a8b72fd1b79056cbd9a3746ae5113379fa194e7df19bfcd8c48ea868164b6a3c0d6585bd31eeabe77c72309ce00e92cb29c2c8fa2163c8873da4a4e1bf71e6f30;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10af865f806fbb81d3927466512d513ab26b5aa59fc5a0173de6018963caea4c21e921c159e45e1f4ab87d5244b24428f0b0ca5a5f461045869002f6057f7f39b13a3ce0e5ed63b8fc9d431cee29e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha352039063b1d4d115e760751aab22cc0edb08a12819e92338782dd2e7191da1a5f2615c1ba5c91bc33f21cdece97a0ebd9b26c2e1251ca905dbd44ecda36e16d87ce05044186fef592ba2bf20a9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9c71df0c353b296ae0d71435a545d956709f1dd5aafc3c386555f4b857ee5891be66fe1ab9ed4afb7f8082ef83a96679ced0636453827d500f8ddeb05034826226fb349bd65b7f818e3145c2c5e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha26e1da06a963b1f61aaa120e6fb6a8846ab3e5d91b9cec727ae1f3684796cf330670794813a447d45b6568b19b36cf3d3853e0d0fdb666ffda674ef4ee0c74b74466679bf92cb4275947fa3f8e3;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195be467b94ae1b93f03eec3b6d960a5181d8932b493031d2fac337a6ca2224064db6c9e0ac4e3d9c338b550ffce9d34677572ce74ff178e62c5aa0e24df34c1ace548633e48d3352ac2d2e6c2919;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48afffc8b19b004d2c42a80067610693e1bd0b7e8c2bf2797508d64ea5057e9cadf0175267f69144f6e03032891ea45642d727c5241ceb0bde8aef7431a6e1ce0040cef7276a119e2e8b601e9d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c9c8442831a06ef94436f5914f9b1f55b2f41219cd3447f65418980b1cd65bc7cfdcbc7191901aa9af1227f84691b615f02cb47509a58b2b83154ef3bf43a9261de9046476734bb94f87b63273d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110a9fa7ec226d4a30bb3fa5e6e9715aebd742923b2066160aaf0410d15912495d03b927397156de97e7401350b1d2a66cf51b46821065e659487a8f23686005d2af5e6b7da60e83aae615ceeefd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f872c087fa6dc52d598b0d155eec8db4d2503c3ba48c7e33e1d3c1f9d1ce93fbb5856f9bce5ceadaa482019816771fc3e4fafabb6ff2f440419cf34761eb7c9e141f75994d53dee4a4ba1608867c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56a18352c12f30c5e2a84d82a5bb1d68178a65cb200bdd9deb583714e38d17e40265358796a7e7bfe0559d706e437cf3d3ff311ec152b7544787353a801f2916cca5a6136b4b874a75998c2562f5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c32ddfd03906183bf412a6507fa3a95a9347f5bd3ff955de0cca49fc3706eec66746c84c270e0c0f206a416bb41956b444e297edfd572273b01791b95c4e0053f4d1a1823df4879d0b318d655cd2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f0d7582ec658b10b658e0b88d91f61c5ba9da83d0e8b639e62bd36c2f4280a44cd3c723000ce3f13871759d94a39a5938f82b8c5653a7c3cc81ad78d01dd8525e0adab326a56358263e5fab60b0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1356cbe3d743bd58886dcc4846d564b868b259cd0a1941aa58948b3418dfa6c9bfe741f09f6b6b1ea782fd86878aed495a10779fdfd092596fd97c55f8b93d7fce64599fce1d15fe9f729d6a0759f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1279d8a8a343269d1cd6e220c687c5fbd1213ebc5480876986f6fe20e76e211fabba5c4f0dfaa6b76fac3d7e8912957340ffde33d26a38c73b102d4d80a7fca047f888ceaea96d0d39f4923e28fb7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h33d1241e442309d5903b0c1bf869f32e032e86e19ff31fc8e2e72023f63012a2109e254627fde0a0e5d7e139125cd254a0c624069b52c9615c6a2c43bc61d3eb8e122a2ccf118a25405cdd0e5de7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha519d2ccf5e3c6bebe1bbd83c1d80ae8e1f1186cd3970fc203272772cc39dfcec3a6df8d1d4a3ed637f8a832f4cd05782bfa44a275750466b413ba2f8c90c7b45310a0df86476aae54905b5929e4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4af1b35f05ce18c72100085f4086f62782a06f88d13f48c6b62331da01fe390686c8935dc368d5477246954265c727c8ab0a8bcca7f6d93883d1504d30f6fff0208225eb401d732ebc4e783fdde4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f89524ff99158523e0692b5eb5baeccb8342868aaaf1c643741b2d288467700ec28deb6a7be3d3e3d4f5a63e876d4af46e0c660370ead6c17249788654feba3a81b6ab74181304652be8dee7d944;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h472e4c661db3de86f8415c8a997fd302fe88e56d75b098a9587cf780cbeeda1a26d9a0c58f5a2ed663b68eda0d20856aaa4260b81e62efaee72a1261130fe7bbbd3cef656ccd6490d7595dd2f04e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e2614abe8e1d4bcba4962401b39be2969ee23365aca860f626300cfa5a8aa334a6947759f0bab9ac70303f2088060e024b1fb5142d1d60157635037bddaf317a30c1f7cc36285a8a56da0fcfd4a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b0247c9ec3c6a8494743bd51a48fc0da647ffaddeac033a0a33b08b14865e90234f9245d0a67853fcfe855b410dd05020504f70ef55e71ddf934bdb51e985d61ec613908a89e380bb83ebdde054;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h670056f9cecf5f39b78d19a61fa447059a586511863b236f83d5bab0498a5c183cbd854421c0720ad68a0924aa50a2790ba4e648c4a7c583fb9bfa87963952ca95b6c3c93721751a8ec2f1245d6a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea9236dc6a64cd527c5a970285cfad652aa29ad630a398259e596d582d6eb4103efa63f75d8d39d86865fa88d1c4e8646705305ff07e9b522334535f9e10df0313d95ecc3210ac40e7296cfadff;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a520eb85dd517c65a334348c3483d54ceef2d6cd0eff48c8d8d34bcc5ce6782bfc51e766344a80b40a79a7bdaeb1e5b284db971d50e342f4cd67ce113d62c0b970818e5922894fbb3c06cd5387a1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he29a5c8c42934fbe7ef9127dcf4e39d113c7129ca024532f501ca253d323952cae897bf1da6da1b6ed1dcd3bdcc2c6c461e7dd499c5d2dd9ccd5239950b2f710b368e809cf4f0c1f18f522132c1b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e2ea6c22563d8e86a1593b4c4ffbefa0e495b01ef7be6b171c38a68876210b937a78143deaf3b0760996bcf1c100316352e83fb71a4a7b2bf3a30249f0ee74b6695b72fcb1d3ce6324a2aa3b4e7c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf2425938443a2da913154fa2a8b42e4180a9bfd370883e66be6126b9e51b2e8ca7dafb71ad3c8df227a1d2d2f6761d3c91f8bc0bdba8d40b686a6fff3394c23840075013115a9efb4235ecd98737;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h777b105ad5483c7481ac9aca3620bec6911a607d18f1c8d565718a7c6efcb1b0d7171233e8268589a77d4254404590a4e2db732d78c49b6ca0c64c983878c30a2aebbe2a14a9be3b216870be309d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h495d9f27184b50e4bd756e33089b66e2fd2f12a89586df842854349bb638acb24787f66e33fb3573a0a2331dd2d5cc4428e8181335839264f916d82b71d3440a955c53a9ffe6dc135a41d8b5885d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e482f4fd0ccbf39ae4b32b4689eb2fa7c9d87be1b082999316c0b81e261a1e598f73d6e01621d38b157907f423d2043be4401b77b08c1ff99eb2cb30216e1b486e97320cb590e7d8dc511e7abb88;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f73894c874b60aca1a310e0b7bd2c115a8fd6ee4acd5c9e4fe43fc7612fd723548031cbd7fd910e23ef2bf690fb3e4954d35cf72257401711e869efdd816527fd30d47b160d9d4ef8e2faf7ea6bf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18ff3eb6ebfa4f2909a94a02ec1ec8464b18110a6f4e948ce9af8a04cced352b0f7ecc8e878ac100f0c926a451deb9261ce59db64b27746babac8001d65df08e2414da3cd1d7d8e39071a1ce93356;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2183a1c5591f9ff6c602415f0f8a6e503ee88eb0c6ed537fa377e525801bc9de3fb711907e3c17f195abfe98a7563742f2df165a475a8fe416733077aa2b3aa3139e83734c179b7eb4a2d3859a4;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92d1e9de41dd836b2442f5bc6d76c6f2cf25986df7965c056f16f51bd2ec012d2cf183183bd143abbcb7fce37bc45ff819628e191be58164936c7383c6de9c6b16a971a5f8e02ac80a37e324280e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f0f0a82a4961cd85eddb4527f6a8fdfeaaa17c2d8ea6656278cab42a8c995a4c992799b32b8b754789dd8c25748ceb80005d8e6d4683e0decfad9145b65ca97d900b1808ee5f0b17beed177d806a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6b4f01d18cfc221cdc824773fbe7b6faa3a1c53e4e68673ce49beca9d917392afb094ab2b4a81af2a3a51936faabf5f18ee25eb55e2793f3ac15e7f26432461dac3a047db19cc66e0649cbbbf548;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h103527b61583d178b7cd8a3a034fc3a10ea340cc52e2063ec72ec526852ad474887ee066e2fe84d2591324936abeac331dc036f2819d48042864e20159a2d9c307eae43c24f23db7f79deb98a61f2;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h146d16e176a65b30ddee4d811609d37a3acc32f5803589763475a8d8d1b5cdb9cc8d4e7a656c26b83ce85c5b7ae3d544d62e86ce4ef4b9a4ce2a9f37df86c9a416db2a3c3bdb08891552f2bc01070;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h860ce2482e770ba32a42cd5b4ba87aa764cfea472c9a4c511623fd2ad30f9409e727161154fdb8707f1036147903b39a5425c10829f4b2417830939564ae4973b011b7447143b916938030a86512;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1905be4b976437ff1fc80c36d222021e29bd04347ec6aefd2aad29816d07d37aba5fe1c315b06c2c9d178cc83cb00e635ca189dec437cbf705b16d90f5f1adfc4cb10c18e5e68e4ff8e828ee94b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h692201d6e889a1a89e03727f9b19f73da04e90af925206347584e268bd9eabfb2cdbed90c986f5c78806e795620560bafca12f8bc68629761bf40dcec8ceb10fbe468deeec28254f18c6b14a0d1a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fba392f16c30fb28b682e0e34f7849f85c2ae428cb3d9f717662b174037c52989e675178042217582f10d114a954d126c8ab86c2781f05dad11d270ceed4cc01c4ce2f23197427bea2d4594c8f34;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f83f498a1956db151d5a3e3f698889b818f5675a029c587124e679df69bce78a0f757c003c74cef647347828938650314fef18f3200e979a4c62245e77f85fb37c598bdf2167c406016c41d7be1;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67c5d1e9f5d3fa21a90cb8c183a0fedd4da8e98fd7d1ecf3e7f7396c9b83981ba846a3b9fbfc5a820ffd46fc38f0c11eeab179ccf06b711ee59e20f262ca21d2d8963687ea31a93eacacaf043092;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141efc3548a3a22401ef8ac33d8e5468df3606a481287ba99c5b652b60becadeb37a1ead8804f19b80e0645ee1b8e3f2c27d0154b5f85c903b200e3cb30c7b961e3566bd1009f9582e017fdd81e79;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1415f366c3e3eb48cfd879e916ab4525dfa57ea0aca19d11dc226060944981cbb8f2be4b434dea769350c0f9179ab49fc9ba3d2674c8fd0881a482dee9ab57f37bd923208491c8c2e2a03220d0125;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h250385df8d8ed782f081e8259673615ca4e142c9f87366567334689ea15e4b7a20e0ef335a9788ce47355f3b6fdfe9f9478e7ccafd54ebdc5291c34437226adec99d3d69345dfae9a51bc2e0bc8d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dc1210c62de2cb4ccaeb6dc6dec37022b68d4ca975e4cf3cb6835ce25b4e9a8750927574013c92203a051e7d1e6692834b982b306dde294d0cab17002bfdd6aae6c94e061829063132852a9fdaa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbbb63a9e30836435ca8b3785bf7f5f7a7f1925f2d0f0cfcfcfcd1a5ed3b2ad8260e3754bacf9f1e054118d7e17ad9d07b9f7f44488f1d382d9b5214182600801afc7ca657d05d379d86b4eb510d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169b526ed8592c7f3438e8f6ffcf6f1417e4cefe8b0724e05190d35ca97d97dac16d91ff7d7ca8f369a630d72a96900d54de2d1473ae6f50134d1bbb7217077b725fcd2e0a58f013e73641d57a82b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8683f53d656e42a486dcc7b2225ca243363436f50c59d8a4075960d4ccf5a6874c42cd9a9f7c6f10bc443b38b4dc81ef2264811c56882aee10a1d5e03b8f46269abdd75a0c9b944f924c42b987a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3b1539f0564ecc646f23496337b424a2180d9f598f05c166255ed4fba123c93fab7c77098123d13e22fdcb1c42def1319b0eae19b4fbd1b40f63d432dd3c75acc53d24a678ea2ef96a9b8edbaa;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161ac43e734454bf94db3065667491cb704c71703ff9db18f827800ca5a294fa71d0996d3066b7afa8e0f5722487aa71347ca0e7afbfb1ce7a9265913eb32fdcf00de792fc34b6570edbb5bccc966;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa48f8823f88b0d1cf1a3c6304325e6de05d4239eef8eb4eff3775b405420a1790f727fb42e6ca791c7397d1c2739816f02569bd0b8d028e4500ff7cb0e81c6ad9162e95bcc4fa376f94dff2aefb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b165c951ba66eda5643af3ef7e45848d18ef983e6b5fb3cc594e0876917b00c773d973a9500263546526e6894f5136455b0d8971ad72ba33f27c06b0d5fa4f1774d9daa5e64b1384b63f7bff20;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8fa203e572ff99456b231216d702221ae6d86e32eb6c20ae68eaa8a4df23a8fca931a42278dbefcb417773e35dc8fdcbfdc340a1b13f91b2ff21916d34f8bbf217cd2d8a6b8aeafbaca36434bcf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189cd5f0a9f44b2912fb1240f272ccbf0255faf00215a310b104775ff9eadd7e70b11ca9d0656fb6a49cb3fff72528dcef5ee655aae9c9438ade12e699162c510ecbed9765f0f38b2bb0d1d813547;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd8d643594676989f8920504df135c34d34a6064b99d461bbde7323ea3f2d68e2f2147187468ed4ffe7fea77c20ff19cc5698c5527755db4fd5da4f9c2aa28b0ae576cea4f28112e98af1359312b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he5acc218231f27f3db9eec9f18f092ca0b390a653383e89712540d8d00a1483bdf93a57d19f71fce97b9dc79cb0c5cc0774d4b5f0cc3a9502f61179a9ed3e0be35e09bcc0f7f21e79cf9bb27754a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h78b3fea46a8024af18c19d7f78e32aa081d1a277ecc1826d4c46d5f13c1886fb0938464b5db8edce8c882bfc6bc56abceda4a42ffa7bc5bf025785514e4b72fbe2b6e57da0e9c9267ea60996fd61;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e9a1f32a3d8aa54320fb2f01538a46a4249b373b70e98184e8a64bd4ecc8a02e54d8248abf709dcea40afc87027653f086427aa05c2a9bd67047ea65adcae2efded0f3debf1e1fd9606a26f6c12;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d595beb092ebf270e5569b2fbaca59d1574bd489f7480154f98f77361c6aa2e63c759abf47e1a4818ee7bb3998e4b003601594427fe053b0d3835c8941d07a4a8a21cadd48a62c929904d2e139f;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171437c73b45ae468a950a869f112a54d23e4acf20ac9b0571699f505a1a718a964326d43c41ffb04e0cd070e1f47cafa3d6e7ebfb11c374873c3f1011a5e5a066e2c5b3b0545bf6ed6d1ea1336c8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h998ce55589a530bc04a325fa1cd4d88ce8c1a27a722b5952255b8798d6123890b9f9ffb3d801fc793875052ad274d7ec2ac6a9e1eee596f34d129d0f21cea20eba3eed47c156bc0ee7978522c33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h197b7cc3a079ce4eb84b90ca12436ccc9309cbf8969226945aa962db122e501fdc535aa3e22409eefd38b5b0ee6f2f7d1c1d5fcbf4b2ce20bf44a61eb166783a5ced9b107cde0b0cf9e58769c612;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8fb24d6e58b9f56038dab2c107ec6b3e1e80021805f2f66a6a2656e2f5ae5761018e377955c82f72bbd2ded91c2b4726065e4176e91e65b8429ae88d2918b58e1316e12648597cd19298db567e81;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13781958dade01377235c3411c703476c6904cd56316f16cafbb1f2f55a42c06d2cf16af9e3fd4c23172119bca3adaf98a09304a172d74195166e1c284d3a2203752490d18543f7e98ef49191d6f0;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1612ba3e91da3ae0ad025dff25a638e2b1bef8e17da2136814dfae7cf9110ba1cf72c64803870300b57cfc7b0b80268330531103877e2c548ba3fca72a033288ab440971ba2718ee64f21c2762f6b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29e47453413f75f17b919124ea6a251a08a22c8f7fdbf57683bb3c0450ef1edec1f4db5afe811ce601488b7b91b6e2c5eb4f106515e4c99f2f968326b2868178cb2d92c32f092f339a8df6349794;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a7044aaa07a026e50ea3abfd3c206998d3720834b0c3022a8e71347ec6a8c440ac0ac935dd657d566837efe37164846e2651d096576e024f29a06472ead21bd1129340202a8e472222f11888eaf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1926acbd3d6840256924712d799cbf93189c199fef358b7bf0829f445b05b9f04ee770c943777419c71700206193335ffc35540e1ecd461b990518e424c3feb07a542e245e52ac8ea4bb6f524f2fb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7b893335988a50f799fbe6e2914cc86d043e8f641f9333030792bcc53b2e8b2606056c9ca23879f1cef4cb59b2faec052d6c91403d4cac9e23d781638b57798ec64376c4c915d52882d251c7d25;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4229bdf6a663910709cd17e18a7cabd3b610039904ac19f5e3b8fc7093a064f6861ff7938fdf1fe56561cb7fac474b04dff42dca6eb5946d7527777b500670af65648273386709f36e7b713dc7dc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d8abdeb95529e4e90993b3f845f1067441a4f34f15fc5d95cb06a3bf4357cb0fa36657c36b718a5f494ac4947d30ffdc6dddbaae7ef402c56ccb8662d28f82f56ae6472b3046f4107e6f81b5c68;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he20b7667cf8bc1df9105de1f017045abdd66ba379cdbd485229ebd0afc4006adf35b5d4d5131d11a89948a2ac57b5c196166a6711ebc3968b8d1ca5bc6e158dd7509eab8bf715da9f22bd6adad08;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f06c05134eb7e57e39c2e91dcec8509328a37ce57239605aedc25271c039ee3e5eb6026f05be80668ccbe62eddede7c3023385267fa75be8fe50d909f65a4c17bc982d19da3b5144a4b252e01e59;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he50a675e4726f6e1e69afdcfb7eca7ed9badd9b99fb7b3449e89466183c57c0b63b146c0a8a310919b048091d121f448a9ed5260682ce80f5755aace04078ebe488453385ec8364991f5b34b5d0b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1208fb92d697011e8c34b0be08d939e7c6c58315eddb9bebab9ec5ba7d81ab61e5f07a1827c407693625d1298f556ed1034d14ff9072ad59afc5feceea5cdad441f247604b975571ad1ff61cb90eb;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a92d55dc76c7b7d8d000539e8ac1994e73e398d13fd82ee394bc627d1a647d2390ac80311f829cc7d3c3d3017e25f36c4fbf6455964588f317fef1d99cb3db0ec5eed4e62fb03e22a23865a73d6c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a5a240d2ec19d1781d01ca35fd9fe9a4deb54f32048fb1cb4dc2831784426fc4fa96a5ef5c76cc5f30ee59b6cd36bc5e16c56522a53d0d4436cac2b89e8e06530288ea31648b193bea17210011c9;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac99c74940d2d226ba4f4998e5db62ca93280366edbb58191d320a5ceb2fe24f0d09d9626036c53d7056af9363429b743f595da3cf495577810742f6ba9a7138b3c6427d0b0f0a00b718ab1aba84;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b3057ce79b5c910a3dd8b3fb57c5a7235ac0f29a0c9d62f749b4404f72cfdabc813ec0b92074512a1336d9fea5a2677bfb91291750fc253d1cd7a342c3ab0dec21a60d7517965447245a926a92e;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e67422b909cac97841830a43349257e2970e21c27ec993ab6b231ead06c155bc2c70ab6872ae5f8f3e2367e47b23dfecdacb9fd54aa140e5ab24bfb0013c1859e041def8470b15dadccc397ba76;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1ec175ac423eda2d23a693a1f4bc6765847e457b59c1ffae5be9ebad671835629945af57f869a9ecaad3ea59ea8ab420daddbf3bf1b821d3056d25272a334d07992ff07f2eeb3e638510f802742;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1260cbc48b06176f195ecf1f7c697a1b78af7b0be5eb83b7d4e0ff5a8987414ce8d6fa9110c2cde480ed0c6e72633921fad27526f79193d7a7cdaf081c9543037e560431625d27306d91508a8dfe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0584e6de6494961681797a43b19a040029b506ae6d0828b8a34b900684d7c7d829db6dd69f19c88ff818b04a3e37d1c1c4932cc2f79fd6f33b08187481d6b10a57c21f4161a0737c22155021c6c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ea30182bc173ca7b936ff994a2111c4d39f33d435857bc1aae591279eb7465f66db0a1c8203e672c77ab8121fa9e96bd80d3519239040b3187c265ac230b1bda162e9a152181ca105415396c5c4b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7d6a22c1985876eade060121f5fc9cb6a33adbb7de354def8ff29f5e9a625b75818da3b665bb13df8ad86a0046a7f57538c10fdfd73f0c94fc048dc6a7bc2bd14a3d84e19c41c57ed71347ae2f9c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4c59bd8effb36d6676482e288aa12203ba301dfa850517cf2d96e226564a7d2611b01c8c1935cd760c4c7d8e2a38f9336e4164ce34093f750c4ff2681913a76f3f07cdaa39548f55d34a01713e33;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcdfa6768d0e498e44d7e5fe36bd3df3cc4c36ef5d82d41ea4252547b1b60c4c2eb0dd312cf21ba1fde248ba07ccc898045f3c03f593c6924226f766e62d38f0ea32008d3cabf22e51b7ad589b1e6;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haba720f17cc134d10f643ab61def18b799ecf52920e369570fdf6d0348e03c08e1555b2682f58060083e15b2b31c2ccc44e4e03e429ed755764730b0bd41f3f6b574d8910c7837d20a56c3f791c;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1604dd4ffe48b02d6b778f1cc49b44b15ea14e97c27aa2d544a05c30db83633af2a74713817eb5d9f28bea99a72f5cba241255d68f31b182b6293432a1f2de8e41d8ddc2673f927aa84c29e23cc15;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17dc0ac05df0df389b42e8c345f47807dd41d139997977c8988ffcd76424da0b2b46c87c34e70f9f6e5f2a57f7d6d94c31af8a62d691da2f28c62e986c3b5fa7888d94248c0e5397efd9a77bb40be;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1584cf027f21ccdbb28a8ed8628668b58f8fb340157ce9723808a3885d33b6b5857c48be1e13c9300aac01f6edf0bb0d929942201c5d9432f55ae810cc5cbe1fa22b757a7a82bd1cad54f14a7341;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h104692398c08b85362a88646339311ca3ba4087265ca41b67dabb097fa33295cf90a5d0009a193a86bdf034ac250f7554d7301dbb2417266af92d785a4fe645f818efd6979c1c716457a91055489b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8dcca18effc453cff7a07de85e703c96d0b75ff5a9c6fb0c1ff94bdeffc3f30bbea75f2a35e482f0237a5ed70a2f195f429272ffd2b08741596892e25e5ae8a43193dd0d484f4de1c585d64e658b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15af84aac72ec6bfc31e5394dbf08ec5f2b700ea8ce95630302c60184a201df06515d08dc90785022c35045237601de59c8602f175f3f9bde20bcb5ca038f467606a254031b9d519b2c90850c7d06;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f8d0800f8f10b70f79ea998c036e6c53de9697409d138e4ac3308313a7925842154e8caed5ba154e20eff3d3ba7ce2cfe0e4e1eca258b11b6f74146e5e5e46c0753ab9ed32929d08c74de1a80fe;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4e80626d7c17cded381bbf755d015e0f13a699fdeb67b65e44dee2ca6fb98fcec8e2bcc175c6d33e32988d094677d8f1eeca8da78f90f90d3800023e1486799aa583fde4fc067895260c485b4e5;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h983cdcd3e4b06184faa3eee2b272d0534e546c247dcb9a7ebd068bff9972c56a1446d1485a02766abcf0f74d12d6e6959f465723a21a9ee728b8e8ce2a4dac7982326e6cb3f5deedf1b92337f5b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc15ef56c36631d604b5e0205acee6ff5749c5edc9dfc7655cfe0f80f71c4c666703e80c39793923b3bb5a7f74301a03851c7e6176cda1db264b0060790b5a4f2b320293863a885ae867549d8abfc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c3f996d5a9dd85ad20f551aab9c62e97e35a102c7069137e8c9fa4c43aa2fab671e629aea1c81ac0bedc0072113ef31093c1f27947210edc2320bf0970d21ff49247d74c442d01e960c63187e2d;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4484fc4ca2ff462c528e49e32edc4d22304ee233cddc9d4d47d1be1345e4a678844a7946b0ceeee9008c16180784e82d1e04fb38e1e01027c1ba042e078cb055b1acf1d204ee5ed7e7c5bec1378;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3354b5a46fe00874873d941d7163d1237541696691b23940e5258dfe15cee4533a42e6250b7aad9aeb3d56acf7b3b11221fa36aa31f629d4aec51d9fcfa7ab1bfd2109fc3ca88bfd8b086279533;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1327318b508d39e81c8e878ca4de090c3af5416d3f3934e038814aa6e4d8d53a16b98897ce006cc7ed2eb6e33872d2a308dfa42b2e3b02a7d409fb2d3d1710b5c35982d2f2aa8b5b00f26dd7ec784;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8023a86815fe8b03342746b83229b1da9a0d5b7d7ba58ea15fae6a868d780c788a03eab1e9717fb3e810ca1b620dc81e57e493bbb71e607d15d8daedf11c53191884e1fb9a167dc9cd82b8eb9d7;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd390d724a2c39c45195954fe94a00a14e20156981cda22c8554c01707c1817cd1e8421c97b40aaf8075387e44cfb1bd0c781a455eb326b8239999323b67cdf9b8450f3742e253aaa7ce50830d40;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f1afc5be12743ce48cd7765989d528a3425097a56fe9e6cef53f7a6de4d2d44de3839652adf28709c76e3df5e49b4dcd3a8a0aa671783759681192ffd6b5fe9c1270773e9ab89f620a0a8fa9ccf;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191e2ce09d1e34d7ff2d4a68bee705b87df7d873364363db573ce3a276bb3b6a30819dc2109dd1b78446c6b2680a61bd46a2c881278026a04c794f5ea024bb443ef438d642af770ab387ba46b66f8;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6737e998f17b012595525f2ee13a9219a90597a39a060cc9150d6320e1bc64ef48cd87974fc4a263f082c45c33491e67c51f1ebed14190b4b01bd6e901d3f750d445b0a809aa88d5fe01bf87525b;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb03ce8095dd135d8cd61aa79dea36614bcb39e2cead08be2f0af2333b4f026315b1cfa2e5c3456705e1b0bc01dad35956cacfb49c8bbad5d6eaa4abe870e79f0f704929299dd56943cb3b1448d77;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h193666fa0a9c03420bc9923f4e7f864c28f52b2dc42b3db05d9a60bcc0972f1659d140f881acbfb469ed1f0372885cb2004664e42835bed4a78df74bbe4698ee399660c4653ccc33b0c75278b6929;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7cb108334b9d49d60a8313d836c65987c7c2084b993ca8fb40d051e290736322f44c5902e5a3f4ea12e186f83ddea7bc6fd4c70766506fe6935a5be631b191b55b8a7f7ea52adc0f9c4857093181;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he50a610eab13a71f74b584adcf2336894a62e2be4a49f7ab0bcf5d114304a8cc060c46ce7ac49064494cbdd51d338e02b9a838d5855c099181fbd99f4d71a6be8bd4c7942c3e96fce1add178451a;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47b8af7afed81f95f2bb97ad3c64d498afb56f0e11bafb9e2dcd1690b1ec52ba31db05b2167c996f7dd792c4e04e73a7815981896c922417f0f458f0fd603c496db13d9bd0ce204e084004e2a682;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b07451795eb60c50db4eb36743ceb49f5f4bf6662f183b54caaf0fb66d448b3ece6f50561fbd6789797d9d6b8e1ed069e04c881f18fbadea69692d36381efbbc00927ded2025ce37c0dd2ef5777;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce7da5ffeffc1065ee5a735e7b951a8095bd9b5a9b028c54334a13ef3335b174191391d0ee9b7511c8844d65eca6b2e08f82059f85525c5a43b2057b80f480cd44ee9fd7a5195e241864729944cc;
        #1
        {src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f561306ce345816ce9fa1e1b01c1588d95d25d2754786982f64b3b21a5fa19c4837e66f072dec8aeacba80834e0dfc2a487fe21514aa09b71d4d5a4b4df0e3943eaab4eff916627cc46ce4e6134;
        #1
        $finish();
    end
endmodule
