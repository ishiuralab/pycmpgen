module testbench();
    reg [21:0] src0;
    reg [21:0] src1;
    reg [21:0] src2;
    reg [21:0] src3;
    reg [21:0] src4;
    reg [21:0] src5;
    reg [21:0] src6;
    reg [21:0] src7;
    reg [21:0] src8;
    reg [21:0] src9;
    reg [21:0] src10;
    reg [21:0] src11;
    reg [21:0] src12;
    reg [21:0] src13;
    reg [21:0] src14;
    reg [21:0] src15;
    reg [21:0] src16;
    reg [21:0] src17;
    reg [21:0] src18;
    reg [21:0] src19;
    reg [21:0] src20;
    reg [21:0] src21;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [26:0] srcsum;
    wire [26:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2746767e8f71e3940ae245f805d56115a98783f4e8090d35ff5d790da83defd96713b5995293be3750acd586eb97197b8b7ab1656d98f009ececc84b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3871d6a1284d5f3adca4394d898aed146f87bcb533cda85a678bedccedc6206f5136107f374b4032b7cec143b33d6c073ef0a447b9c1ba21c7b7c5d31;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda2667d06258986ced574f1c6882daaf8219477e8176161cb45582e16da357005abf10a5c994596c9a6aae6e1b179693b9632f98b507241e771fff369;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e5a39251c814786eebf906ebb2f87777c1d717db4b3059123e35c68269c0e4f3cb593b788bebed2187c7e147f06b6a7846f9ac8d0f0e2f0390517147;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56b5c70462a05c171dd95e83c0f98378d29172a881c81fde75c57911b421dcfbf097cd685c92da8a443587b0e3843925aed421fe9b7aae29dbe1dfbd5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde6063e00483f76fdc57e8e36ce35cb7ef5312367711ef079c631407f17a52543495299cac93bf31dc6ca78a1d8358e2b914c76695120736ba584aca4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ee20f10718f55630926d9a9f993c7d20dc850985177ade28f9bdefbc52f3a1237116b6db1e862f7d7f322313e4be86d6a501d3bd87fa5b9d67f356e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5be77bcb13f08c1c03da0e201a634d255529c607de5427f6ce511acbe900bf365430404ae24e94f54835e5d821fa806db275ae0bc40e655ff3e8574d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5db2f1e1b709f0916e06ff0637e6d1c8cfaf762444193262c62b6dce133b95fc71b2da8e4a179910164ffa5bebf404d4f096f8e398a35d7c35fb86176;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f909f83bbd6d1ffde8344d25bbcbd6e7d6af3539ebf8f5d2044e441fae997d31438318b11edffc6c3e33a2b18f168e3e7bf333c7a5ba91bb72a58c23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0e3e8a581f848f94cdb3d1c1af93b87d2fea5779042ec5212c1f282d8ca5b30a705c86f0140b33c80e6b6729a85ef76d86f8c286053449538c1f8f4b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h997186e46df8f451757913785d264c214fe1bf3e3624bced0a4b9141111ecb1a51dab47dfd6573b73c2508590d016622cabd72c5f2d9550fefce1b455;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h409b249567570ef0c904c67c05894df32aced7d4a44b36c270d0b619678bb865d90b15e3bc8baeaa60fcbd01bae7bf1bf4f48b254709d80eea407fd1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h654525183b17c90bb97c00de0bd4391a541774f97e9cdfb2249518c4aaf79d946c477f2097973dbbec083b376db76f50742e0d0f92dd3fbdca0bdb3cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8988ecff1462f4b963d891026ad22d42fdec17ceea39e09df1ddcd3f555ce31ff38cb971e2c3b7ad713edd98ff61c224059834e07cc949a1ef2269716;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff63d95b8bfbbba0880e8a655f84396966b9a39f8f0501c4b6cf955e498fd3b4b448afffe36b42012787dcee65b51b363a1b9a12c93ab3f5a912c8697;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6df436c33ec0d3c2dc0da8dae001eeeafe0ba556e678ee498f25786c7007f28fc67328f141d8706e5ed3e872672d636faf2081a620c7820b3fa03890d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd05fa05f7e59e85c943b053a3e5f3bb5bcc48338ed2ad226d6af11bf32e1424d86385aae97c5250bd5072e1efe2fbd8a3d5eab35a056aedce65ea4ec0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb646e479a4f58004d0664aeba45883ba45e7e6f5980fc15a45cfcb39a2babd0f57ed0d1c4e79c2663d33880940be9ab526d8a2539df23757c8d95f2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e4b5e72ed3b0fe808957d3a76b1aa8eaeefab0b449e61d0aa81db9cf6373deaf1c199b93d42fe11c369e51468a609b7f21fcd318d45b52d09c038030;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4dacb2e4eab2c54bfdba2d2ab2fa0a0908398a06171fef12d72fb9526dcdb3b626fb4f1fad0891c4174cbaa42a4f4a6092e5a8ae62a28185bbd9c262;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc729424920194b1371cd698b5bbecf1b69dc95c5811fc002570b796b647f8582458d0bc6ff6becb40dd9efa9df40bb45e04733ef0f7f5a0b7102eda18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11520bf0ffa0cde2400a8e277b62213cc193e023f91a31f64b05209228edf3e02f423f3eb0b9e75e86ae64aed7cbba878c31f2fa17c3a8ba08b3e9c90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h916bf5ab0b606c563754e33093bc4c5963df77c1c4b9a2254388704d120dcc006dae630ac71946f3af0dff87a89bc95f87d47446bea50a4a4da2af66d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14e7e7c3b1364b47c9bec8d4b41332bbcdae3792265b48b8d8e1c488dab0bd9f8293b79dba61c1832bdffe7b9cf13edd5ccf3fbb78c88f95a63882872;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3b69d8908649e39b695bbc4172f6a9c58a953fc7e5cf48ed6771078301386f031e6e582deff26ab7932a17f4e0322a4c19be56b2a5ab57d8c45d7704;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h433ae2475e05655922bb04836cb3401e0343ef5c948175340e76f40676da79cf0e1c4308eb12c16d86db8576662bac78addf332a52483a5da0a815917;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf9e3eaf478e9522b0286a039cbeb04321976e66113f366bc4cbd03b896abd75fdee767f08793014cd8dd8e4bc84bbf50c47ac6de0b2ed17e1c0b8992;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h352d0363639b63d3cf4bf9fd4eb37bf67d9e2a80690d0aa4aa20527f3ff14f5860dd47762a9aaede77454af7364c9bccbc5005c25dae8c9c752ea44ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88c91e16a0de62944294098be06df25cdc175c29a967ca860307c1be6483791d7858741ad52de458db16636f6638e34f89644a1f77150fd84c88cb70a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he957fc0c9a0f83bb4aff04b2aa283e0b804a0ecc30176ab3392e17a6935067085191056ff65bac565013a015956881078902936964f8a4dad02c2c0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79edd3519a9556b255c0bb0d18276931934f15cdb2bce0ac1a149dcdcd677f8ecfc4c36d12b4a1d4e2cd0851b8b83664c28f3b53d74c8df0e6ad8534f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d664cc79915112f51b6f675a6bc06c3969687d24fc40e67736d650028ad415a7a317b03d712fea6b7517e8cffbb430c18a542246863b301c772fc128;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda7c1f28e2347230bf235dc7b11beedaaba4d3405d22fc834c930804fc0e69b6c79c66fef74edc8b7fd515d80e71af18e32a2180e0e76d6c7bf8152e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48f29128889e7320333ee88b1bd9b487c670e5330a6d6e484a8a8b20450a01f17b19951396266e6a31d52ae38413fccc38645c7f8c3dd5c2ff187d0ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8aa578c91522cd8a069cda2ef81614ef480ba96e3af909c5e33c4a0ea8f862451ddbf4d9870860d615f17e49742700572a4422e2812e33eaf2f602cb4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78b2109cf262840b979cce7da40039a5c9b1c0457aac57be8a71a81e1387d4d1e94d4e2223ae2bad9967bb577b6908e84af0c91857d29559f5d44dd43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb95dd827c4e19e6fca5d422194427402f4a2c36c5e44f1bf3a89ea88e5716e9da50e375684b52c265386491f32e573b4440f4cb87e0b206d1c8ffde7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf10f16511f52209e3e8dd4085851f01a28a302449d9270345eba52938236a071d1767765d0cb07f2b34c7aef977b398d43af60b84c7b300d4f664ce61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac78f69a2f147692953287bb9c971fb63a3dd689277da785727f530e094ff52cea6189d69cc99f21cf695c7b94657fdcbcd9470dbd50fe04928cf0f25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had000eb5f5387241814fb2e2fa588282b23812199650484c7ac0fea9b6230a6814bd7d80295ebbf811a4689af47d4a1e214aefdc3355e7bc355c8a489;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f276a470e417a2b7044882e1254ae981793b3e3bfcc9ef626a66752b7e402c5a2dcf7124d3bcf8428ddbc1f887ccc11d4b09fa4ce9cfe59bca16aad8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee45cac0e1c25a0c3058d45a30190b45d2289c4c0251662ff410934611f99e3f1f69ded6b99105f25d93470996a26cad7d68e7df9aeb32c6c1c0532ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfe0b1727c1a532441f44b161b98fe2806756ea54e5440d6a7281a12f8551023708b259fdea3e91fa0d8322fe3a4e8a1a063792e6e807bacf91dd0ddf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3a3446efa4430fce6e25c2b6964a3c93ef7bab9853b172541adab6c8227b39e8709ba17972256ff9bab006490b9f1f491200796ead3f0e561b49170d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2727abb86b3b97906703a897b2d2d3f4f44dd32c36676819ddedef45320c0f075fca27d740dee984ad984fc40ccff061e81a4172677e5a51eef46ab2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d38c3c74e3a9205ce9dcd0f2cc24323595243edb150b825676f683ed2ec18019478b2679e92bdb1d893198184f915152ae4f83617c4544b5f3d08371;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12a28e6b94530b6c3330780b34f971e2206eb516354bc1ae84ab7d3f91b33a4767b54604b444bb6cb3306d7f09c13bd1db15a19491877385107427956;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7538f9d77b92d692ddfa2b6e90f8af082d8b2ad142bddeca13a36aee1599cbb1e4644eaab6e6011117d5b3f793e8f33cc5879a3600a42e48215301d9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfe3c147aad0653481191db718936253fac4df4ca9ae13d568bf437200e2aa91d381dbe4c155ff25a456635b60fe45560cb25f351ca8029435681b682;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb81a8ff4c1f7ed276deaddb8514dccc92bd66593c51228aa29871ce404f64c845bf7cb02ffdc5461734aab21389d9a66a738967d6b5758f982639be2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0cc5c497f6cac23b0537a86fbceffab7b3d21ecdc592f5813992b89038e2ee3e3f9198e0a254ce71dbceecd514b913a1c85a9d015b151f97ee66a3e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6941ed9bc486c024b2a432100604fd683a01f07df8de84f69a17272256227ab72d9618f4a1440507836fa09b1ac62c9d9c609929c2347c9e6c6d296c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec048276dc45b294834a1b2b46527ac313f7db5f51b252871afcb8cf59f22016cda619d4114ba7e6a16da8965cc0380491e094583f1702d10d1bcca1e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc06d8117a2088218b17d6f10037b0dfcbde9fe27ed98c71bb3382dfe651e1a74b0807347c9c05dcfc51769842adf2923683299be40eb691ef89985752;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62faae8db313add935a8fa22cc5416857c75790db0752246822951f36f202b7bc16e42306f672d92e9617a1fd740d920379759db2e18ddbe7547c83e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36781ea09d916e1a883024f1be0b8c27fb66ea9c125e7504aff23677405540105eaa8ec3621f5a5465064917c16708e36dd203352811da2abb1600e26;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd91597a3b2bcc5bda586f3b2f8d7c35d50067b3be662d8b876d7173df46d88b231ba3cbb81e2766501d2137436b308516926a59cfa6d6b0423dfbb05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3d628453751d8f01c15bd98d7916cad07d740cff95c47154d3e620690c77bb29f19a756bc542a9360cd5f7fabb19d2f99a1d6b22ba4df5bb8ee971a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb723f470610abefc5a2ebfecaef05c9a52fc462c5e2a8bd8c60462573173802406ae75a15784069c506061710549d2cb39ef6e62015fdca518da22aae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccb5a4f612596ce7be5a91cfe343c834e81ddf8a68a8c549a22dc342cff63c27e73368cc7e0da1b85dfde53df67e64a273251b8963c93f1d40c6aa64a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h983942b615a8dedb6d95107a040fb841160820806faa6232c2768ab7a0735e24ac4c48af90af9b5bf3734db7f50b0a23b5a141e507cbb83a3678eecf9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27ffcf21c4dfe301e56a6687531d0d1c20965348e195d50a9a7565e50e5ed4e9db7dcef834373514e45c7912c0eefb5e316ce8d16badea9bae777ccae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h514aed55eab59331c174f5058c8b9c0aebd5d2e2bf6e394a227edead08f4310e567e3d080cdd14ca4142b150c3a0cfa422fca9e38a3b54aff5f554f78;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8d90353ebe4dff509e32c320e4897417af6c12eb6602b24dce106ee41844dc7345d932e8872ae51646af4ed35ddd804bb7a34993d29168011e25097f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5806a8019525f0ac7bceb758c4b6864cd496c8e009f091ae1cb74f2dde7daff70a1c39d8c4678b8d6f5efcdee0fad29966f0f3b94ffdf37b615dfca2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1dd4149ee84755d7ba0a2b7d21648b516ba4f93826e06247a223aab646a0b09ba4770bce1a69933924217327c24e17ebab5e64b96dc5728accd6d3056;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb94ed4cb3fdda8e9adb61d16e969e728e7648dfa5b4a4423420fd8cdce88ea5a79b40ba3b96481c5acfa1aa6140f25cf1a59b6eeed952d9b38c22a85a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha084e06e8ab7f3cc73329dbe6f7fb9f4ef609c9082fb4d417202e38d89d7df1cd4e3f5943626a75e43ee79ca21e3b238de5881f55be9d75a63c387463;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h412f36a4555eb2be68a472a1068eeb12dd0694d117b2fe58790645b39ae2a972dbe5464745a464fc7063de8718af217115808d74d59d4a545a41dbf87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbf761a9de91bc20afbe62dce0fd0b33e0a342c3c54d3b27f97a32f4f9349bed609c99c2f7de6398c1eabe0ba7cab95f77b29c0ebefb9105d445b4f28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5989f290a9e4f94f0a5fdbd36d8fe2207f6b26c0843ac06292b72b532326ce0d0b7c21e060e42ed6914b213fbf5315729757f140277eb2a8d9202382a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55c7b1700410a7027f45ac5b8f76a1cc285834a02d51e0da56ce6ce2ab127711b1933351f978ab2652dc52a76bf411315d8229b30a8d2dc96752cc3c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31ea3d1f884b5a82a88c001df041fde0a173cd662e19612d515a55f6dee7afc28d66ed12c524690186696ff260eb9abc0d28662165fe429d9116bb7d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd52aafb6ad682377ea3d71903e690080a7ef7a782e44f0299923ae79f81894861b940192c372c6e2615bd601920088116252149a8a73b515febbbe711;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h989f0e2479cc7b15283b787321c622853827f1dd0f094d6ce45b96d3927360b3bf27a8f8c41705b8da9765c0106744501718e43df6632bd55ab325c96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b54bfbdd669ea4778fcef114702611add0263ca4d6423f1df38a8c6c32b13d549bd0aaa09fcfdf731e39585a894c10dbad81213eaace451b24bbe6c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a78f9f691b197279adae3d3f8872e4b4987a7a8f0c7bff7e82888a5129f1ec4fd65083a6df85f37983e80876986bfb97fca26db0a11b59d44a75386c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb82f1ff7862b8b4bcdf5810e570a1419d522102ff63a688c1297d067b53f18812aeaecc15779dcb0fb1b35ea038afb87a9c9d1aaba9621d9c01b7f57d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd67922a30a96cde1db167b84a3b6068b4599078b5801b1fdd8a560bec05571505a848b595c8bb681aca237821be929f0147def8733c0d74a54f9f02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56e0e6976265312b8f91dffe4072cfffed792bc7753b74b80e34f31e162a42207b733dae713bb362e3be2e49ab8e4363f625a938764c307e6e0ae5efb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71c7bb828110246eb70656637a882ee667788f09c3e9caa7e8a0a6950504074be6d30b089b194438a92724bc7d706fc9b6dab0a18354577d96923a1ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bd4a9f0bd160dcf85b91f45aed7d2a1757299049db3c7f9c5711eac74fef469e7c71e4bf1b6ad6c1b1e194d5593c0d62d94bf20a7ab1deaebdecbc98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7be30a748f2f8b789675ea4e322ec2062b16f5d18c1b6ba46bab27a3a4a251dc7e35e91da97e8f9d6e38fd9eb3c656d7d56864d7e00130b81f8027703;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6bf589992c2dadef635c974d9591efb395826f928fbf6aab98ace229454b01ea52633603c196f7ab736b925e98183f327458aae7a7886cf12811fe5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ad2bd36e372e832e7382b67c79e57f2fc3363c00eb949714f132e45ed77bb5cdd02864682fc82038e7e5520e9d32f1f837f33524fe28e088f6d5fa17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65553803913418f71ed13e85ec68f0d2509f98d68ea8872bbf1aa0538d053daa2ec8f4abda10593164ed630af2e38d941d82987a95b2d4b6fb16e0bde;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ad635fe41ca050d9880d908d40281dcd2b3fed80f40dca42013e93df1158a443670a9239795bfe86e31b5bfddb82b3d5e2d84be7a65b59751dab1610;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcd55d72f243568e2a61e7b7e1943e68aa803e1bd92b4ad048be216b1c589893cd1685c2de4e44ef650ee49b3e0d699a776ac5786ac4ac8668540e0b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d908edf8cd77d6995dd18a8b3b1f54f8d7bc5be6d9f9cc70e9ffe35ee29239e408aca77e3127e1c5de26935b4d2362c64103beadcd623459fb540b8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3c7e8bdeb3ea4cb7e4e2a38c46eec2f6ae9816c734b0b370a0becc31ec3353fe59a5748545d3e0978969c493b81e18d72d1141fd52af3c1324be1a4b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a491ebc71f5d4ac5859489876ab23bd5f1e588df48781413a0d4c7f7f4456314c79ebc12e56a1d5cd8271bac15921e018e52305fdfd647bad6e955ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc68c02c159ac05f52cbaf2b6921c83e9a68192374a1d425f94a56b7e398fa0c67a321d4c5811a4c165d6a8782349cfaba3d448a948d00922a9eb1a3c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6aa75cb795bb3595e5da362a20ece18dfa477984ba27b14b32e72c48493bee79ca3f1f3cdb47cd8b9d5b87702c4a7813f1bb7f80cafa56c53ed85204d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb9e910c46086aeb27db3081606c50c3ce10ace493e5c67b712a90c00c458cd1b2890a02db8e7a31a44aa42b9b6802941dfbc957ab44295a086ce82f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14322f16c474e092047a9c2d6b6e39df370766b815d31c3784bf27e9d7d98e3d50f9f238d042a931ff3ccd62e5a54fbcf69803feadb6f4db5edb8ebef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5233bbd342d66d6636b56afe1f468fb94279fc779fa2567b965acbca48152fd798cd140d058d55dc5a1f4230a7d76d167191f517d41d2f6781ff5d47f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h367709fca3677ccdcf435812021dcaf42fc4a3d8ab0ba544dc668b3b635e5f16a7435b49cb054caed484efe1c51c55c966bac48d2584b4b3e563727af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb451903108f33fcc1504e077646e1f26221fba94566056138efab8d3da36668443f089439c34a05dde8f1fd89c2663a24b9d7915939fe311f046230d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f9f8d341a309abab8ec0b68219a11d585400e921d1ef56135bc6f607e781b0f1804e279cef3779d73d8dd0c589b931af9eed2ef11757f361e1dce890;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31e4cd0d070a1d0bb80d5fb08beada3e59b67efdebb32c6e156dfdb0c47c964dbe5bfd36cf9b851538be70debac63793c47affb65519357cb4d364538;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haec68e7b49f8717d05e496b7ebe3604a63e81c4c333ff79c2ec52b24e67e547704a5ba3ff5b9a0ce714a83ce74fd295293deaa411e05bd33070380558;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24decf7b856e9a00bb5e092fe45381c6ff004cccf93db5affd9746c135fea8eb85562b831a11827e11f71cd42d710fb6edf579edcf288c034c7d647f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdb1f3dba7fee95269bedb9f655670fb1defc332636eb07c3841edf535165b371d721a7f6beabbb95d44e6dca64fc8136b3ebcb708748e3c14a70a66f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1df4b3a37d846261a89841da4fedca9b0d19822e801b64972294fb05f975fe0ae737fb8306102b1f768aa3cb71188a87eeaed009b564cc80a97c60af2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had216486bd8bd8f1fec09770d1451db0774fc7dbc8010dff77bd2e1d920a2a38d43256016f32ad9d692aed832cb377c63462a8733a3e5e4d76ad247d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a2e834398d4786c661037566560084aff5eb7b9885e5bbb24e7404bfcf8f040031c117b3316e5eb3282684ffa960a0084506467056d3b91b98acf5ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d03b0381b28d1a68747e865ed13b265b82b1a4f038f4897375ed3bcb7e179d2e02806c8c3c5837da6cc42e43ef51f34b20e20f5c84d8031e3109b9c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h230db3932961e4a7c997c0649b1b341154a85d48e69be01f9391b299b769a1d4d9b160b2137851ca2517594d439cb7469f041b7db2ae52db38cd0a6b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he23707faa04b027f99ee564eb04b90782e1622e424b629a0932b45e7017eeb4751e14cbc20965b02004e534bd40ccb11adb182ef5b540ded770e4d78;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91e8aa51bf89217701c1b24184413592aaf1ef8515d7c902d62d989bb8ff1f2cfaeea24b59fe9f816720139f5557f4ac9e00e758e722edd6ed4dd257c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d5354ad2d0682c5877ed65f6554eac248e7548e090450ec21258ba7513890fae8cd7b00994146ae126cd86948deb8814a7564173fec6eaf65bf50b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca945fb617b302193f74a57486fee3f482fe04afb87bee8ce2ae45eaa91e8a28dbb7ba879f2f6650b887b450a1d8e763039ed0f0092da2775369df7b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b71668ec08f9c255ca598d224ab2d6889148f8110fddfdac0b37d4343c1aff17f6f64812722e1bbae517ae586de29a86c2991171239d12394e206e61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf9ad0744ec9cdd3cec54c940e0a7dc9278e13d8c80872a635bec91f6e9df04f240e614d6e9feacd223322a880b5beb5f26081a2f80ee9c6c85ca8f55;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd1f815990f166900c3f783094c9b8e0375b772f267906ae3f023afa1c4e59b54d8d75530ffdffd87b4643b95a321b64760c05c9bd5cf8efc472b506a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf75efa97b6071d8ecdf38c83df23c793a7a204c930ad0ebace49d695fb75cc59291814067047ae1df1d3ad3b8cf06530615e62da48e6fd04110b7e7f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a80d1e8a3142dc43726c32e14b963ebad48eb72620f46092e73ef8a1434d8f034939d902409992469be8c820d26fc6f70c6521ca73f263bfe6b09c40;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18abf4069d27df57f8d9c814add6746e4c3f04902c1aeb4f5a16e314501db02593e88a6baf56b3e97cf73fe8a3b5ec7a91afbc3e07a49bb1d3d1577af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h355fdbca147120c441b57ed1aed4a790f1eb8c24c5dc84e2dcd1190d58a2f4a058181df3ef857e4d6136960b2ac58bd0e7cbd988f520bffd0b46dd12c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7da6c645e0c7a51a0f2f672f2419fbd393440b03d281454c4521244c7a0ce4b60490694c6576158c6af0797f7212b0a3690b89baa39cba9b730d039a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1141c108c50c446772de79376c75d254766bf47543068bf66bc2acb73d3b763fc44fc3cceae62419feb576bffa212d5389a5e6160cec0c6a77f056e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h787fa8b6033b9bcc3d9636d9a7c5517576ef2db125bf58a768cc3a00ffd60f5d2462a11f9a729739f66166e58eedb6c18edbbb80f16d9a989f4acf1bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce59b923b451cb3c593257261c9509bddc88bbf51db37e486bf28370688e1c43ad9bdbb4296a5672593d2906a66c2c33e34c873ac955aec8b1fce4196;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15b766b77bc4ed2369a6749b198c22c934fd2cb16a327f9e18bd4c8f4eee4a2f29b7ac7b86adc846460f741e25eddc2afb3e40add6562da4d5c7dd6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ac8c51301f78343242657deea9db3543421e9441bd34ff20d559a2b724acabbd6d3dc7c608a7804afdeb61069003af923e9be05df8391e10005ac19f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81cf744d9ca103c53b11e56a6543726d9e8346e6e2689d6d21df2c51a302de7248b938b6a3e89d1f2aa0ab12d1a09c3c556da54539a7b1d73c303e9de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8aa2aadbd637eea96072d4fc59789c9f66609ce0abbad7361efe4093e994dd37670784b25f4b25d6e98833670fdcc908dd0c49d12325e707945158545;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3f675d4938a1967646fa72c84e221b7a9d96bf0081244080e1e4942b8e0da0e30d761858a8f21231e92c5d2892c57e5d2e91e2fdb7a55559e21aa790;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ce6edfc2f07076372a1d27c8b148afff1faf5696cb9a2aeb34e02f1e32609b88d67ab9ce2c982a07e44fa1de29e5bbcf238e9e4d452e5be860f7a144;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1cdf2a430c83488a941cfe7b466a420650af9178ec3aa25a6332e8d6ec85c1289dca435ddb388eb9d522772607f31a8eabfd4931ce352c7a35960bad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1684fb3059c4af77d3e6e49339ce0ebfb42ac8e77976871f5f9e8b686978738b983567e02abf1e76c9e32adee784c62c5aa32d2325e243aceb6a8d063;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1a9f0af725352cffbf469acec02e36e932a92c557c23f6c70dfcd1ffbe3cbae9e22f763eb5397371ab708523d53ccf925281b9a48a26a4e7c66a861e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9effb3b75e0c172c93e5c41902c598cbc71f6435ca389556cb84ba81be1c4e5105b9783c88cc32832b96ca46806b7e536c0d810b9f5023df7f2e0459;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccd6dfc288e0a247acc308b30d740fe11bde5c70b362f9d2616ed2312662b89d5a8f3f9d1d38c7be4d7b1f7cd8abbc63fa4f3b3678088cfd83c0c4463;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab4af1102c2676eade7a6fd9cc4bde579e843c29a80b174f883ce315ece1d1f76caff1322c998e2426b1ce50d18303dc74ea63901102ec8f04f4ba4fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb96af9b315361b1253003431cee05b901ab75bafa813e95a50ab399fae89975462c3dfa763d0409ec7407453f32a2137296139e8182c86fa0247904fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b1baef4b8273383961c95403230f0b0975646165df1fa76738305685efd91c24f702f8372d85e48ad81871b35b5aacfae0e0f5224cd258e4ca60a7db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5b2fb62186b2de3b1be1299153616e53ce117a0aa6707697bc0b5d80ab2677d31a6b5aec4fd4145e4ec310ef9cd9dad1687a8a60c7fad5668deeb706;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93c2cec2e2420e4f7283550f72c00c7d312fa1fda1c1095ff8f56526e9883908351f72c1a7879de5d0b151ad2c7ccabfe44557c47214d6b3b97798542;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2fedd973529d45e8d9be06fa87311f3c597ebd7806356324e571e67de6846f94d20ec65b13a2eded93bbdb733cbcbe15044fdbfdf358eeeb431432c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62b8152efccd08d6427d22e3fd6c02f123c467aab6eb499c733cb1d248a8abc9cd762ccf0529638732a908c8a999b5a013bf9c13a72db13ce7644b3da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e28b81f5bdd5af764998aae57a8e8e0c82b8805298322632b6c95d163c7bda701ded842209256fc75a1221696bcbe0987226dde83067241fd3e2b12a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he764ee1063b73ffa8b1b7b02b0307e13ad1362b66f57a8ddb2d2fc4843e8c0abfb5740ec16e576f04fca79cf6b12127331410d836a6f9fbfb2f290e42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd5f817dff59f8abd878f8af8f5f34924023a4180ea7ace115f92c91d0400f7d049e3038f729deafab6fc273fe9bbca668c5ab7b4977d43a9b36d412c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f04d482169ec0072f2e7fc8bf926886bb5596aeda3606a7cb8e8c098d14ac2f5a3597bbc34adc2dc8a2da635207b97bd15af7bde554464da74eb0f10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc23ef28825ebc43fd41088d0be0a82d48b505525b5185548c3ce7f44cee102d67fbf8879cde91ab1bb193a86e58951a0091a0b2fbe531f5cf6569d2fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he109fce43564af2d5e02c2303e9ab8299006c49139e202b14f44399d97a40a9034b8ea6bc00f81393a26b703824dec232516472104c7201f3317f5a62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha094951b8db8d603ffb7d39700c5f914113df9a26e2ab8c69f01e576ea8c17e11ba79368185c05e13a276470deee52f05450d24cdb94b51e5d04e80a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d5705e53cd6e82d25d21377cc9a880c4ec83d05356241538ca22a1e7c54fd36aea5bf5582c7ab12973dd3a79ecfd10a2f98b40c1af46a7c6ddcb80e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ad27c1d273ed49caaa2c9a65e0e789bc77a2b836696c21a054f967528c50f98d410c66b8250d2f03d682bd325369ff26ae2425f1555b4904e220a65e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25aa0410118d1671cb00c29bad3a1ea8ec532a2e8abdfb9abe113ec068667d1be2c777dec1ce6b70a25b42068dfcbd56d924e0feb275a0e05f0b8e255;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2eefe6fc89a731977a5f18c36c0429a154057da2b796ff45298985b808ca2b9743f02462cf17ce58b4fb34e4db7e90154f055721b99e03a63e88231c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fc081fa31335a0690a2d6918e6b6668c82a097ab5dd3ee79708b7c89f324e0b662e79eaaa5fc86da8d41a942522cd9ec502579e8ff42c135b13aa75a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4db6be1adfdf1a68b58afe75fd0f028252263ecc6da22deed39ba95e1115b5497d7f1ca7228a3d5e7d4cf187ce3de553b8dadf4c53758c7bd9793cdb2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c7f05e7fd96b4da8dc307ec82cd20de160e8d34cc9604e1655696b057bdeffd900de941849e9f9aaac1667f6f1905b69cda98033f080b811ec45ba2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf42fde0f38631ff53e4d150c20fd4fb0eff110ab6618681fc7b0b3d35fbaf0b67f34fed8feb7986cbb74bafbac5477a3960c6d456f84630f3d953815a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27153c2c57c505dd2c2247b6a9c482a8ebb7891ba8a4f1b282788010b5456188f2f82e00fa6ef9cd7b649600d95c73535b69922cc0df60504427ecacb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda434fe2c13d14acb6f450d9fe066a36a1387d0ea19da43999a6ea3b1c509e10a885b27e0c1122407685567bafe898f433536212f55a17ae4eea6d5c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h541c34122488d54a2c1b310c3539df2e8cc07511756f3118d29fb9562db711ef64f0432da04ec3d0ff2f356c380f859bfd98c8d48d94694ae7a84a66a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4949e457697fb8419180ed88d1efb956e5c6c9dc6ad23f6cc02354404d9fe7d3cc1ae45b2da19ea430dec3b78a35d6baee5f84a12b3d9c48c9ff032b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9da94e72fec0f6e3b7e4d2af3db49ceeaadc5a3dbebdc320d5213ce533f98cd26aa565b50d51d111a1a42e9a0c3a386cea1bf9da3d64fc0694efd68ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12312e208f469045f5ae50939fca75e05050fc736904f7ab1a19639da9ca2199f691a29aa53cb8ea1aedd7c88c938cdf1199b1d0cfef9839948414b97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41712450b22fec1fcb12035458e0122175fd1749135f28b0ed0745db9f4a5d9da085ea405a386a3e7d9dc97966ad0dc4c12abd0ac634f021dfd093336;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1d0b6f585eafba51ff5430fd4e59b45be3ebded61784df986a50bd4f393352a50e74b48fec541a4e0d5bbc5a58257a89a336aeb425003bf25cdd7e95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf156852a6d17ed1a911535095eff876d8e5744c86faeec0a327e3ca9792d08fb814129544005c5c1a1b16445705fe11963f11e18022ad0b973911332;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38573a367648eb033ab45e523f98e30d83242cc659607ed9ca0455d26372e07fbec6cb3b894eaeaa6baea5ae4d7ba4ae6969ef9b05d614b203da2441a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h347e9eae4c8c448a4a9ceeb84fabd6d5d507348ede2c6681bd98f586093f8c7b49934ac50a3fde6db2389d85c5b6fecb468a25630f40b610001069c74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb52f4a643a6b138e618331fbd906d7e2014df358972371d0c32041fdf7ccf82685866707c1a106ccb8d52c6b6bd0725ef942c2a782c7d3e02b464b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2a743f4193165f061ed93807ee92a607b72f58a41689569e7d519a913e9528dcd6fb4884be87523bf57fb072a56933f1f993f62c7af4e1390d55a476;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba070ec011e5ab8220c75a6ad63299eb4ea94dfec11092ddbabe5e3e03b157666d012c70220fd143e77f7f6ec592fa51f69eb5f116545d7a651177d1b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c5e8ee4d567cab62e0e5eff269a765d4e51011e864f347e0f4d24e2d40d8db3f13454215cb2a36da9bc413c571a68604249acf800284cd18e929252f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb84cd728dde19e263194a0c022fd0a46a594d883c8cb8c41c4f9328facf53d64eb2c0bda50a6339abcac82e11bf6c1354e2d66957cda6fe4ea5bf1be1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha29f3374cce7a24901677aaa342d7015b780d7b0a85c0461f12b68fc4094eed5b0c9f68955b9d5dd437d99cc4a4daf66b2494c2566f7986a7e2b972b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha07d8146ab43b9061ba4b5188f22f8d711243d70f37a0f02fbd3edb27bca09cb2d1a19267658b716a149b705a26cd85bb550daf9646f7d70f50286df8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he32441b2b3f4de788f97d91ff5875f2c9a29d90f9bd45dbc63a24029530817335e8bda0d06faeaee71042df272fb913072feb956a9927f805a2cd145b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5307bdf334fc755b5b799e934dbea554a416e455c80f4f16628340b18dcc1180b524756dca5a828f1a2236905f69c745379a616df85853f3e9e7f042;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86892dbb1bd0855a9f9bf6851da1bb53e4c36095999f3d0663a794a68bbf41e32565d0229035c449cb9b275e463c764e6f5990c2aac01989c7709860;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88219a3c66ab4f97e5eeeb4b206a4d260fb9a6c5e9f39149fd762ef3394e55e8fb6ecaf8b8553ea7db364e2d75628cd07b222b06d660b91c4d8ea3519;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha262a5b9375d45f75fd2c117fd10b89b65173f01ce7d4597f9bc669856bb48a93a5aeb114644c9f65c47048376321e1f075b59a9fb503d7824e29892c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he79b8ddd183c1498fece693d4f7e07f2371609e250b84c830dabc0c6155606c6b131b9c076d80eb5cc3afc4cc46fec4df22d8db8954d260f3541a842c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20783c5d0958b353eca9ca92e943a6ae62c56c9fa1e0b663a8e557e38046b1ce0703a48b86b97ca856c5c04d54978e3fd5f3fec1c6c957230e4ae570d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h957b29e68ccce0983409e90d61c82c7124bd4b86a864c557ac6199b401a689a5592b67c6ab68ae7bcacbd66a46c5853e55f789e207ba8a71f09d5c592;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd794040c06d0d8a4afb586f99ffda224c28e933f357576a75099c6ebd7f7da354ce08ddc18451195fd5aad8ee3d3b34fc90bef7248f8ede63638f3006;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14c49ee1ac4eb08858b7661d56b2baaab58476d627c8732fb397fdaafd2fa26c4e5440a17e70157fbbc522c91f26f71c044c9cfb2566dc5385f781406;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9579ba98589df7b89055cad5bdaf957f2e817b1044544fb108f8710e2668b2985cae85a2bb6643bffc19ab26c7a05b022a4e21b70d9ca8538cfc809de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51d2fe6d31254ef87e40a96afb3072f9dd11ce1a93ba1375bccd09b7d24ea05235ef732509f161c15a764c6adc87a5a55924b0dac0b202b365f50f84b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h776c5cd82cc35810668949eb438d0de187800071fdad362b70922f0f06d05cc0223d61a11352a93d8e4f8342ec31fa0c24567a59788835909e01adc88;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10b849c7070b552bb48d9cfa8887f03f7adc3decc97a009a6e46a08ee91829619a7f2cf274a9faa3213d7463cc60d8450cc04317920d58b9df8c07b1b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d35391fcb2343e14657b7ab91c0a6705a0a135bc765ba95f8a2d107434e68e6bdfeeaf45058f4dc4ebb47b49e3e517f9456d862a9a6efc4daa3317b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bddc75c47a02973b9da376a9b5925a35a0a2d56d0d2ccbb3d6c92d0011bd4b38af8324589275ba8f61ec2352a8aab81fd96f78b7a45b332f240c64c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he39d82d0094099c540c54660597e0ac1049f72a0a970456ef51b6beedf20e9141db7e5b5b6840c67080cdc35a26fe2b82b479ce72f413a49cfe4ddf7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cbf2b399522bec6b9bb44e7222fb525c5a1f885a39d9116f78eadcf9abce9899bc1f84fba17ef68fe4ea4e56ea82df1547f2a1360a8f5352a23be885;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2371ef71f8a7adada28930a46f12f26eaee57fa601be23764093869f01a98a3e0f27a2347e9fb0c0c6b9a7807128bfe0e39771f9ecb65ef443b7813e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1734b829b09a0afe54de6874984eb907c644a5add98c6906ec2b57ab555f0646ca47a882ab6c10108f569a08eec2773d2843e05519fae3310126fd9b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h979be597729222d4f3160cfbfbeb2494425fba64ad683f3cdebefc7d2a4ec0d69f396f4fc55ab3c8f32e543818090036ef962d93c75cb1393fd3da115;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbeca2f4eb0052085f83349f33646c2df59d29f7acd988cf014c3d06bb3952bf4b9e9311bb16378d6abeb7954dfa6902fe19cdf1bbc5e399a9403d6211;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17a227aa139218929660cb23359ca84c8bd5d3136fe81eb50f40521dc837df0479c41cacbecd8e8e3b5427283e097770988861536b587b8bbe6ca406f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f6e6ef0771c5a651c747af157f234c8c93be59c258944a8e9d02e6faab4ba79255e995354d751ded5de85fc9e08030010965dcd5158da4637b6888fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86b6d2ada969db746b7ff1415ca5969fbaabd5fbc0f4cf9eeb7ffbfa83355985ba34a47cb9f82206e7fab87c42d999b5f0f702a0e5c31f93ee582a004;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h786578f7a396700af3ee6dfd3d5eb079f8d6bab2b56429e1cfce86a95da58c5de81b77413764a998d8748b780fae066dc17afee1c95d800d45c407055;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc03034db6e9ba5a581a944325b2d0ef45c343939e793a1cc6ed2aca381cc3d7706a5887ff3593f91e31d730d4fc752d231133f1aacedd2f908de3f3b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94c92c9b60540705876dfd470d1109f9638ae349f472b68d3f0b05d2b4233ec796c6d628cbc3f6947f10810c838bb0744da6da054f83385a087814af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9869b5047154a2d4d62a37bb98fbcf9334f9292482932587cf2bb161edd851125eb06be2688a706e64e1a5dff0be3873664c4bcc366b6541df15b6ba1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17c9192227fac3fb9eb2c263625558a2494bb1f7a995c20fb5c708b4bcfbc31ccdac281c1604e449df9053795e03f1eda2b13fb30109d0678947a8855;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd004001ac732fd3154c8cf152f5d472d5a9c4bc69ac9d7929eb45546e16e644b57efa19bf8c4860964c5f9e7a1d618c54a3280c98d8bb7a4f5ad8559d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf66852d745329b879420c7f1e0323095f00ed9feaef123f3599cb5510b3175e743f9708266e9818bbe0fda85b57fb41f7fd11888d5f8153d9ad17af72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0c6506dd95734bf35ddf237c285055dab6a58b84299b54516ce7bc8c21de1f02bd41d096722ea0370ad469d87c7065e436829f957a40d7d6df708658;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8868f1ae6309b298c185bf00a6be6498e91af80b0e6900699a65def6afeb8a38bf57f734c79c890ffe1666a4f8926233a6df6ccd18ec1d8e6d7e0edc7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b5c2fb0f100f3ea19f5ccfc96b012c6ea5911cc29a2eb109ccdfb4db3473fc1a4464f4695a993b860dbf2c425e69d99d5e7ab5dc5a6b34e45c9f20ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb11ee0db185841e4967a89ac56d0f853e103f1772db74a60a8112e6e64f218bc9c5c5744b1bb83e760978d433754cdf6f817e1aeacef98256d4996a42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf17fb2acb388cd2861acb042801fdcb2e7b46281d0e7b112ff859f2b12b892f3ea3346a82d759f42a6c71deb93757e11b9459f9e3fdfd92f376d0e9c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57e55041564acb986bfac1a3556c3a0d0d2da467e54ceba618e0911fa1dab9ca1db333336f05de3e006c03e5e8f307dc8578f79518b7b76c70a4b4bbf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12dd330c16c63e1213cb7df6212a5e15b7037a0600fe5ab5b6af6027d0366bd6f1a844188c7fd22f96885ae501af197f5aea945c9bed5e28a94e64177;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9b6ddaf2ded94a4fd8b502cd4d5764695de72ba7156ecf4664b9bab52e6db3cc5e0df7c5b1a2c0d8eee64dcf0033a7b632c3fe846a44d997fd247ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf52d177d219b1a654a2f401fc95db91b4323c0501e2887bc13db72975a72765d6e77fdf02724ad61bc7a6ad2e5e3af4bcce77f6fd34a63c2ac59c3964;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22d3cd6188e2fad7d24dcf4c5699d4fcb36bbcde10634eaf0a15ec835adbd0d3c3555a5e7bbf9318127089d813cdcb9ab976f3b0fe8ac8cfd2908cc77;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h419e1173dadd2795e9cf917b6d4a95fbc12152bbee93645a7d4e617266d7d77ef63c40516701ffe09fb82046520fbd46f25cad2e6e618fd3847dcab6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2e9f18b83b6438ce340e77415da60e3adca35441ed676975e3fa14d5571af33c253fc1ebe60aa4d7d7601fd073c97d46498910c0bedd1b8d1d6a4b7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd78c07aa8a24af11e0b8408992beff68a57f455ee748a2252c2ce23bf9277288d62659d196da4acf339f43d1df01337f4415c3919671451bb0fe3e044;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5520fd12981f53daa20274fd2038ad3485635b35b7406e24e4e3314f14e65062e9267049a4857aa0fe14cc9e03d6f8b93dc9a878294bf3dc25ef6bc9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h306a8c54f1195047f5f0a30927a85f1effaaa38e77b6d062004c20eb4b4bf014d7bd25869f8e494c3dc917826ace06d7d1954969e7b1c734823c98051;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53e800ef6e9ab6d601afa28fe3fb7a9cb7d85b05ba52395e4a03f36ed608aed6b7cd64bb08fff3707e18bd60afca7087dcd6e51836b3899fda2c5de86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9f22041517c9eccc4e65b47c8cf505a4eff62f8cc9b0282ef44fd282e54d1ccc35f96c6ee435a7dee01c8aa37c170c7a6de8003f2a80c71bbe18fa81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he928363a4368af8a5ccedc3b32cad7b7215fc8f6206e424cac89512c9b410251ebbef6d50fe815ccba60cbea9f7077ee148dddb39b98cd3b02f13faf8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he83bddc731115d2b4376bac209d91050c8b7fdfe942e28c078dada0dc39cbcb83bfeedaef8293a94e4792ec9ff424a578db69cf87855763150c5fcbed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h574e55c1cff877e497e0d8a840071db39bf89c37cf908f6d02f13146549d81d72b3df224e65c516fa681fa758421b5dcaa44aa097b6fc7a4ccb9d292;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2a691ff1310b2cb7e25ac3ad46b54a1fcb47f07a05cabc8e5837b5ff70aeb24ed69187cc07a9c434c840024acc26552d8127984b12cd080847d40859;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc38b0b30c73c27b17f155599dc07e755193f632908202d68c9f82e00484a7bfa1258652d718dde0c1b678ef99ccea31fb086218f73a2f851f1a6e5358;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20037762a86a770c2e3fe88d928c9e503bd90693a95e98be42c2cb9eddd07a8e484b52bf8cc1b8e24ef9defc191b99e1ea0b190f92347826fffb6dee4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h258bd02a957f36624d7665eeef80d7ce4e920657f0a9dd67dbef2e6001f40109c2ac7d5aea320579c6652fb71aeca504d3d5ac853fdc2aaceedc4358d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60c127fdef66c88c6d8efaea45c7d05901a75d17cebec7a5c3a5518a418c22a0cdcbdc81015c92563fd62caaff585ba10c540c43b4af4ce155fa73829;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9779add3e727bae0ae8bb464b9fa1bd22d1466bb287226b07a0004842600c0a15ff8734ad6627fbb3fdf57095769f5fa5a46c6d34f4a46953513e0806;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27b53c53e902f5d59d4653fb28f7d8ca2558daac6454357701ce0758f2cbf2c59cbbffdd7c23aaf55c1f2d71b57c1874d2ef771b0b1df72b7b37501fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85fe9a255695536a605c7754db8d3979fdc3d745b1288f3b326b5e14145f47db488d44d044b6095498588cbfdbf346c0f3300a4981b9ded1a4769ba9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd1105041fb7bf07f314e12df321664ae2bb1f8ee88319f505f511ae6090f1fba3e1e66b4d2d23a7564632827f9fac276c4233b3725284972e4f2b170;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d9f953053869320c47ec310d1549bca117f79b0c403e159a50142d63b2749a72f68aa4861648af09b42904d5ba0e6c466025a8c7f20a9217f9cef268;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he49509b1b8a4cc014cbd5e75fabc6d518cd55b0419fbc015fa51a8d54f38a0ab5ec8e2cdd47919973743e14e7b0cd6974b1fa548420d229f143902dc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd814e7c9083e792b9015568777d31ebbd33a418aaad04526bf881ef8ffc27cdad5e50cc63d0484f308f0ed86383165efe849f9c96f9307a4debd6f08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h513a47130924d9eca3d0d67900a1fb3913e5fdc173ae35a107bbd22497a17664804217c5d7a5d460ad3c95256c5408c0603356619fba827ee1f3bed07;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde936d6a21bc9a027673339caf9b64f95fc7bb8994e9337e6b25114b556fcc395b8cd1adda0dbb800db3c53f6b131ebfb6150f39303ad3a56d08fed6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cf63761103439645df657f1399807119a34d2c67981cf67661e6d2bc0833dc019627fae4a9595254d9a86de11e68c295a8df8d4fb3b9c258938f70da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2408c77cc9e43417507c575f5d44aadb8e60953fdd8c921c3ae9abcc3ee459fe52041d0a6b678a4e3ac164495a28421eca05602847b533ae9b16bdbb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff0c6cb7997fc2fbeeff99270176e641293cf1d98731282c3e5bffa4e14cb8ee7717ed08f3069865ec4a586698e8cc6867de6c77c4d9e79a8adb1533a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb60d9863bf0e8822a78128c74924c427b1a852fc320804a89f594c725eba05a90b69d82b4d03e4b709073ce9f2f9f6a78b0c9a5f161f739458cf5e97b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafddeab19b850f82bdeb1fa197fe5bccbe3b8d42a81b579c78d935ca57edba1af4bbf8805e2b7be1caf91bc5d99782102cf71f2f16fe27bef5516d143;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe9da0a2737714be4331d190d3e8bc708f456e4229c75ebd0cd44bb3446aedf883e370613789b9669c09a808dcd1099af7a075b669401675d04258f59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39caa70132f063a2b8f4bf55fc1245ea88d03222f3d8a00a5e801795a4a494ea09c6d4ebe2036ea173b581c768b35df7165f2bae71a0346fbc866be29;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h648c9dcf881a3456d93a8cea28827c26cac31a403d99bb78fd2fdcaf097d83cf017e81789b6c0fa2b313a2acfa1e1f2236435cfa9d4b9e5f0d24271a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he136bf8655e7ff6ac7a12b6d10c00b340aaaaf3ab76c35e70a0aab3e201a97ea46ea1d879f37cdccaf319f154c46a80e0faf7f27d97d92eba749ae617;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he096f7c7168d0ab055f57f71cd6fb0ea6e38d15a34d0978efd5c6ff931d85e4ea3a6a6c262e83cbf200c098786044ed802757e43c3a6717f732e7fe45;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e3acb53880479b126516a4c1b4296ad66617aea66b8a6240399b162741b6ca47cd5b8796e63e118bbae07672d964d491f25df60fd3b2374ff48c1ff0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4f91263fda3f47679320d7102e3078d95ff6ff3bc9adf2a288476d2a3f5e78d726097cfd3862dd019982e8f6242b92234162391a7777e1e435ec359;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f1760253912d03e3196893c695e74df7f507a2f9c15a89666fb00442a6eed7ce1f5b6ded87896462c03eff0c59d22a8e72847bdc1e729e6b06d2604c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h709ca0709dfd2acff93c019fb513840043768258e24f7f922b21981bfd865238c8b385babee53c91a6783a1c047af1797e020818b9b2e098ceb51495d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb77569e31d19304a3a969c94902d4c5e865204c44cee47873302980b03fb66faeeef20da5c87fc83f22c55e9f5f64f4524688388748669b39ca1f8621;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e23d05075c7e108d73b190aade1838d60c6eee90dd85b19278628cf43a98a38c78114b5ef3d70112ee2655b2fc5474c90dc97aac8783808b9e3f8d95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bad54ed516396e1b0b35ac91fdc80a02e080dd22e14cfa5c03e8bfd4a434f928375254146385f60e53fbce651a35ced6b223a0ee0d55a0cdc157f00c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h259e5535560ef16112a3b772d312b7577425af47547b174ae833516b8356a0b7a12a2d27808ead571bf5e0294a90565c5fda643a5aa7796eea85ef5f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5001e5833d4059fb5cb295fe8b9aeb8485db3433df8b89e64a45b7184262b9fab21b8ec1fb26f4c5b84249916989dfbf9e7ac83477504a8f1a0a58333;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13bd59a191996e7d52a1b73cda34049df4fd78275e6539ab4c0c407f2e65a4ca5f5abaa95e859f86d4361bd39be82c2295925979536e22529e31f9c49;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d5c84eb63abf5f6a862103334b3b209bc9044c0dda268f8a523b1684f2e863c37a36b58950f5a39bdd18ff3c1636701397bc80d5d82529fa67b655b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc568ad06cfcc4e067c0adae6aa4b373dfc9a039d7f46b729d5545c73e4639a64543cabf5d9b271a0277ff91a378833cd37878e68b4d586ce3387f68f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe8b052e259b48fce4af7f8accddcf345f986ae45f7f6604618ee7a1b964d2fb0b9c271a78315d8ff26baa9d788b6589ffeaefb8ffa2d5b949d0ef721;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e9f88214fa0ef2ed4a964a03365e1ffff113c1cda54d5b1d17959da5f0bca088c893b7d3aab0c353fbcdb88d886958ef273e855667c6005afe107d41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7463ec5a2b37509487f9d13592024d0d21b04c5604211c6a6b004f2e594e4ac048d6d474dfcb394274adb6855dc03734e0c81ea1d4f767344068a45fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85487e604f9ff94c393cb6491076b3946e1b31ba0a112fd09cc1d3d04b9c4caf7fb7f73ab7d0a22cff6135c1665d739cfa3d565a2c67bfecdbcb2440b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4242b4eeb0066d3d156e5b5092deadfd41195c16a3fa5bb05f37f999618bd6be2cdf09099d0acc6799b4c6043edbfb56566d26041ebe8ad92e6fe1ac3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ce6bd3995ff00742f8f004d638b47ddc1da7aa6907dce41d0ca66e583fdcf3c7c1678d498b989567899b7042818a8fcaaefe6d6762d612617e724420;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6beed104cb54ca9214e0b8a451a485bc85cbce635e6f80ffbc6710741a168ddc9f0f9aa28053f992b63253c6b7bbe2a30da9c560cd159c644c78375ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9be1aed3a1aeb1669db75e4704a3d5485fbec5152f6675771ce9b834c657141a2c43540f39b6b441cc6636f84c80a98f92b905f59c3b73c58d60f529c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heaab652476cf8cc8470a8e01c96d5e617ed3a6c80fac4fec8dae5a700293194732196fb5c39f16ced3d9d8b4bca6902bb05e3ef34c7ec3a71f953dca5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h999b6113ab6edf633359c971698d6acb2f532100fc0e530000dafe1a11cef27fc04f018059d2e122a349b8dc7f00b183f9544086e275f61451d09bcc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebfc79fa58b933f2a96dad2ac6feb8ff5f33e1c150b48f0a5b9ce7e5db87eef443d2e00d89e1f6916d69774da294400c82373b43e3fb40d537922cc5c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39b5297cdda927ead6e44221872fb03713745f0e0d790ab0c99001798d81a896a6d8149fa63476983512ecfa84955ce90999f55151e0c61cbfe53f378;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8776dc28acd95a69779f472343476f525909bcff8c0e6e6afaf171c6843d1a80d3506774104137890cc5bccd251de3815cd3699582dad3aef79112e59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26dc6df7f4bacfad1ca297ba03ca0980b95cf9ce0434a4f490e49e546049249b1134d420b77d7454b928095ac9a100ecf56c67f1adcfbc9b535c0e8c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf60d4e9bd55cfd5fc960bfe7a8b3879821b35fb188f909874b58089febcc303990af8fd9c2392b019c04fa91b0b07318d5b061510d09c52fe8ba8a0e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a1b6824cd46281f0740be49993d35ba3017059b8cdfed129decf3e935a4e17f75fe6b571be63c36c6674c35cd36422aa7c67998045f039715e31d6de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3427a851a08fe34461b9642adb90c3df4c310b390c2e84a9229ee71aa627fdd3aafc24d6a11fa01972023bbc44d20fe9a5015d80123c7732f46915a6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22cbd33248bb25997e77080532dfa948e2f1f463d52de3dc556dfad9fed9d497c9fac22c26847b34937ddde3578b1429d8bb6d2055f32a4c03a63cef8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea78e1846c8796b1669f6e82da33999403e263c310f9e3631cec1c5fe818eef98eab2b1efcdd24f059b5542a358d24549eaf9033168fcd8137fe0b1e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h599229558560caaaa6ba25a8eda5d9f6ef3762b331c18d060b6f3669af1ed36fb2994aa124a86a8d57c3509cdf9ec336b7a8749d556e13571dcf25dea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d479739c68a5930ce573fed55c52ee8821286c968708c083c9c5d4f014a99513c4bc55446072040d7c3c2c820c6d625b03a88c5baf0fcd275084318d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h296901bb38ed82a4017ac21ced15319233f856537b4c942ca0b5f904d8fd2a36991faf35e2592316c41ad8086e534414961e7a4c6048893960c2d9f23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c409fe3ec7fc41a7a8b3c96fa85f91545ad50716c86fdf05db1e074dcb199a77d292176f7afbc22fc81e19575bcf7035c2864d80a57f5fb6dc21bb1b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haffc4ea42740fffa4e392f06a0ce171a14dad694bc2fe74b6ddc9afc1afc70752cae38097a88009f606492a3ef783cfee439e19f80cae7c435eb34999;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h536e9e7325df41113639e741d5e9e4754f881139aa8807cbda0ba501ffd9544cccf82b1936e8fb1dc27bda3c8b7e91b4f0b2d9a476862817d25f8c008;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h432b011f417c022a3cabcb7564cb55f3a4561b57ad054b6746902791472af2204163980edb7f10d0c680138e6715c1662ec2c918e092ce135641e204;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba6b22fd2df315eae977ed8b7da665a2361fec612cb265291367385723a4c6e302dcd28f089f585c4dc6d594d4d13a8ab208c29d0394925f339003c45;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdeca50fac818cbff0a98c9287477cedf69daef47bc3a612a08d24cb8ce41a02a1fe60735b9814fa7274d2285fa2252de4da91ef73fd7e7f3f3d58cc3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc67a7a1e0e794f50cf38cd7a00b125cb94d605036dfcba13ee0199002b502c14eed4a41f476dffc8571b62c1a3fb469399d03cd2ee4940a79a702e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84f452993ce2f19f6e001ba71caa20704c12cd06ea836ce09d1c466ab171ee4dcaf838a9c3d266bb184a91e047dbd61689d276797272464ea3063eeed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b094ef84487f8a44c2fa2d292c537008b6a51aef00c7e761f6f7a435b3c04ab3fbc00cd789a1f49f52a43d9790114afc6e4a3aa7fadf4af33cae8415;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb4dadb95b5a86cf4eaf08c904b7ab27a0a3facadb4b3917b5e5fea014e83b0a1809280446eadc540a5cc62dd2db9b8c2d1d4e5718062b2af79ebdcd1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c7a4d956d36fd335ea0c225d0e050bbbaf35391aad15d81c4af846280fe45925a91572b3180e340c9763245eb8e3511fd911343a0d70794bcfffd841;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h205e437a2562b29ce88fafeac97b1a3029471ff50d12424484ae71df3e01b17014fe55163fc8f3de8aa3f6a1c55509b126f747cdcb5e9baa91f036a5d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0fff3943e9a31505909f4812ebbc68c5eb8819cbce73166829a130d90eb4f46afa42f54bfef905fc4b24e4f3407686552dfc92ab95640cc76745a1b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9308ae5b97a147584e4a18f3d529fbbc65a92d4fb0f09a9b17fd47b34ff7729b521c17690bbd969c1337efa44152e07d5a79520650270d7816f5be23d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3acdb44ef6038cb2383d83e7f1aac921794fb37504de6e5cdf0ce5442239192fa8b787937f19b896efc597c1d3554a05a6be2add3bb96775a3104b171;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea0da5aa9272c3a981976a23f10ac7f479404384f49e9cb3b6de3487bda9c6d473006321c1afe7a51dec5b631908f458b1648897158e26335c8642bef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2060257f0b0f403ee4d068a59ac1475d63fc13392a953571becf6c19761174b008e9e90d7fe77bda6e0c766d2c02541aa01fd36ec6a5d1dbd003d38c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc38af61ef0e8d1a0c598c0297f613201b34b25a3079c9b31f301061446b23136e8461df472a7b1dbfc3dbc9ad11497bd02041b2d428ffac7b4b740b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88a00ddef843bd1fcc5fe66160013046322c7b271cac444421ab72a2ac70633a23d92ffd13c086635e664ae3e340f63fabad0f20b5903095fa34700bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b54c8f738954dd94dc00940bf16ffd5b5c3db601048ff6e3f3600e7e6d74550a0da6b4d37498f98606e9695436cd7190ae4a9f869952ef934ccdb6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h322437966ae864dac903b3d801b91d51956095d80a8f286b4dd8ddf4ce26df8731ec4cd1e083811939c4e9d8ebaa6d0599759b92daa05b3e270ff9a7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3335ae5166bbfc01f7f30178fa7ef7f2502f35e4daf44c40d3a64ff760af61079c8972e9220f68b346bfe36cafb18377f18f5d9d902939906a5c95f7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45ba910c16850849bdf804373d45510db32ad9bccdf28dbf055c5bc3699a081a1617848e31ec954ed83d2aaf80a5b43e6444d5b5d5674f9fc8b29d004;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9e4872ad829364d30f6e13f44a82ed6f2626eda447c27cb4dd9f1e9970221111d4be27e38b0bab0efed2e66d08f1c744277880b05fe6b6f90be280b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eaca33eb3abb37afd55a767d1e5183e96847c3b90f2fc24f6a612a689b991698749a9cd17a6546e11b3bcbf72993d9b1980958a8772a0a777b1c3629;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bd0b5de08ead4db18a88126f79787787f1d9e3bda2f452087e0aafe70ba9a75ab78209259752f1bd65157291838a3c3116922b95f9a145dfb59719e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc60e0f994b5dd627f8fb98ef3bbb75bbdb4b9b6b063ba46fe8e548cb729e74d0324f4aae020907d436bbf90ee3686a7bc2d85291b541c6c83766f5264;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had80a8be7b744eac066c03c39bc8dfffa300ef06d81c26dfb20d12daf762bf841a7c4f4a3d2dc2aa6ed7f27dddbf3e6a0e1ac2305c381d5f2c3584570;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h629b41698be240a6fd01f3a7fb709755fc7895b0a6dcf40b628f462c6663ed73c8ebc4a08e09a9639fbc2bcfbc893ccbc548b9b1aadcbe17df8049cc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bb83111a084a99c95218dde668a99c0db39ca1bfe6d4162ba0f65aff1642c647f04ea90e204cfe39a1c9f70ebe9fcc90eb23e980e922891eb5b5000f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49e303bd887a96117eac534385c311c612324ed4db89b7b85065878874a334f0dc318525989aeb84c952cf0f4132d12be51660723bc21b51b4b0c6ab6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e54230d21ca6b177e385a646f5364a574a388f803eb7978ae83d1a5028a966eab5fd4bb9f3dea538fd391a5472f4d80c2080f6b126e00dcf49a1528d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f1bdbba187453b177fa05bac9766a4af3fdf0ea16250c432d36b1487b75cba3683a7a09db229eb7ab2dc1be319a1f7f8b0ea668c7bf69fdc291318b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38f005ed4197ccbe202944045db0d54360e94f63268adc2c45643eebd18aca67f1551c3cd42c9a90f556342e3b168224ceaf306ffd2114f75ae39cb6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c27bf6d925cb7a6fff8acf2014738c96777ae5bafd7587334b6b9e16920c409c67c0c80488779dd743e886c31ed7d276469ba1e44b0787274fd3e777;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h882ffbfa155e966d2c5f4e8a1de6c440635f521fa6fd828b2737307c833eb51bea94a79df9de668fc20346ae1e3c89643a16230ca669614aaee8fd0ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0ac1353f3e0216aa00ca1879e0233690fbde74ccafff770b5226e3617d3af4a5865fb7b69af16feb78283543baa4f1cb0a84a180b5973cac7894f7fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe3b3b388a15aa112506d9a41693a7db141ea6cde219f243e59e4ee3cbbbc71d523a3ebb6eb0dc14fb8a67ea2a1604bdacdbf8e67540b9bb2b7e75ebe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca28b29b2b0a4eadc48eaa7b49b03ef55edcef494eaba5209eed42c26248fdcd7dfa96597e466b82c52cf1c1648e4d0cb66ccf05a3a22c076b7cb24a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fd40215e90dded3e1346c28e83d6e6b5f5b8e1b4b2d0830b81f7c34746e68866587c39ce1b9f572e51c6c41965545c42282075bfe3a088d3066ab0ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6913c0dde7ad4ab8c3d84f9c22515876cf929557bb6cd29ed1eef35a6b572486dced037c2b862558682dd09dc4c0413915f4f3f55ca2bfe9d90e7048;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65afa0a07e39dae3367ee204d1b0d7b130e0ab38951fb14320301278d8fced22bb7a7585535bfb52ffba4d6c527e95bfff1653864f98898537c02e715;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d21059522e2ff77f0be55ef82e32bd3b3e10270c9a457f34b38dda771d7a1772b8f199eebcb778dfe17e5473ac69b88584c3b01ca05171cd1c223a3d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf07ee8814397e1011d7eb8c255c1634772995417e056ee01efa546807c533cd97c226ca196af7a586dee1d8826634fec486869bdc3894ffd506ef2d53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51f692c4473f753c7dbe387545934b3589d1d6202a9dc66f30a666c8d7649002344a26d19b885a6b722b9e1ea081abb5cabdfecd3656fdd960e206ff2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha84d8d6477f17eed58e03691a84372cedc6f1baa53fe23769771e4187bc2daef280db89c9e454f7e76024abeedc7441eca184c694cbdb010913fbb5ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7897782e4cad4e99b881d1d11472f86806b5f0f97781edb83c5aca5718067997fc4c83444623682cfbfdf7ea04a77b4d1275f06c33f9f2ab1b9edc220;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52b7ab43fea8b4eea87e2da7535314da03f05cdbee98ebcda5b955f5969b6d3bf1c0dd52f2e60c739994d709315dc38f4a026822633ff433c92cc9aa9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h258961b7466a6c395809475fda2f7e18591cd3b051010acec794185ffedbdae698d86dd262a68f5a08cf85ff7ea51e6048c437ba9c163ec16a89eb349;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f0caf54d13d49d7554fb0234ac93ce6a5b3579ec83194d5a271fbbe6abaa36603b171b3ac95c2198747559e3cffad8c65fdc24959066b5bb451f2f89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ac36dd615a85e498fb27c8f13b92a64e1765936d0d9308274b27f3b6f071f1da6d8695886c00d9cff82e6f15e29e6265c59d0e8dcf80c510e91b0b6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fd674fd06f9bd6d76cda0cd339bdae7f0b11685a9cbb29969fa7ad7bae49abef7504d8be30b14553eb57713488caf9cc4644442c9431ffc09278ee9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82e251e9b0807c6653f4fe2b98eb3b4e32dc8a5dc6d7e3591718e1268557c598ac60c1e07fd741748a7ea71f0d39f7ebf02436e18de90c2889310bbd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9f9bc02eb84daac103de762cb03c1836d610cb9856f2aec0d3ac549524e69e4340b3911d69558e629b4e58e23d26a4802caf6f5e9ae2075d73789c1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1df046723657f9908a1af275eb46eaed75a0e0365d4d4156948dfb55fb79f3bc7e86511baace7e204a1d8c31fd02517b29f68dd6980c1eca767d0634b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8be879d26f80d7646a2b91a1f05b3828ec21dba1e17de461e74cbd0a94bcba7bf4f18ba13d5bbeba584b1c721056111fb68c25fbe851d9b946006082b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c72e855e65ccf61b74876b076a46f600905cbeb981680b3e60e8eba13c1cdd7da2f09768da573d1d3f888d361e89e2ed354deb6730fd01ee624e771a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h946e7c54506773518513a39e2096c0c1b9d5642b1ef92810110b2da1dfe0ce3f2854cdcc36dd4fb1d67e12757047213338a01946d6715749519c527d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he85a8e52c6a9dd33f3de6a447ee669783e4c9cb6efde284e77aec18a220cb2865c094e3157f3700eb2babfbaf5d9ad62bf3e6969eaece86c3c487cad3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44028ef83da9bc28906c379d4ce510b54e72eda42daa60dfa4db893ababbe7e45d2c7c116dda95ab756f698255040cb9ea8d14ec78a1eacbb76112987;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7c782874c6e5b6a3bd6a0d614dce0b3f23d1d94280b61ff2c03dae12bebd08022dd2c8255580fe87dab9969adf776c94d8e4b76c62ecdbf56e79cb09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1a8c636c13c5ada176192132f88dc6b6ed5663472d2dea97ab587b4462aab28b2ff39fe2ea84499e43855758951ce35a3c93a2c4675d648e3e09d1c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ca58e061721481d3c357a73961076a1700b52ca78921e919cc0820826202713d7e9b665553ef7bf060069b60e715567f0224779c54cd18c782927997;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e649e3b0a489d0307724331a73ebc3fd79b2aeea2d1e988e5eead9f46caa77a46118e128caeb4c0324fba1614ec1c692af7955730391ae02e71c8af5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90ba75c5b9661de91f9f3a1f4ea3a33d551335a37f624e1501e2ece268b199d0e29424e2e115024412fa82e7234a52bb08297183921c71e073c7dfcb1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h461165ebe5a3b10a40f55e90268ade72bfcff47fd131a6961875f1ded512201025e867af7d72448ccf36e05b0b97f37bebf57adf69a1f67380ea630c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ff3dda45650cba1d9ac5ac39d6c420098a70adad5d7b06344b929577025a24b5ccc0e37a0ccccc851ba6f6bafc37c1be5b7bc64c4629d7eb58a5e5d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e8a8c228782d21c9e3f2e0d7f0b87e5ab9f705b8d0c9dd7e7d639f7b247266420c4ef699847f12464b1ea91b7dea0b652f31b19bc6cfffd8b1e922b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5369963df70c5913bc2e55c20c43a78a8c34e0cf3abb80305f35a972473a5c16b6974308f9dc54b9355e9267e69181ee0ec3d18f616caebaf111071e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c0db89e3866372ebbc4be3a77ed137499c96d70e1d55acf87187a323f773bccaea93fa65a455d1a25e31d72acd7c47d8eb049b738a5cfa9e8078fe25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb34372ec91981095840ea80d6e3ebeaf851a604549a2c38bd9a483f54997dd23df873641e3be13bc6453c011e0c1c741b02a551bfbcd6745fd00fdc97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc99970a8db0544cace6136fdeaffdeb5d81040b9b7b2c727753df8acec60f8c37ddf4e15e90e95f4c7b9664d456d8f0c119ee264980709fa5704323b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86b8ecd35feb8d4f05dbd70cf6374ccf9ed11f1e6947e443fc518ccdf0e1e73db4e304552ee0ad7fadc876441aa83c9900ad1889138a1341cc72e39e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h549721d3869f52f0727d1593526cedf3a2ed16cfe254dc4c808e2a5e36e22f8dc8f847f88e5bc16dbdf2500003573efa2d7786664a219af89438147eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0d8787690855d5ed435d1936465ff5eecb837b7e8c3be7ef42fbd6efe742d439bcd8c6ad896e2f5ab787fac7e0cdb147f50bdf2127c16d343d58b784;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h217c6ef92e4d6ca5c3e7ed01fca36ae6edff71a5b5dfb6dea50e16ed93b17fb032ece706b5ec89e38bb065bfbdbde0327252f151a87d30b72d06a314b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc4a102153072b281782bd47edce0b5727e884bba51818613d5fe9612a98061be8379bcf615303cdae5e767d5cf7f77bf0f2b332a3b7b56c66cfde620;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b0563348018e42bc7c59151aad0b2a0fde682253102078239ebc8324fad233914e371faf9a87d0e087ece78c190a53074f5af7ba80bddacb4cc5af4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f9e7e88de1deaccce91f744d37257777af57bb5ad4abd5304d0e6d7744412a5dfedff332f7f8019d3d9c76d50307c4f01b999146d3e21e34231be9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f9af7182f17dff4b611e61b3a3789bfce5b8f165410b1b0e938806bb904d7220f3ab247131b2b960b7396190637badece4b935627d9538d8001ddb87;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h362142a12ddb3fdb4d8bc3f5ccc75404356d5c36ed4cdbebb895e97d04478a874a462feaeedd2f9b84c232b18be43a925f022601cc83bc0383c68e873;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee13f6d4c1ee844916892683d7bb6606f311a28901e1c5e6cf2ba47e52dc52efc61d2de38c10094bd4f2b43ebb2b3f349cd50e16b3734ee2b84a142f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd56b7dd7c148776243f3b767e3c75d5d6d7cb5bbe619650f52396b6032c8ceea27ad44102b87fb4c317d34ac8b81f994e28c7909a5a6ea3d446746ec1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53afffb17f16ab1ea1f47c2eb7c9791713f1229c998c4b0109cb10a4981d83540366adff591f78ca781656010ce82df450316a6f2807a16dbceaa1ece;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb206d628a34c9a0740d4d90254aee0d9463fdf2ffa384f2748da0e729b4069f1e4a6e42d75906d2bb3d6eda4fadf71009fd6f35e9af43a8f3926e57e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44c873eedee0716c3354d706a89480c91ab81579537298a3eefc28a6841be4e91585d38714dc109ed87880cefd38076f001a3003ec3573ef37fbfcf49;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75acbf1dcdc3dfd04c88dbea4fb72012b69cf2b3b0b2e7698068c3b91adcd2c2a0bdb09f1d2370fe9c7c13f441e7a8a1909404919bb08ea4da29c004c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha53ade7c5d8a73a935d4f05a769dad49cb21ee68f784aaec85ae02c8c746614f2c1eaff5b12554cc5a3571d3753844c03694924cc9d39652a33a98889;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc60dbef67c4255ff48027c69e5e9c2ddac45f2c2bcbd69f7d4bfb4f49493be3d7058ba9703a9d038191e7f90d18888198e6d2bcec064dd5fa974ed5b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6000ac63ac87634302f7b5651edb733cf92b90d77f13bccad29b35c0b84ba83426cac86df128028d00eb138689c8bdfebbee4cc12877226a2d070deb2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd698a25766f1ebf9ca074d11208c5528f402c2290cdf88c04b67f39e6da2c6e79f7c9a7a8e183915e6c88946ada756e7789525c27677616b16759a50;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h613dfda93ec04b1fe195fd6711bd5ead6b4c7dd99425b5e6b7c6fcbb4b5cc88bc1f77ee56816ad9a481b7e937a694f28a79447e06d48099184ea76931;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha864775ada267780fe76e2c5a8844ff4981c0e103af596d4c50a58c61faee3895e76c2176958d22ffc79d8b89095d717f430198333af6d54d5e51af85;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec1709f8c60e10626f5ae0a6eff5a71229e6662d4b9aba1dd0ff9a2e2e5f954437feba6bae751a2fea84d113b2da3e5a7b2b8fddb14f7bb89438b6940;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ed12b34a8efca8e7555dce55f011ebb6b47b86ee7bb11f5020a50d7f2a9405f737834ac4cbacbb1031c9ccb692c59bfa5e704ddd457b0ae3ae4b9df3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1c7a1fe9c5b4d42dde4064701362d06ac2625cbffbdf6064fef47d3cb6c260a414e85a0c30516e62b9865fe0bcd47d404d104a9364cf9ecf224e2922;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23329f3f70ca9ff521d126f216de3187e257238024bd5ee1242df585c8466d961cbc8d5b7084bdca3e31caeb1df3547acb0b8564eb77029a425f0cb3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31ad337537442ccf850e8f978e51d651e6e539135468b06f0177c916367aa7729c0f3fb9852360e2886e533ffea594b213b5f64115da5ad5ec7a6cd91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h109d7a4370d1cfa02c7aff084ec05a1edd90aa05365ec7acfd8a5a4b47c0dd8127ad3c2e7bead5a5788873b8bbb8e716d8deeaf829fc56bb893f5f91c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85cbcf05450b83bcbd4119ae7cab0d3710a8df49051140b5f812c21d3d3fe4b23e5a2f1ab14ed11c175f0599b30ddae83083a52c05120a9e59320b508;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59577eceb9531fad8fbe8e965c877cd4658cbae9f262ad64871d7ade362191e1589edd4005c4aabe3426e25a5ea903173b45af7b494129477895918c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbaa0dec783a60d90870dad6f08024be2a461892d3c64d0c3ca893ac0f20b4c6bd6e58a006a164841b40dd4673e016275fd74bd9b24b5e222e2a5fb8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6432e01ae659de7945a6bb798ef3c021abcb96559fc6f8722ed0b3a6490c5ba4236eacd9dddcc3e531575b7052afcbb6a19065972f086493d63fcb008;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he985e56d74508cea30b4349dfbd05a977dd787cebf06edc2156f4460f47eabcb48e896b38008a90e8e416e6ecfd4dc117a777b2d2561e84d88423382b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bd86ddedce7c1afa93958c1c42ca6d19bca507d2d96ea4dce010e4588f86bdf8e89797e8d9dff611e4cf9668af7d8fb3558edcb789dd57055b3e218d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eef1759375afe19809eb46dc691ae15d4b804ac6fe7376122f9ac1be2444f0baf4c37cc9b76614cc49b8a227ab804102181f52c637f32d476b41f05f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h621a4d1488cc8bcdc6aa4702be5d512c1068f46208dc6bf12ee6265f46e8402d4ffd8ad9f09cb1d5756620fcf2adc4ccbbdda25f2de9769c4a2c7416b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb06c0cd9da388cb24beee00c3a0baef71d05e2070cec64a05f14c2a818abd14c58805c3ced71f7a96011e45dcce6288db9c52739766352bb133cc4df1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3304bd6bad14f8778e3e7881fe444f9df1139f4bed5cd27a9f1f8f07559177ec8e42027881504e6790380a28fe9eb72677865761933c9678e169b3c7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78796472a83126131fbf07a017bb943af7173c72500d904529aa2fedf29b26197b863e84b9265fd73dc71a11c0036ca79c49d47e2f79b4ffc9a03431f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a149d94052626008fb607a2abb9f44c050049742c76143fc21674e4edfdfabde058db5fde19d0cadef0d5fc215219794b62b5608abf88858622f446e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h883e70f3bda248b0ea1b445a1e33d5fa7bef5896b4c6a8bd43b182432b267c5ae7b7536f7d51e1a4d9cf36255c5914d23fe2d33d64c0e8e7ccab6125b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1d9ed93207845b4d5db00820cc9070b1269aad13c41380b0db1f716c7d20b97e3c5474a7211bc4844db9559b810c06ffe44219079a0f5bb3dc6a2c4a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8414b5abda4ce7d456eea142895095d10ddc3de73afd96a9b82a4c59640871641e8045029b3760be3a2d12484bded3573ba0163efa1c57410a13fcdee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb52183a744a13560da76e36676ee0f32296e334f9238a69cb23c1932816813177fc700d304f39c37f70897accfe091a7dc45ee8a6c4b2ba3dd61b0342;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ccbafd7a79bc9cabe81b27524110602e332276a60bac9759c711e21c6d9863a104d6d73bedac317bacebb4b09459e34186b933bc6f451dfdb4e74059;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81fff64dc3bbebfcdadf13d90c3bbc109f019ea40dc62f69758465666d22c6e1bccb07bc7f78dbbc75d55cc2189eb9e349346d5c5fb2656e2e22bea46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefa7b1a8918a382813496653dfb908537ae6e4fe1cf39aeb0656d6e9d3e019d304ff92eddf50a8353463aeec6b129bc2a738baeba267ec44214264012;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb47ce2ebdcb09486641893a3e7bf9616dcf5c11bfbb2f3682c9103b75fe695b27bf9d5b201eb5f3b78d6931a8523c65259a31ac10baa76d263216e7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4d606d419fa5808c5bcf9764b3273cda89e114bb372be6ce6e455a875afb140b37a557b6fa4982d3a2cba063a1ef42356acce91bb49f2fe0e82e02f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7157913d922daa83742a46024f93f1744490eec6401db1937f04385910fe632140118153bbbc7c1715acc00a6d02d6df4017ee1cd985b2a3e04fdf09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac5a503095f69b8c2167c804c742178762a9ef2833385b358bd212c8bbe7690ad84347ac91897bed1a7a53ed56e999e0c08faa977bb27d2db5d22180c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0cccd0c7b2fba6517842fcfa1357092ce87bf0db5006a76d4e503c9a436fcb46cd6b54b7d976c4da18e5bedf76d5a2c6ebb0aac6ce39bf235866ca3d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b5b367bb5ddba4b07be571010c9402a9e30c262f6f2362267b04eb606b9cd2edcb5034a60eacd4d98f48188b6eb37d80a6c7085557bcd36b45f8e570;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h534d93a66464ba7f11ac82cb984b75049ee38e1b042d934e7b84d301dec8421cbbc6bbef229f383a920c8f8e4b38cb948d1f90e029c099ca4634a71d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb8e8e9b31401c2762b790b6a3606d26935f1e055c7605bdba4761e745e9d989f29e70a562e72326976722c28c46cd140042d0b3633b1a4eb006093af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcac083e103e588fc204382109020195616cf1655cb1abe298cff8dab8a9b731aec171fb6c4f2aada6c34e5d940ba3d5d2e8806b2fdd4f484f12d590a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f5141c96dae589202771333a306d3213c66d6e7ccec4a369c96d96bc6deb79f71cf66adb8d4aad69e6d2e6668b91c5abaea06b8a8997f64c09921b28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25286744d50114ee6d8b996399b34f4e128845979469bea7d1b1e794435adf6bcf3efecb1a21c01a2028ad3ed2958630c87ba285dc52387f121ec048e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f8bccc2bebbef9521f637e8b289953d464e8571873a3965aa3b699e433fa701ceeebb2896fda3ddbb9926bf571545fc590bf3cd946cb4d5ba02cde96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h550d5bbce027de75aa9702488027049ef9816c76b58b141818425534f0cc6284e9ba7bb5fdab13e53314f5cf0037ebb3722bd9401c21f882eaa15c7ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3662939d859fefe3bf5a943d991fb6fdb2164307cb60ea9c6c52d257b336b63bc0aea331f12ea6230b6c6a3fd5ad4607aedd9fca54cd0eb398ee1cbd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4eccc0e8e12b87f0cce2d29607416c97aa3195d911ad77afde2f1d278b307f1690056e2c63c0a9408506e0fc833cbd375d6ae2102f8bb77c88b63f19;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0942f6f9c61fe4078c4c0e31da8c4366540b53f974108fe982bcb362a094f22ed9f5c03f16463e06468b5715a1371f8b0e056a256ee95ae09e24bef4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd4824267da638e36a5bcf57e30fd06f6356ec5f6430cf90d85e740ec42e97629690a4391916335e2d4d79fc1951c50209a104093ef99df4fe32207bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf16b6b4a8f4eedb26656507330e78afe83f0c8672376316fb47a7fe64708501971adab15c46e62c0a0b6557d6b20e563c2be856811f711bed7c1d01d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e55d85a08fd561baed62f4547279f818a60d25b9bcb88136040a43e50a2276e216a0ab1ae209899b2ee292d3f76f0642470e8220a82e05cef3226f5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe29a2f2ab7ddb697d67882a04b0e0935b6ba9fdb3e23f603d6bd4f09a499426dc83ba3d971f008c24ad112711cf5189dc0900093871287344a692f49;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he033e870311b0a63c214d6a228b5f2d1720b9888667301f99f72f58b45a65d7b4a19dc4c816db1c990619af13d9876da2ddfa573cfd98e86dac91d6b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd437cba0bdf2d4aff493e6abd0a24d8565b6897fcb0b7426e0b171459d3cf65b9974dc1a5019a0193348006798732801f55fd8d2800e553849b61667f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60397d8854ab32aa28ed77a313d50dd27ccb9b5059f57505a71964741e3de3845532cf70a3d095ba483e48518cf53bbc463d973e9080b4ad1b071ca39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21da7cc551eaaff9920edfc7ce22e51417e61b464f7ad99f3ab5e52628b8b1da8ed64cd5c18428001f112cdcd2d9d02ee710a9536290af4260afa6dc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdea6dd60b4ad51d71dd2075f4756874a17b1f28da10d171ba36338d0f26f41c7a2303b930b23cbabd129d1fdfb923a1d9231333325295fc7327d316e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3676b33dbd851acc5f64823875d83ea77a1fed6cd8cef5062aa87b19b7ca2b2464107dc78cea6ddfaac745b25667fd8b77514ccca2c0e0451b320ea8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a780fcb7164fc3931b4247853083718534b2a32633a3b2c063565631a766be881f337a20dd7c7525e2c415e050b6cab6ed04c8d75b81226651af9b30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44fec722bb80067cc8d37b04ac4f2418bffbeedc1bbf54a53f5d77872385b428b2027b7cdf14765a7a2eb3928bd29d287d00186b693d3d1f6fa6aa802;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bdcdd231524d56a005262f3232d8aadb732afa10a1ca21f0f51a57a66a65a6d1e3c90b0302803adb7787a15b0ed9c20a0562dc11ae0572b9b69f53a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h916051b97a531f9bd1442c5913a638c40d44a06f60eb26379840bf5fbaf63746a72d693f19f72d99d039b4820f6a23bb788de07bcd68bcfc319f319e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0757a33f56c7a872c48c157da3b73c9da404c123946517a80a76b66f041e6ce3eb209c2a39fbdfc8e0914518ceac5671a87e22fea7a6625282244c11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cfa289377249c98593103aecd6043b0f1fe93e1a1938d5bd476682959d74d7ed0e40f6518575e2f377ff38c84662a0ebffad192abec23d0c40c13f17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf57912df2338fe336b7d91262030a09cd4ab7b2e374291d3cb33cd6b22a72e5efba4e4255370d1e8d83c660013ec2aee87b1a52ee869fd156a0470702;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h955100c13654b7d54f83fc98524604df69b5e9c7377d81b8f397cf15d0ac641c85d50dee88ac909b029740d270bcdda6737af0d0ffa0bf18105e5ca25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2d97e7e6b48b17a3705d62a978918635e28a72960839c50738173623053d116d279c1032b821971fc246ca138736fe0f07120fe5b41bf2fd21d8328;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cd6eeedd008997a21339fcfb59803678cc29b1caa95274e581080837aeb8d7225e01268227221c0969c6f9f8760e70aa4c166583b6d5ed55b6a88451;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2cd519479ad0b1090179103157c67bbde693bbb9a53e333bd330acadfa6f3bc3ba93321b9702d5f62afd2ded1c93e4af1982da51be36b131b1129e47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaaa29d2457ec604ca3dfb5884c0eda400d643262178028b6a6432c814d6191357c605c1d76a13bff373a3fedec7aa0f1554dc0a7ac0c915ec8ec3f5c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b96e1da6e948b0fc5aa065259ea35e395c458fbb21803780d51eaf415da8811b4df0fead040702a393f6a49b9f46a8c45dc473e15fffcc93fb735b09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h237d4059407a24e97e87d5727b412c7e7cc69355c8ad93be9dafab73eddc652ebcd841b7efd630951006213a8e794fbe69e893123ece7c2565f0af35e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1298204192ca8344e6b543a7d33c4bcc43d26751eb1622d8871c80a5b00176036b95dedcf1afee7f72dd21fd870240e299d5a6007e67040c1489d3d24;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb574047b005d5c3f9651f7aadc71cf2be000aeb981660815ff7e1c564cf3235b76469f361ecc382496dcde5131e670916414ba2db63df36c877a32c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee6b4b19f971d081c7a8f761d0901a4520579d76b058e0399cc31032d813290480fa0f31853b7ee7992740f9b1aa00c9b6d9dd1e5d0ef17c847eb8237;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8438dde991fe56a47ce6f7e50a11380fe78210be3397ce27c4afedd60a82a85b375e440f77ef2e05aff28eb2942a82eb54a40b9cd521f9ff1caa0341;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h859e70c2aa4f4ebbb70026135f30adb401ac7a6701b123ac1dde6e18efb4cdf7f3566869ff31d0f0d5f5602233152b6b6f586a7271f93513f0c466eb7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5193bec92f53261d7f76623dc185a7075439602599a6226f3352030824743210d9be165f84b2e761528403c077e99bb104f54e070bd7f11d7b06c71d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2625d6bbd24d42c0e9b88c971dd228c427a4abf4ba58fe7dfb484a178afc2dee9c72b030a69b9b7f4597a628fbedc25adc0bfab5bdbe27db59d32514;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54464f089a8c8f5f517a498559869dd8ad2f242b91487083fdcad8ff3f877baab62ec26320dbea3239971ff33d6d0191a7a87e25809113137fdbdedd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59d28d0581d16803a99fd6964c7eac6fac2dff03a3190d7183e678d6f54ddbd09f63a544b3bf300b8123fe9c5fcbfc99900bbecc730304f93899e3a69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1f37f4babbed3d2e5ac2283979c9eb8aee5acdae9398536eaf96bffbf9e9356e2255a92dc4f9b02987629d8d1fe82752727a911141d5df6b6aa83b28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc43b4f2a0f3641c7af9a18c501a4448b1bb73b4539099b624ba5e1a04d793fad39c5917978c0bce5df40d9cbb09d935b92e46b87d62342f15223e76e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7ea085cb4f27e4e577262ad3de5fb4151e9f7dfe6c2fd8d1b0726a17538991f990d09105868d688705c8937cb193c0693f2f374de206fc15f997ec08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e8b98de2aed548a9434eebfa20acd0315dd86f75efc2f8404151311ee4dea066617544e53293f40ae567d3c4f660ec367db808d4defafaf25cc174a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2f2b3dc812802ba21d847e4fece8dffa88389e51cadc2f2f29e3925ef7823662053e0f8fda829a8b77aa2dd76644e5075f73019d43e5dd1a0bbdc37d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ecec18180d03962584a0b9473dd38a0350475a27ad4c1f2389e92cc865e81cae8c937b1343bf32e16cb47d0fe2c4de6c51c5a7080ed7f6d3fd2c3f38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h818b6f2752f7374bab0c2ef85d292bc3ba930e668c80a1821e6ffe89e400aa8a225759ebac62f6963fa46052c730501538098d0d59046636484b248a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92168d93d5a1425be837fd162953a5439eb4385ced667654caf5ce3c7cce83747ebf656c043bb5cf61a31e8e72e287537ddf56743761a0ddfa94de89a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e73ef19156fb2b6c5db4fab23bbf796dc5dafc89dc7de1102e63825926d0eaab8e95fa96939161b7def42c67082a017c8174fd5f8c2fd479517b5b63;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h883087dba608e37b8b561981923a91e3c52be0d70eeccb659c0fdb05f430f1e619784b04e52eab5405f8284dc04e85ee4b7f411cbc4262209a7fef61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37686b3b79e18e335cacabc6f389807cbf5bc99505c9a1baabfe4b9bd8e74fbb2a505ed0c04c999bb1385aa486f49253a5df80b53f3341d2056da2407;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2aebaeadb81f82781d9cc284494e5b50463a448708d97df5b33a9a36079c6068f0cff927124f3e5a70ab2710304310b711217137834f4f82effe00cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h360ea27e182e78f4f4bdea48fc921938e7af2b6e658ee4b23b234f9a775fc41f3b0215d4033a20725e574f2d10421513f2173773aec210c7819c650fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h692ae8c5fdc6a6d53467cc96209a53151c21f0311f6d71eae1c8eb034fe865a2967e18cf76b81b08383f03eba7fd66b4e8ed278b9fecba28b351f9ea6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6061f89a03ece5b61578c2e310ae21a09e5710294f257e256b88eeda5305b9e9b7f45200f0bb72abdfd324eed9304d06153fc9012431a3d43bf697b05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4e5d50f8cc5fbd80a8187093b662f625b68d06617f21a03e286b48cc78b9e53ffb7ae71c16c04fc89773271b51c114a1e611a4ff243281d1a76c23e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c156cf1c75cbf3e6520537698f20c9ca81ea025950196d13b94e59bbd71ee00f714770336d4ef87bfc30e41eda058c138731faf834a3e88cac59a890;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68d272713d6706b93b9f14961c32c007b5a8627ec48c145996e8b50f1eff2914c82323b5dd4565b1c2a219e9516ad03e39d91ce7c57fb80ee58f97c9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98eec3fd9e1191c965218b3fc3b644da2134efef90754ef16990d45a75cba9bec20e1b3dfecf097a435d36063596dbaef012854aef9d4e89d23200df4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5368049f9d8898b096bf9542829371e3b67f428def2a6991745c98b18d2b943c56229a546b7782c77b76e75bf48f787904237d01b59bf9cf2b558ebb3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89078f9893c13f66cd4a261d315ffcf51f81ce477b427fe14e9d9bf36b652a99789d2b2c99c45e4ab3a209cb3b157c4fcf90cefd03115af55fb823090;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1ca93ac07123f657f9cfb8a856b2cea14b790f65fec2f219af2eba3cb6352846da5df595a512aae3e53a1a324987fbcdca34af93ff529197196e7029;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c21ce2125ea353cf35bff26b4c1c101c89e40d30a27cdec908d227bc5245705ce54a20530effd0479290dcf6d6459140f789af4b9e43dea0e524fc7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8742660be1abfbf0d8a8cd9feb048fba4776a8a72332c0b46918978cfbd2231c9943efadc9b14ca91d310afb5a4864ab00231827ebb74d6d293ff1459;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he18b2decd7e907b388c0e5bf1a839b5c13e765ed79187f875540bec3c625b694814d4b0a8d29ab8cd6873869ffab0ee590042c1b97d2b112619db1986;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbb13548a732ea00d878ab98485a9575216e26267669204836d67830532ea7bb210bd5587cfa26f86bfd0a11e2fac2e164643cbf9b35cb8fde7e49a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fb041bbbbe970f1d943caf872748d10c848f22630668e276d5f64b782322cce7340e72f3ea1b0fbf58abc8e267fc29e7439c35d08ef45b6644bf6b05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h118c777050a20507c89d2ab9a16b4013ce228de099a504daa6d8a20ee866bb9758aa47e1edff159ad2059cfc6faa0e9241055f8f5b0eb1bdc99b17c30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66b1ba542f2b6607632d0e209f05fc9d7055dec0ad131ebcc14a5d826a4b47e6665a24ddefa91427faab44b3e067c8e649af9862ab5e386ea630ffdc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f1d799555e5cb9c04523b55ac87e903a6d27817bf5f4bb56eb6704795bc7f089bd0148450d8e3cbf700bf979dd79f49a17677976d50c59aeb9f4a9c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15d623d149d645fa11170a54fa29563553eb8ccf786ed3de8081f0e44bacd7b4fab76e9af756345e171b640ecae462d036ba49bb4bbf8bd82f986b357;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h473ccc22adecc8071e15fd9afa765f72c9fdc78bc30d0264236b8f6e893d53a7bb34b23054c1473469b740a5f2471253deb6633e7d9f8fca965266b74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe8ce8ac1e568c65c64f477584fcaaae50c7b7aa2a5091fd25f35e96ffc88ac34da28c90b166ba601325bfc908c3958308336929cd3cf2ac1dbdad7f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb40325dddd7c68c87b06cfbb383996f7bdbf113ce3d5141439936b6ed64efb8270a6e3e8acdd75a8fcc05ad560af5352e403082fa7e665f01cbffcd7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64fb879e465d412251adb7361b03a7eeb80b4b8da24b16d363c089ef2e1482a885d9bdda57417dec3492970cd0f98292a7a9317da238be226bb37155b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h163faaacb66d14d57a430450720da0ab180f90757a71aa0982665782a75f079cadfe6ebc5f23938106004171c95e92003f3feb26726f2cba29bec1b4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6680913407be85625fdbf8ce38ff4481e9a8654f1be32ec79c06009567eb11cee5b89b16dc3c73de323ef5318afd7f6388125a100a123e21ffcf12d7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ecd5a428500fa015c9a392e9a983f5cde4d906ba51c2c1aba96fdd22920580530b106a693d6f7ddf006427b56bbf90fae7656e392816f8d5a9620812;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1778941cab1d2dbb2361d8bba2510cbd49a7c1f930b52775c4aeeb25fd214b494f97688f129659bf374869c07aa271d9ea3c0ad4e7a6017d610490b70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5601c24cf554222c64f661d145f585a0de5529cb5a9e43791c1d11400660b01267167815d9bbc1bda599527f5fa50fce0489204bb9a557aa07c11e1b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8803ef499e2afcc56ebb6104d60fbe2055985b4bf56e46dd758c36e1460f0087f4c1c4fa44733a13b18707924d99eb0114031da8265598bace9abeda3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c088e503f0fde83d89bf55cbb6091c2212d001ad87aca5b06c78548a938f0d5f187b019a1f7b68f780015c343a4f2d2b3f5234a223eb4fb2a6749439;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8e5450a426a6afb982b63900e4a830d2ec40446cd6fdf706f7acf3e6e45ff3a1118674b4497bd6a1a191315faf8496c343f383f7612fecd473611f78;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h387c9c1d7b0c85b2ed867bd8337c4ead5105abfacba360b621298d47646d5c2782b2a1cb45fd63deb41d0a179d816d1d17293347774fb9f6800ddb5fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedd9f1c2f41c05f44fab1e6e18a055b89e9802e426f527145013f93176b54716b89fb70b30a4437d0a3a4a37c220a203ece69c6f63d765ee10f9a8e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d66712abcca9b1a13779f670364e6d9399d7af5c296937ab66ada91b8cb2650af5f27f45ed80d0356a781f5350507fc70ee7166984bd3ffd6eba5e93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1c8cf17123ff7ab6a92eff9cf22b80bfe3eaa4a6d7d0ddc4089cfb49c782db8c6497bac9e41c5ab38e1831a3acf8ff78e7b04f634418aea477b01163;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a9a4960a616a4a82c52a6d2c8439b82e1536f2d421c9beb67b6e8b66fd3242daae616728404c66d5aab35c81a68c5df99720db7c250c0bfa9f8d5af7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he79db7206e07f0a350aab72168d6d593236b1079404790143f6c9bc85fdb748be348b028aa6dab8d10569ac0c32e995d12d4d8be1153e4a5e0f5e1662;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb4ec71fa8e022169e04b2d319d37a9476bb9883cea83eb7ef1b07e8a0b7520da15ea6ce58ca464ca01a4315228b6a31333ad62e5360365efee444c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1dba76db687a190574e93caca5e601c530d16266cc54ef4606403fa93a9a5af8b76366e27112f791b4616ea05e8a18f9b9b8cdd81b9fd6b6e601169b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17fee00bad955a768338415f838761a32b8f97f86cb0449d7cd62e76206108dcdf1d3384aba0661ec9d13071d0c05b13a32f71c61610da333c65385a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab2d9e97b7a27d9127ba3f5c0ac862a19539d44a94f6d680191d3787173196fe4d47335c6eadfa7acdf105ef16c8e70f316f6e1b339931d4b8bcaefab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7d6605ce32aacc3cb408238c90b37800cb70132bf719a194d2f11619d1687c3de810a65e02d1fa4cbd2e78b5bf8279a45a135c0b0e2039a6930df278;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43bb177b2610aeae528cc2e563549a25dafa27c8b6507aca6778a02ac1e3aba016c867e159e35b8dbc3e5f77c44058ff05010ffebcb53240ac2d1d0d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed84a61dbc476cc7b1c93fb2f62cb158a2314b4ec78a7f35aaa0c908824cda2af643de8f057bb2ed89aaeb0c6d637532481931cc67b2dc4bece64b075;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91eec264b289e273607147141e3a00ac5936ed4b6166f86a694447049528dc408912b322ccf21b4ceb4fc18b0d6c4dbc46f1b325a1546478a05f5237;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb188ea48e95084a78e9d7d789fa996d10cb1a0ba9afb44dffc29ee7c8261a07198992fc1e6f356a7cc8ba2076cd0ce96933e579827973863da79ef122;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3aca1ba95983bfa72b0d69aaa9e8540e4dfdc6ae435d6dbe21448a8d3faec858ea2daba5966f708b020bf57c062067973713c0a2cef6a143a321b98b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5793f7cdb7f23b32c783480a63b5cdaed39d58053e1729a807eb9c19983fd6e86411bd78105f4ede575665259d2c12e895a920e15b69de3466342e64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9ee18ff564996a85656fa07b98830cca66c1c717d76201919a9ebac0142340598fffa1d977ef4442c7cd2c3d2cd39a8fa68f5f7333f4c59a59ba4ed9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd1915c6ad3b139299455ec27236e044e04426d66f8b71bd7ea80cf7c32f1f5118e17edbad02f12e1ee3a8e5729f9c70d4140160b2cccb681ea1e6166;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b7ff207932fd88086affb9672f1851ec0f26cc4e6c5a69f2b2b34ab2e84e186e8410c2eb74e8947f7434777d174979da9241f9740247b7150d5fb267;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63d907cdc424fa619ba7949566f63bdfbae4b8876da6031dafecdb03e4f513fe77e3f02911c2dadb9d6d55655e1640e0efea6296103450d7b74ef52bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9cf6c66e925ef9f465c3751404bf1b959bea6e894931876c58ec93d6dd91884d8f93be331351383077e16856550af064c364ca4f9bea9b635ef210e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b9d81e71e38c18e21dba98420945e1bf84e0b62448512d3fed95294a48dfe0dcfd1b70c826c63a3183f700d451980e5bebab8d277a947fa2cf566a98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedc11c36ca7e1c70ea82d73d1d77fe52b3db1246ab3ee944d9a00f495753e98943f7c2c2bdd69a0e320db9aca4616af137770393b3988a846b67bc5a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15cd9a09dd85883a6f7f1b0167291f543d67b2aa27a7d5ef73fa50e176e81e2713ec857fe8df9304aef4de3b2fde531566e955dff3891ca790434dc93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc2d3111192c9fa02875f512829bcfc181c5376046a1d7256d0f0a4c0bfefba3e19fca557d65ea0bff85e0702e935c897e0a41c7368922b6fd1402d9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dd947bd2708053f5c588eeafa5fb30e6a48723b62bf8dbb4d795513b18f6ace95bcc8ba6a2e65ea6b503f2f587185cc0e68b4eb7a253562142a33a55;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5865fc164fff38ef286159ca825dcaa3b6089ae29a4adf023953104edca6fdf2b6336300958c21d5f104044e4a23885226b746e553ee06bdefd7b02d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94e36be35d0e23ebf57ae2d7da9513d72ed509320a818dbb5c4dafdbe0d97646bbe8fb99bfdc1663a598ba1331c591be8679968b61a7efc88603b66b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e44f42df705d79a83832383480d4063c57656799a5d996ccebc906d97925d962086e913abcb61d1defdbbd013e843dba46af5254c46bb5cda9a86467;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f06fa753f6a673a86bf3d012c76f44f2616d129be2b16e4aa0a341936fd5b207516fa569cbb2baa7d6416773ea4e9a4d1bd47969af96827759162d0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd57b90a2fbd821289ccd8c35b8ae5521f3c4a5c2c10ad3a55038ab3a69040b7ab179adf6fb80b3d893a6346e235eec7fdb21ac02a359eb7cdaab39507;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafe34ab6688a47d6283e1a2ab7e8c17c480138824e0b5a3642a5a085cd6485a046bb459042f12ddd18395211341e8233050b92541f85ba0fbf0e9b099;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19bb220c6e82f2dbc5972c6b633da2bcf08d489bb818ae05c078c1d373283999ae685ff342864c3a75568c53208d15c9c95f10227785da89e8236e998;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94c26079245f165136d43102b911745df924c0c7380d20c0e9f680967a26e8132868e0c8ce286629835d7b2362241794c5f6440949b61300039a4181f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb580cc49f6eb598f0ec92fd4d86d50e4f01aa2f339015d1076f8fe49db969211c9cc59c72cca88509caa1f5ab16ddb09ae4dc0e8486361aa3c94ba53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed13f9f1c6cb5819d1e0ef04322b2c13d4ae62831d55b5dc7664b6fc678c0f3b2ea8c370ba6f94ccbf7faa8cddbd0046db4f8e9c464c34b5f06162301;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc4a3f598689f33e2708159c00d4c25abfed1559b3bc5b1b552d01da97a587d695155e3d0b87d721ac4a041d4744124c93b9b0a50a284b3ac1b9092fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h563df4e7f6c8410091ae096923871e3ef37fe8f56d0c48bcfb08508239f52a890cc9b2e6656b25ff4a930647e456ab3dd2c442f48ec9b7e1f4f644bab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cf442a1d0ecbde93804391a5c6af6b1ca808f6d77706ff69171587c1b02b85cab712e41f76f0f6246506b7b00f651752a3347fdd4780470e47c44604;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e0165f5bfe1ec1bc176d54605cac5cc5ce8e945d0a3a42819ef29feaf670df4b900666c5f8a91f8eca1b3f88b80595db4e540323f7d21e824556822a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8be40927359e7127ac519a2dc7bdecb821a0283abcfc477e75309a4dd588e6b9fa76e9e41d87e8256e1a7ebc6b277b60c2e83370a033d360aa0fdb97c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4a45596ee771073d8c0188a9d739eca8ef6977851220c4902249ef770d1258885d2a92077461978016c725e5808fd1f03087bd30e2a5d95bd93bb8d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2acd292d30d4b6ae87cb2af82ad342b1ff7cd96d7d14c03303625ef605dde207ced0c411b086e071922229b345d83092463b04d29bae7f591eb0a0ef3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6af44987d88c642acece49b758bfdde906d604166c59f2d6d7905f08b4e8ac4930339b46410cf4c90d9bc21835694b9a9464cc9e6c3ed2ab17c7a6cc9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa208de56d3b3ae65b736f9bdb820c73054a7c493a8a8216f394988b7b836a8ca67ac7081f44357260bee45c600d756f957edaf826254b1e398bc09b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1360e6e9b2e74816acee371f0edb03d04ea7fb74b5d0ab784ac9b6bb89d3b28d53553051c7fb80beca3e1beb66f28f807de7ba6813d5a103763c578fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58be1cd1ed0b51eb9acf8a3a40fa69bf2b326f6a83073a2b950775d66b829f8bb930d13beaf79e4827d62aec9a47c5843d176d7f325dc81a5e1130974;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha07fe3fa15003892267a05d646fda9a6b280eff8e7381171ec4f12481406b8e19421f595ad1bfe3c5a768f689f5b8d4b030adc11ff3a2962d4ad787f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30937c4e61cb719003064e85917908d955674454b17654f595976137032dfb3c6599cf7499cca56672ee3bd321beed3fe26dc8c842db4900cea79c647;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27281ce3f5de44035d409d26c402a08825ba251809fa96b42e674128060dfc1ddcf2ea8c5fbf34ecbc59bd12187ff80a86b580eae38828d912a7c56b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed399411203004676c2d46350c70497521509cf5dd84d0208c3e7ed97b7ab051c157424dac147390d0f402b2788dc14144ec5817f8d72d11999b9d72e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3395880461bd121c5fb2d17ec67dc1fa0b6707b99218df1b95e9c05683d44713a1431dad08531fffa8faf631c1287a4427a4156d78a2d178cc7be84e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb644d760868590dea458b209d8258e65e3cf5a27a8c189308cfe5010d8ed46b5662bdd3c0b528437771ce58d9945fc1564e2096e978d12118b4a97284;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f4b54f7bcb0ca0a2fc8e17d42d5a533691572c49a613903b02a9aa37a9a3cdda71f37ac91d9ec122edee88656b8c876c99753bec3fa8514284f2d142;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h644fcd85948981f59bd61a352b00ddc170b33988b26fa5e76360d652d8371ebbf18df6d766ab093d55bae54d204a18bc6e60ea2d091deea8cec47d0a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b495ece587b49abe65ea9a9a268e0fe7866da2e22ef162f643b46a4a68b278d236ad2db64ba460b72e4d4d076bb7a50033f63882437d911a7c80c91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75f28a6d483e07c8167da45b5ca8b1606e045ce87409ac2b65032ea99247b5dde733904ef82745b2e9e20fe32359e8178b20e02cf7cde59dba9e61e30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14f8e6899e38829b7fbffe3e866ba671e2c692cc5451a995e041a0e0af5614b1170b6d6056902e9e75f16360c4ed4fd7e8b5545431727dc3754c98631;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53934fd3a417c1823b01ed725860932895df0ff8235641bce49d2c3a551595d24bbcf3cc5f46e2d31bca4e998cba8c8c22e35251f164b0888c0a90e05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54d390831d43e551a8a307d34454c03ad01998037cb83169f47aba4a045f11571d8f79c2cc69da8da1e6a4556ced4b4308e07c29621131ea216b7d980;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc49861ec3f7772934bfe81665b61df004a8688755eb6987e407be67793ad248ae036b07ee0da752606a361634eb9275231d6b1af4452885d87b0c1f60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5d812ab3fa2bf5e22af1e96fceb0300c0de117ec8db01335996b9ce9af5826d747a5444af51d7d0d4223033f49f85f9ede90dbbae3bf0056e9332067;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31d414adf50f5370a7db846f0b5db567e41f00294920664f7db219305e26e9c2361bc6fe1fd16833935c9bacdec872e21370e4780858f695d74398b4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3956c462a6d29b3bbb58a0c5ed4cb2d30bb4af7e253f59e4b884a1ca87670ab94d529532305a7501447745bb0dd25ec2e01e35a96421349572f21a39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb89dbc95b8d50dea39f46a553edd58d6b3183d770fd395d3d1da438643bddee3fe0a0ae184b76810a2f65bc81c3a209d5d8d547f5a88a6f16a6d47d9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94bdc67e91dd1194f3ec46cb0910548fdc3afed2dfb3b50ebf4a2851db9e92f1a86a856c2a8bfe2d613376a686f76cfd6f87e283e9d78552fe1babdec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55891a6029a604896a70e5f2897bbe30004217c98cfa7338d8565ba9c04a3e98af9dccf8e03ac731ed0a16a92aaad269258a6deaf799b0decc0c3cea8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h991d1aae7c5c06e566c02d7939dc7a8e1a20383e6f320bf05851cf709a87e7ef0f2c741e5efb9a9ab92d8f7017f282e9988c984b918c1e02eb1b52272;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51a07fec79e5e01e6c7af487c0543fef12c98c4eb3fd20c5f6e00f90c77323e499b572510fed90f636bbd04bba8aac480c422204ba3f02edd99ca789;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha49e3c0d1076d2413709ce01669754d7113787ec07e814f34ad7abb8c5c8b3311d328e490418832d7bc35961192802c3b5c580c69fb48b2ae12ce78be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc742f77c3a70f8d29d4ba2c2cf83a804ed28a72941859b7ea850a4b4273a1326f4d05f53e7a1449e1f7e62ad158d692c7e956896e763adebc5443c92f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3be371528c407b3c93b2a3c8cfbf965bf8c682af460b80cce2ca175c9d1d53bacf11ed8562ffc23cd726314e995ece3276103aea96208ecd7e095e39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h194c22302eaf828aceef48ec64ae72890ee040aa8c635492c0e08c96f8a60e9cc0759335b9b1a44069103ceb0e242bdccf6f6ac4bf0a53fa2fdd9cc95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58f2e6b3e315135b9bdffbea4ebc2638cfd634a3fe0a2dd5756afa5a50809f8f5be14b54ae5a1f8d31177d17db1fa0ed607fa4e96755ca3610666fb9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15b6072401630907f429cdba8b258d51640186c25f0dab6c117bb0ee26da269cef017248ff2ccb9f741734d2730ca9d81d2cd846131c2518c270e4c93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc439887866d8dbad635a0a128e3283b5d53a0b4f3e40fe33544ab69be4052287eaf375390d7e873669cb0a4993744c98af896c5d7176d530a36a3004;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d5e0c3fd2e32cced49ae234fd8facab4aa5a2c22ac941e512832efbd5eff7081bf81870a8a74ac85e3da3d6ca33aa4bb9c9043782f94d89392c1526e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4deac931b1a582bc27c84b07e2028daa30405838da8dd7a79509d5e63b8fae30e2cde8495182939699608fdb9b7765a0f4b5efd85ecc66357f50d9bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49f2991d33c10e44a21de31579e10f43bf99e743121b7bc37a5b4b39bf50d959cd8b8fb668bfcf0ba2df0492b0471230be350c279c3197544be759313;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b6ee0a715aaee44455481e9b8288f9ca99b438b3aa7c05114cf61acf6dc7199cb2b27b55793f9a340baba64dd6ac6d27d916aeb9cb4ef253d291eee4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h926d93052fbeea95a9936a15a1e4940f6e96dec09eeb8b22e51138314c797e2c1eb269f4ae941030f9fb67b40fcfe0806f3ea2039e98b3a6cca651fd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'head4ed9ab25e018628795c3b809f2bcbc5cb626a930063790fcc18a28eb1777682b331a3de269800cc5d34b273ac1752f003844acb5c4483a083b4ea6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cfde56622255b7d1d29fb4ccef309cd71a36dce52109fa6326c488cadb049bba71235d3ea3ddec36a90bdf685a481758f4a09979d4e488307662011e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e1ed0a4c7424a9c54fd3728c6d8c27595e92edf6cb6ea76dc9a0b24aab89de10d701e8cbe6d2f908cba80cc63f022ff38ff3c7321a82f069332505fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd28fb8b7b3852c023fcc4902b1ab1efa1d3b04d0759453d7a083b301bcd6e21b6aef36e02e884cdcda8cd3494d1c7b080c5fac85c5c8c9582eb8c70f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha866ecd4f1ffdbc64c8d2354504b69c89a4634c99e6b750dc1005927935b299691b1d457428daae669b70ed516c2011089fa3e816fba41d0c575ef976;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6faff08584a6be0cb7ef55ad5c24aa3ea3e00bd5771611d8b54740828a4b957493259fae1634cd6d5cba306ee7e4e5cb5dc465c6ff5aee1e4f0ff7418;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h346b850fe9cb19c69639064ea3a954dd6aad8d494fd340684bbce8938e19d0de97cadce79251d347cb3f7daace4b8cfa64b19a46e9175335ea8befdc7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he27bf7579dad20c95163349ba5bbfc8db18e9a4a0715e7aa7d26ad7f33c088a288332220749348760fe0f93905df14de86f51c87cd42aa05b899d7ff4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e649df2725526ca286065fdd45dd9c0d1f25e37108342dbcbf86722fbae99024beb8b87240fab21eebc325cfa90ac2374b9513853faaff1699c3ee79;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha172c526b22be5c39adf68e8b6de74f98f93333d06701b1c6066f4f01167425e45a69f335d6b64bf8840ec6601eaf97d9f3a9959e6d6c1da4d1ccd54b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he458b2bf3cba83b6a2ee737a16afcdcac1ceaf408909f9936b613b4f2746890b0be92bf9a1368a7ed043c0301bb870df7176cb013eb590e77663c3453;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc10bde6ab93beaaa6188fd49f31b33255bf6e09748f0157886a79a19c5dda38355dfd87f857749f82d51085141c2dc644fe4ccbbbcebe076e7eef01a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6356094d48fa0bbde33f6848654f0034a85b7dbbfced6fe43728ac5636687e83b949e7fb4a842bc40e6addfeb2357c147348818e71a6ba0214e5ff35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h327594a80195f31cc0564765c39cfeedf89b230162158877a13483fb78e9634990a136fe7636675f6ff5e87c9af83abbd70d2144d70abebcaaf38370b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63882e3f2395f78edd1a9ff2cb6a0a31fac8068ecaf991e3c2df34c1dde8e4a5fd4fc46de3d4835d6064ca7e9f1292ef5af5dbc42ce3d51b650a50501;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5afe2c274863bc0eff5ee0a04d9efaa7891b55bafe52acc1e0da6e4c6cd117d4292276bf96c850656cb65281fd8a986153ef62b80495d078c209c7dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h713adc14e217fb39bb63569010d62c75a72ac75ef0d81403aab20182b6e954eba77796b39e8c97cb5b8f4761d5b5ea5eeac931caac048b9fb963bcd22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h446d7ee4f939b0a8dc580041cd00ca4c5aa18541c0f0191cd4cb0840fbacd071f13281a618c3af823010b1b9c101bd0144f792bbc855fc2b4a78f2a62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf66bbbf6caeb914840cb7ffeddae0c76a3e87e97fb5afae57efc379ba242754dc360b28cc5a3c12b6c7878ec3ace5bf0920eb043d898ccdebd3a8c470;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h247729bb1557fdbda2e486704ae20559a8dd43afc58048f3d06708470786e57d3742982438a842ab8c292cb305e07e533b13d5cbd27a7b264433ae6d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he33b06805a60c0b4ef50cfd7b0246d262229090b62b25b4c538a67c7f4a261500daffdc0c016aa4814148da86c97ceddadf8edaee4c62da4b9b240456;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3479d217d661fe1fae80e6587008035d88ee9520dd4fe1c95cfa55a017e261a553a28dacacdfe1827029b28afd4665e849fa40d1aa54e890e64305d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd79b733ce626b922542f72e11b6421ea04f49b511ab7c66919bf9311cd41320cdcba1f4f28b94b95458ce7b4a4912142d6bb64c8ed53dbbbc1915232d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7afc0969266f9a7fd1fe0f129ed2af1f2736b6d29062df4a28be3ec458bf1af2ab143a5b8407839b63a82aa2a3e8456b20953d9b4cebd5cbddded8f38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35e8caee9ab7a185e3cdf85710a65526baf2bd30a0ce604ec81ca6fbab23183c36cc1c354524e9aacf82d9fa43d005b128222c3c54078106f9c4668f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda2e038df6843a2c0e21b8e88f6d71270af6cca8c6ed8e9eab4bf46153668e915c99a3d726c4c5af272a11944fdaa3a9efe579b7f6c095c1f190f421c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fbc4b7b96135a534dc380185d6f48d67caefe6b7161a84b188d75f867eb656ae8b23e95bf2e9c945e805c7bb77c81d184fb8574a513dc127a207e400;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9389fc5447536ae0c8969d32dd4adb81a97aeb85f23fee95943c13afa756888e9a4c8d931815826fc0e20468226851c28155d7b40c9b060b135b853dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dad22acf5acf373131620040abd44710c23633a9dd8c4de968a3d0575867ee1d62606e5d67002531d588fd0d2b33e8b03273c1fbd7d40def6440f02b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97bbca00939676954219f36b8ef9012c59696a7928c83d53dd45b44efe699380a561800ec49a3d8df7254268c6bf1ca9bc731bd985fd7e21813728802;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab12711cbcd631c441bea35dce2547182c34b2566f9f141d8810cfbaebf21eef1ffe25e61d29c90a9e1642e58bc1f12fcabef5d659051b60e28546503;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb64eafe256c5a5fa26cf21455df746ff78c89edc49513519cad515546f057b2ca594eb2f9956579c61068131e04572e55b4d93e1671e6a8c4b0651e4a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c208b3c2e02da2bc855188fcdabe0c255be409cdeedebfd9f1f00f9aaa3c7eb82cfda62d03d54c46da6e26749a60e4adc2eda1c2a3de9a98384dd82b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57f32b87a801d268251faa42fbfb6cf2190333e5dbd86c6dc5133da1fb572913e758f5674b47e3e99e2af4c62632c268b5b46d3730f7315ff7aa5b2cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heee05e9525128a5b7e3ad13e0fc10c363a4805cfc767c58e2a32d070136bc8d7d450843e45dde6825ac5b29c5eb62c92e2e84dc98e1ca82e6df73ab4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf3e9de16d04669bb596dc7e1f30f6561d5ecddb4a70c312efd6624ecc91a4a12699ea265b00be00ce10808e0e0dc6860028ed0831aba4958adebfae0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a6de14c9fa74a68924a154411502c6e2b738d37e0b19a011df69c6c0abb94dffaf8c8099582e262fbd91add36def3400cdd09d2ab9353d14cf952640;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9aaf58a9200ac729497a960491de81bdf6ef133c40250241b2621a50127c05f9581743562339cb80d7bf115614a00c8763f8592dd3eddc1436bad257;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he69157f43fa8b2bf3b155984e59c415c1931d1a9e4dceb7e4c51c1fb4cb4df32f62ea5cc71ac2c9941fc88e4a5149188e8da188b43c514fe69de13169;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd245dd73da535c86d1572a3649f9c99c41e4021ce7a37ac5bfe6ffe3e8e62fe5d9b1f538e663b4a7be548dcbdc9a8a123d9c3c0ab478353ae963331fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c014323f97a6968705aa0ed525e701a845ab43c8144f028081cce7220e864c9e1e26b864cd68491c8d2f1524b66b993225083d2a67ab025c21b25566;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf647994b8e3f2a45622b03766e96b595a10a5670bab90e11d1662884cf1b07de091b6567deec8792e3b68619aa315ea643e4c63a9f3ec0592508e5df;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h103b62cf84ada5cf18a3227b236dc8e9fb1db9076025143ddfeba1d7a62d0aab1aaf2137cd4408d06c9358101966eee6421daaa17a327c28daa21f3ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he91b8805008672afeea621811e0eef300a13c1443c470915c6439f7763ddf4906b058cfd4b4c2bc587faede4046fd94da6fcdb9c448996b25426f75e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2beec6c1f83f120cffde01c8af9c8d903759731c934e5ba37db9ef9175fa8ef3262d8b2f618b382b6dd9eec995e5807e46fd571672fad6b237c4a6cc9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c7b3a9de2cb2c378b740788b05cc5413777584d2f9fb559d8b4982a3a6e88dd771a9f49b3f39ffcc92a240c0234d01a3bb953155376241782b61b687;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7a529625c3765c101b06a9e7d6b412e34abfc8fe22f2b7b3d4310ae0d5ec8aed97d0ac4501b5bcce4989df89f25f1eeb70a3cb091926d44e3ca70d59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h748511a71afcd1c1422e80003657e4dfe0c7cc1e144e56edfd5d2b9398eca37d9f2f3733b681fc537ec27ce1dfeece96282c436adb67f241a68e3660b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d58054b92b1ff6d3f68ccaa426cd48405a23f23b7991f333f70100fa626f20ed9a7c29813caba2d74877bbb2d9a33b7d52194a1f9dae13b418abf48d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha33fede847eb5cc525b3c28bea71ec2bc20d8a1586d491841bfe65131cb421b6fcc72b2e067c80937ae82b005851d80e7236f66817e6252203a4b81d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7253262015a5ecc64b66bbc15c7054cf3fa02f0559ed3a7e6b53b9e5fa833a8b52a8cfdc3619ee8337cb6c8bbb48218411d32d871e06f9aa26fd264c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc438c7b21a463262a18ee8227008377319cd9a4b37000764e6ceb04ec33f1825986634f6f1b38b47b19a9c0fb88da5812f420138a4a71a1d0eafa6ba9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h330d590284a6a0a0fa29c4e1e531a6fdeddde8d64da2becfa4bbbffed3b50577704e0b2d35cf894036cba48910f5b6bd2ebf50e340779910af4acc671;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37d84efc5f16a46ce8d763c87d8d3d1d1f9ba437d454b7131c0c0cef7f5eba879aec20dd8af2d348a1bfa7e4ad106df29256a821819f05f48066ee4f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e1b0a5ab5b6cdfe679f9af58a65432c53fd938a90ac584d103bf47e555ee23327f983ac3ac33f1d611be8a8bd781f76c7930be17061b76609766dca5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebde84875dd403142432f520424390deba2a330cc7fefc09fbf1d7db4120b1ca95108c0a34ba629a7d047fe471acfa88c92bbec72ac00268f1fa3262f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7d9284501d3738f53e809594e55467f008ab21bda31463f8a57c53222d83169f26882f05dfad2f806c5785e9c7d58ee2a8ae29e8643896e51ba5a7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d3355c2506528b87f1ac3a27a5fcfdeb31ff82c6689abe47815b980dd9a4f9218f4dcabaa84b5a8a1ab896cf9c57778b770f7db4823c8807f81aeb85;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedc08d8350d58c5f7589a956118ac752a12b789c2b0b41c2c795685c3449b67b16269a706d9e15e97a03b835e8a139c7b52155cf301b75347a43ec77e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3be0f2a5bc9197fafbb5d6948fff391a13b75f81b5e8608270b6e3b23738418e64f365f2c163fc489efeb18bfd92163752b62b0c01898a1bd628475cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36615889f5b7598c8f10522cc78e012a3f8616b0c21241987d727aeca951243b419891805a326c4826ed2109448d08489f0368b2068c5d1be9d18cd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h309b2cabf5c4fa762f162b1af3b908f29c9b30d7ddc17de40f88ecb86a0bfb73fac6cf9234beed18ee41ab0598b6ab1cf27dd5ffa351a6faa3268b149;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7eeeeac0b04e0529645a00c3650be8708f59609185cef954c04576e5f20b6de5132f11d993a6442586dfc929d6aba87b7977cef30bcd58dd9e3f6ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b13701f8f1caa8f0315842028564b9d2a6cfbba9778697b6f0d0971978fb0607b9015ff677519bf338735bda4d269d8aa8dc8c15ff37f3933cd3e05f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf0de5836884c0545648061362608532e40ddb29d0b1e2fa1900e7ab6b8da90c5ac57566f42a48ba7dbcd4695fe71ed241e0767d8c482a0d0c2c48b75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bdab73d26237871f164f5896909b79416abb2c3c3dff5fdbc0f0fc78c4e164b8e937d004623ba97fd61a5ce268744502ea93bcfae08e04064ffa5067;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91953ab73fd0c8f981ddb4a46c79d2fcb35c4d8c12e60116d67243f7bda76144b5814f4229a68cad9a09214978c876f66c922d55bccc94a45c73c9684;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44ffd4454657ea5812ff3ad9cd15fdd96549847640d7b8b79bc22a7fa69f7123b93d370b7aac4aed12038698bf060284756e188757f17ba6d487d1f18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93f61c836cd2b7d1d4498001e1834fccbb84691395afece5e6d4c452bfb61090cc6c0960ca528bb4985289b7597e5f6b8634a6fe2d098680235957e69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd46576ca937cf62ab01d0a31b8f1c309cd39344b65b30f1d37615c665b82ead138e73e6d2e125aa97e5773e272f99c80e99a6aea8a12b49cbbff4a39e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7bd6369b811da019044f580475e243687fc46a39efdccc0ec2c7c08eb7ba583d14beb4db75c4d8737ea3a9b807a6285743ae7cf1d723e3bff0d8e786;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed2bcfd626a06c78c4875a5bf4b29980ac8033a324e39459fc5beb6c7de996d5b28c10b68bbaaa276b1318a697ff8197d0daaac23d628dc8ddf18bde1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebe5ee4994a8416d238b8780f6dda3f9c80cf18b2ffb39aa28a16eb108730d6ad04f01fb54247483322acd91495b1ceba8948d055a1fe55005f7a17a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78e413b26a2cdc2b26243c81d81fcbd65445da554afd685e64973474438126d24a3dfd5ca66f8a2a0933be3307fd477f66516bf8d50a89321940218c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb113923e6367d4444a53d4ef2fcd135ba3c38da5ab4cd1590fc44a5bbc355ddc1f2441b249e412aa8061055ce33baca5a7071253b1ab85d5e865ea7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed676151fce05a2617ca0a18838107ed983dc8e6a7e2eb8a354610e8df2ec07be269c1d7ac22a766de3ed8e96e5c4952818dbb9e21064fbad61de530c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h712bdab96e8feb553259b70ff2222210ceaf070dc5941dfb091214fc24d37eb79f3093e6490ed5a1944f1ab32fdda55e8a6b670f902ad7fe82e671e97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e90d176874440bb3fe301847c4a57f24e4a2043cd563a7379d63873368d22d52553fbbaf59538d2018ca3b78d2c798439c4e22ef7dc06f5156279ca1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcac3816785a6f5c72379b8fe82672f05c989864e8d79b3d9e58253157f4f849b4948ce2c3a3b0bc774e6bb23280907476d5d66b189a46fff62c4ebf81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88eb1c7141350d7635369e67260a426a5e2f6a503cd0d29ea244a7eb4f2a917591d34ebec27cf1bb0953540469ae0cc7ac84b25d0bcd3919c5ba9ba6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89a8991b5665cc19f44a7c4a02bdc56c75b0559e722a69a64d8d5ad68d7b981d21a00e774c9f852efbf5c225c3319c7f9e467dc39b4ab86367d28b008;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd79f4f44dab6ed1ef898e8b939359f095505f0f45155bce2896929f7f4007c4c1b7b35118374a4de4fe56e9bf69fc488cafa084118df2bef44f0c70ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff806260e4935d6b0757f2925fe458ee3988d277ef61fbacf8788ee61fdf08163a21efa0a56a604fd5de877da29c235dfe26abf240f4f661e558c9ea3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h576b55abeeeb1fc3b3eab8ff55737b5f85953be3037945a83fb82c0d70ee2b6078f1f974abd63a95e2c783abb811a49009f9b043436c97cd0741d8a54;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e1991f7902fdbfe3a2ad7d3ee2f309cae1ef745df5f6a5f8a31f7552cedb7aa42a79323e8d4253c7e96d94d4d06fa89d6920e79dc06441dfb6805832;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf53d5a51ad25b342350d70bc79ab2743ddcf4544a566ba829534c91e217b7133b6f55d17f4b9299237ff1aab9b29fcdaa89731a875dae859b437e27e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9579b08d60dd3260ade582f5a2ecdbb453acf2c36d739c542cf162178b86efd84fe9ed1f224f76824f5fe466ed3a51ef2d93793dd7db5613242abae51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee04f7752d3f1a383d2bf2ab5662dd844a096fb63965afe64147ada9d143535826606abb86cc00993d41ad42cc313528d155f01c43efcfc078a2929b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fe23453a3863d996f9b3f038ba6e81f6a60474389b5aed4883ae699e125af158ff5cb9b9f651dd8b7cf700c0fcd720f13163b3f15723071b995d5ea3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85e7e073bd9ff0ae0a366b30f31809e01dbb1b1321cac63bc72680a71839d4023182086473743eb959d18ff92b85e4156af222f73ed394c61206e21f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45245a142a12458a554799441a6bd2b3c5b69da71788b3ec0cba0729394b8361f09b53f649ac517a77bc862fdfcf497d4e91ad424452cd880344aec63;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcffc7375948fb072c28eed4599938d688611083d1d101a896554dc433828228463fcb81dc0df6b07726d23747f84e95b8267f7cbb22d698747b3d1542;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h906ed951b293dfd80750186b0fa5803c9467988723e1184ba1c1d3cab8d987c55bef678a582b8e4f023e65b7eeb6c596c17894c49190e2c7aa9330b14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6210acecf370a455dbffb93dfe66dc1bee234b84d5770fd513ce07e1b258798e07d6311a8d0cb1c388974cfaab39b55cda027cdcbf7374e22afe73f7e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5ec3cd84d49034c052a358a365a20cfc7ca0713a7eff8285c0303daf9d03fca8053ec34fca52923d1e2c1211473ac0506b0901bed2e0b62e365f4774;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43375e9c92520f1ce55db35e56267f9ad0af36a2cb8ec75ecb7c988805adc8003f2ed170847f41519a298b348bd82aa6360d2df71628e2600ed6324a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h581e3dd1c0ebedd5e1ab908f3ca0df1026f5200532bccf22e95adc53d7f9c2b127e3a13ee9002d0201bf9020e3dd4db45785ad470838d0fae0ec35e76;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbbbeeb53c524a1ae95c2c23d8edac1f7d396ff790a6da0039270335cf2fc00c9f56832a843f51a8a80aad3b471c3fa6a77f2a52e51c3273172d957f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he878cfd2cff91e5bb5ea7d4452765965ffef35d902ae9905988bedb3575dff864a7da2c37405334c2d42d3d20beecd821f845c3ce48f966df80d47968;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5892cee2143d3bba0b18cd50cb6078bb11bbf2327b72af1eada419e0eadc5dd0847b413cdab1c40cd4b3ab8bc98facfc579478c194320dab82d86bc1e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h433314b7bc2514aedb7bf937300202758fe1088219cad31d6c57f85593ccdcc3ee5cc92e560b120145919506744324585d6ee156d57be2dac1c293fa4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8113c173ea4913b879b12fa7db8c7033a9e2f8e79d97dff187c19ad8409e3d7c79d46131205e04acb85ea51d8524502a30abfef415d39098dcc9302fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he07144bcf135d07450af0356fb30223364f2ca76793a33401c82e6ec98952d41d1f7b55c3b3403326a0d9f7d4d1af6d9eecbd51b2bcd24b6e0ec4f58f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3887a06dd1e02e541506b63ede2c269bcb8612451deafc7b2f1b586f47564d882b0fd226ebb28795ef8a9ea9ae799427fb7321ec6ae3c106efbd43dfe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h629de954b10823260034307330141b3f20d4d66d660f634fa05a566edc1f0c6c4e5c442c7e9c49811455363b338174b936a19c6bbff1ebb336a66647f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4439617eace86cc32ce7d5c505fdfc97fa8bbc350d6eeecc69cc586b8cbd361dcb9f5d89e5024bead83270b1547ab220a1497eb94045dd55091de9ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h451568f4ce5ae3e4c18a37be8e5d7b472e8d9f863ef90c832debbf4c037ca5080fd5a5b5f5ab712282b1eb5b7dbfbc1997e0f569d9ab826fc4cd39fd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h933fb36f09d279f938426c2ba71ff87b9bde6753d6e34e35d8f2b9785d3fe87e38e3e6391a55ddc418f12db7106d93c0b1301a26b50a32a90eb0136ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fb29e55549cf24217ffedd4f70b4c3073832c61728e54383c2a086678abf045c525588ade232ddcf6e6cae10491de0f8e58a4a290306e2d56d373707;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8c3f570bec5ecfaf3e915b4afe56fbcc42e7e7ad04000a98b2dd2690d14f59f9257b76a15ccfff5dc945af854645062232164056035d840cb2dcc236;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24197e89d1fab34e6df94d738148fcb62266ddb8a9d407400c152bf09705055a7579a236f2c95cee1fb4c0fd1051f7f4e29d6a68abd06057b90c266a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8f7735253fd32a817c5385bad1d74fd41b410b2695d8c0bef4b5f7dd1f8981fae94b68c0f5edd818c89f83b29b1002446bbded6b65079da4d7e4baf3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a23af98b54e73e2279bf75f9b24e7b28db0b5720d8e75b4efc035f1f34621f541fe1284a8cc4b495b534d4ce3e5f55f6f2f80a09c56175cfa0172c89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0b5e8f3ffe1448e47ae5242cb54e76be3e5833c5a5ff46e234eafab5d8d76cb54275d2cd64b579425b339df7e52460c38d86d6fedbcdba9005e84fe1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7ecad5970aaae4e3be6bdbe1f0499eb337621aae701302687e329130c0159d4fc277aaa2ab2d10dded21f75b5e10d265b965da3ec3de50f0444e47c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae39259c5941597fa27e3d35506fdcf1574b7aacc73df9cf056ceeb8dafaced5d6b5a06eb7a38afcf315516c555c025d5dfd80d6c10ff62d9f96c083b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb85f3f7e19f58a85290a2267552e959a9e8e35fd8497b3d7b93ad3bd9d6aec553e15e5343b773d9bbd200b669c12ce6c40b59d1b0860ab89a1d012873;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc43c84ef957603ac2ba34d796fb13a0cdedd43d9ce55aa7cbe94912aefc172834e1846988610fa62e390d632074ff177ff554f01c8e31a0bab480f61a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a89f300f4f28ad36bfed4e6478300cddc939c06783374d5a0139219d8a35fd4cb1e31bd014b0b2d4583ba304a53d8e1de163e121a263e554d68da156;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92808e7af10a1b62046e25fbdf5fa113efac972851beb0dc33817f367094b8cfeff5d0a3c31aeb92cc72c33501bc63ad375c6bc8ed3c30cd48fbe01e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5278260ddd53cbe91cb5cfbbdeb81d0362f5865c7685359d90ea95a20304d009aa222e1002a40a31ad14337775b1bd7c5cf8efcb64d80cf505dd24c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4401cb466463abe7713796cf1ea23ccaf23828d892e0169b9db34d7494f497e0610393c235be034873c94bae741879fad17d8bbef15403baa277fc63;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4f06b487050863551844cf475eb7ee766c37eccbdf23120bd56d8310048784e63efdc988775384ac9149639a314f6c6a96b7fc5baeaf8d550f733bfe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bf108b06d4c840eff4e456ac25bb0fac9134262a4f985da65a22e2557920cc183f155d859a35ecfadc89bb4fc72057012ed10eeb4a1a21e7f611b32f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c27200194888698d28eece46813245e8cfa8d6872f7b1afabe8c8cda8f1c0403e244bd688f502c81f157684b5569012c0f3f7c2577882d2aadee582e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5668ecdca667552f4089042518280e2db68938bed169524c7f08356a01dfbb2ad785f18a75e1f8eea7fde7b5a70204bd0de6b3d4cfd2943db5b9ae292;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5c0db2ce2dc4f1c43e8c744075a4ec2852a83de4d03199fd8cbe564aeb896a8184d49c9582b77c2492385b6ef8e2cb1e5d2995386207799606a19aab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd19dec3a616bf4c84a99411ae2d876c0c3fba864343b24c87208ede17eb91f6744aefbef547212a8ecdf7130664afe37d704de96314b0c824ab30e56f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f248fc4d85f2b691d2bf123f7452fd3214881dbf0e397af4eab37747bcb546669bd78fba5bb922d68baee6acaf9d3972c120d1b3987da481c28e1c02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h434dcc5f2ab5d4eccaf4d4ef7304875efc1512aebf59fa574d274f5a7d6b5c86684e682dd7b75e55ac9f0585a9efecad3771585bd7d146bfb30a442bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28969b3ca345f784bc6188f03a5b700ff2218acf858c7ed09adecd36df427ca7575efe5624861ca8c7e5c56ea4cb29fc65a158b27c21ee2259baabf5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc789d60831fc93ff82b5ead36c43d9bfb64302ab33143045f9161d3b02ca9e761e073f4983ed55e6b36a83ebe029d6cda50572ff570bc67fb5cce85e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77edffa3b1d65362e01c98cc7609d61d4650efcc53c27bb719755134166274a8e3e20d80cfb30dd0533df69b74fc40775ff14f8c7dca41254bc65ec83;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b3659bc0f1d5877ac946d77a7e17172fae4fcfe338c4ef32f2024180533c315e7ffb9108b1a30d40a737cefa6c7c600f27ea29869120403e9b581ee4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62859ac5ed16fd672384d76b38e8259b6431617d1e26b54d197185628627567a2cd68dab42c9b85cffc027a531fb6e3f5218bdd6d0bae96c136f9bd8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3ed1b1fe12f1b4e9fc5304c81667b601653a45745f37291fcca22cdebdbe3ad1831d868d1572b2b883490c07e75f601d2fd9ae143f55184fcc5369be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ff8b27be279d8d7bb50b490dbc139f7657712fa1e1094c77470ee61f3179b41b83ce3647e92fedc170d51f5633f4590a1d593e369dc9c0e806a664a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ba97be439cc4112562832bac4779e005e4bb9f710cc0c273551e8f5111a0b88ade16002725430e035be26a4f472ee87660ae36119f283960e59caa12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bfd63b17b06f75bfa370968ac5301fe76e1794a34c181faeb177322fce7a2ab4eccaf625353b2b5d5662c39df8626186187da669c901d5a37a7f4103;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcafea7948a3611095bc5397174c6d066dc371e0def578ae8ecc0194fbbeaa118aa564431ccea74bd62738c1d105057a099275c7db78a1ac99446c860b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ee546792c71d85ea8f47a0ac2f1656837308247bbed0a55f20580f7c93cf07edbde33e8112a3d700d6fba37ddead959c0167e08020f34fb5319d4435;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7927c395f9803788dd4e0140951bc10872495c6bb305902060392404ef019ad163a2d55043c8c6669ab8bb69a635ba3d5f34998bed4169cedd54064a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f5a01d9f11a0d0dd9525a76d47e573688acc8eb477fa543ce6fc74d02ba3a4b9fa7addeae82c49707b6d3b44bd5a0b8a666ef32c67b4e53b5fcf8dac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb5840a772b13ffd29c61574eb03913c04b99c93ee7b9933ea00ce04633d23c20517cb8f1039d4b8b971e0d3a2d8da11a2faaec2109f46e542a9d1992;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58c97daf30e620bf5d415d84d2ad319eb7f3d9b1a9b9dcb4bbb6386a632ee142f9f94d46b3e6af1337bc5c3421f2f249e284fa8f1af18e210085596d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2959a5328113f265d126661b6e5c8d470eb840ea8e2116e711debe2999fe0585be87c7ca0a6e2f0639a62c64f3e0780cd8926e211e4282094f7271ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha14346a188813520c4cd5ab92d5c0c3c92b7c9d3380aed881b8458d7c687d21a11e89bde264134a4913a21e423a5dc04075910c239316a4f726c1a850;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b635e766c156c49ff7d95adae0eaf9507e9b5812331fd665a2d02c960887ac7668c9d62d49b6c34ebb3b9aa6436bf8bf38894ac70d8b9648b15668c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcbcf8cc7b8e4f561844567afb96fb15dcd120fe5ec22f22eebb0ffb11309f41be8635a6773f33b829ebf794cc3bad441289022ff48cacf7ced2e2df0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cc5934ef1f901d70e67c0e58e3f8e426d615b2b5eb5b3a25c599f26d9192531e2c546264fc158087a8a31cda81ed67b1cda6fcd88665fb4ebeb29d76;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd47403a951d9519b329f982c00c929b24b9c09e4ade9522fa71dc83eadc22b02fc658185dc0add914d0879fcb9f278be6e250ec21b6b5ec5c274e7da5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc29596fcaf6d6e1d206d804d843f4dbf79cbfac5ec86340f267e7bf4a0b66f00a83b7571c8fd5f062bfb4858228a63bd95cd185cf60f5e78407dcd14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb55b29cf1b774ed5f222c429a5a2fec41560cf7cff96b50291933d70b9da2859c4c42d179b50da7834e9ba27a0b50d1bfc1cec6300b8733fa0b243054;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7377d97674aeb69643e7c175fba2c076e072fdee2be505c812bfef8047215edb8308b18b2b06e47f0def8b01e4b9ed58467b806036512d9b1bbf72b77;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdab48b6ddce0d0d70254c505018e955a6385c30ad01b51320b03025b8e2c5b178897d4f26cde07661a47c7e9a84cdf6c305cc1c4e6bd9115d928dcb58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20bf52b208773eacdd75b1f98bb8afed09f6b4f993006ccc3ca6b3886e3040d6c4fd2fe45c7364cf8575e3c15d0e6961cc786011684ed1a3e960aacad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc40e7916ffed1c1846291e4c996f838d5430615b46f08364750ec1214bdc36d53246a1f09024fea1ea71b2e57caf69818e36a5c1b3906571f44e1533a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7db5ad1003808c43d6dbcf4259df2750d36c0b09f390c25ed9b5ef6d702d12f64dd1ed51b9ba009955c18f81e573b540d6d3ab9c03a3034c3beebda42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8020e47d7b3930e69fd90729a97ec8cec006614aac212b323ad47e5acdbe609b873ef10a5c83f97f74dc060592492d939531631355dd487a3ecdf6837;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30e59ecd569395b88cb77356779f9696a0d6bb5eb410526be620843c3fce2c6cfbad04c3f4f039ac52c995eef57f1c8245de800dbf2db6156f090bfe7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4ed75dec0f724e3d27adaec5ee07c473b869351335da507c2a0669c133bcda35fd95d4d1d7627f2f018e2b97a4ff8378a2e647fcae2dbcb7343b7e05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1caacd67c9977b80894e376f4f5fbe4897db683f39474e777c2716c1b62541c915705abf4734dec0d80cb6742cd03edc07dbd10a6826c2ecd763310c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9745b50f39abd90a74d1abbafdae030554094150c7f0f9fc1c651510179d5fca48a05f682940258d31182b942641f826d29c9f124c37089417f8caf20;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b8a2acc73d1f2f194fc246af0462b6036f3ef84022c24a1cb963cb95dd651daee7543362c49d2300b52a14318f63c512e8aaf6903f080643336889f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he84ffcafdf9efdf5357333d31efcc42024bb0db2ead4111cb63fbfa1d9a08c6ffb5b1734a1c92fadd05424d4199b60d5bcbaadee7ca8b8333ead736d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15047518afe1cbd3bcb2264aca642ddcad455b969116e020d186abc7b494a8b8341450158bb918371e265cdb68bdd0f98cf576a8d1c344f09c1f1a8a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6077a160aa9f88541ad101a198ce935b5a9f20dd7fe15a8d5c34f3a315168cecfd8004ffc570aec1cfad62f7900ccca5146425789d3de2cc45574c34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d758d12b8c6a5dd2853c1ff93b78004cff195e91b02edd744241d71b7755b8655877f8aa2c7e28ca5ce17030ccf6636b2cd05c34b9aaa89dd230c116;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h492b6b40b45db93e269768f1464df89abf130b2120d4c04f02ed4257d1f788e607906deb64daf88bfa7b6c267dd74f2a0b88d535e3fca93889d69a38e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb90e6ca9e1d8406245b22ef92053fda678889c658aa75e3eb81b77da8d061493bd4c660de2f38fe08024d43cd6e869926331c5729fc652f7295b8838;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab10dc851c6252334f5644cb0b540908a5f6559322043fa6f084fca9154c40bd61b2bb42abfcb78dde4bf72b1b3ddce1ed8cc72bf2f0d36ce93b1ff48;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec6997f5df48a91a40d482d2278547ae58214861958297a17696d4856e3e88fba1cdb5fd8395ff7fe537fc74ead954cef8a989e15782d0b18e6822023;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd810f9d53d2c7d5a2b6ee05aeef4a1e07386c30e50023ad62581352590949611d2241e77d401f29f5e41c2c4c77729d5cf10bdf387cafe1f97bcc066a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4be09383a4dbcad36fdb9ea5b94334ec601f303f55dea2ca1d48603eaf792c93e97989716238583c66ddb5ce740ed003078038f36b1d218b40abcdc0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86e36405a4cd8c57f3e1c42995d1a4ef39c66a6b6b3fa890207d203757f9cb648febcc301d0ac300e7f22a3c561a726e7b2ba8059d7dec0242b691adb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80110852c09b5b0e22723d96509f787ccc1c0ed810e334b87ecd88708f084c755610adfacf9b3476266ac0b3314c2bc464ada9c19531f2e45908bfbeb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cfa64168f2de66d419e718aa9f2c4a23560dff3a057a764592dc1bb67d3f20cf3da08c64ce063877ba951149491ee73a7634d667e5d31ee77c19db35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd13208d0d5ab943c9df3ba97773fd59ef7986219426e2a987288b7366652c7056b882efb9436a0d5c25d024da3ee5f32da6a63d5e88255559b784278c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c4cfc061b6e72bd2c370f1b07519129d337cc1278dc05b9811a04f40b431d1cbd726050f151af4091d1db269dfbd2c63cb99f11ddc064307fc1f86a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38f6a58898a14e50f0bf1d9b0f86da68dea5910406805de22ea9350845bb9cb43c8a28602207f3c326590d40c59196ebd99054f517166984afa870666;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h203841b1c29351a6730507f560a2151724d2a9d7381808751180003cf5e00d387de87610ee3cd99a43d502b2cfac2ccd3f1defd19b05ea2becec74583;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd976524c7ba6372f6d8f72eda804928a46d8a4690274a039b818b56fcf5904a589573d6625f9e2b135e9329655bda347c66cee82db28301e34002bb01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcede58129e0eef3a771684ffad810eb7e5c7c21fc27bd807c892a0be2ccbc52730abb3a0e080a5c14946ac75df751504f116d0e8cb6369f0b65f9d76;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc22bc2e20559da7691f30f57898f0465246f21171e4ee8a3008c60191e92a7349a7cb543441f9d30fba537c9d825284da4d2ca0bfb2f2116e0b8606e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc16e29e76e90fc0399276abd81af2acd90e70112b0a0c361cac74f5b267a91d32bec97816d13de923d4d6d6b675f42ca06c8ab1a421744c358d0dbac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfde0744da42b025dc1b325ff5d29b988cb1b2b16665c94966fd0eeb1e4734ef1666d53acf2bba40002cde67aeec6ade00beb9837cedff1df0b8a7fa4f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64248129baca85eaea29422feda75ab208d5b4660ca83d94db373392b3638ab36bb4a66a2fe22a2d58ff53a9db8c9d233d22e4395cf8d4c6f6693a16f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4e969b3709575b8b9022304aa32fd929623765157c959cc5bc21e209b4d6870c605ce86f359c1f7cd8106ec3dc1542740d2b23b18182e3c2c4d9755d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4030f5b011c243b329064041c898d7be4ac4ab444d35712d31879de522459dc98c3260b29a7d0d606f66def379d1965f7cd0551c39dedfe591b29a2a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0fcc67156c0ad7735b159cc46d27972a87cffea9ef69e3b6f2c29103ccf9b8d90fb21d82baddec6c08b9641bae26ad9905d8d5c11d09efb800ab66d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae17eb74a5b72bd533257d8d581609de3a3266ed6f7ca474358ac246c861fbc836fa983f48950d716d9799ba2f73647305373a31458f333f5eb007708;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3076d6af51f4939daf868370e9984aaa8d3fabcd08108d2db5bfbde216da89e45d407d4a24b4c992ed08e89271cc0b0e086c9790577a1be83226c32f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc91f1d412434a5b0d15369dc75b6d6009cb74a4e84a642ce4190850da8df2c902d814b3f1e8d1d022a52ac998fc6c8a42ffe2accba9cf45a739be8860;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc140f7ae6104ca8a6746dd8c84791140aeab4792810bf48ef7de2c6521cd26cd4f8f369e5d8a15067d06d9b7d8664d53160e21f64e17a704520938cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8a14bfe51df450de6f639b59071d46a3dccb54efe08c649e3239d8fef75e2f12bc5b48b3b761eaf7b83cfdd09a55ac9f4c7f2c5fc4e3c77818e11928;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he002b11ec434cc02993d9fc72acef507c017b1eb4b23100aa4ff42e1821c684ff2007b52ebd3e5863165a382fb1f317519ca6a433f24da068ce04bd65;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a44b83740f17c31d6b7a958f4ad2f06bf71d3673cac16f3ffaa2f58fdc913917e97b3bf47c404551d18fe1c24799353d0ea47756dd684d7b55d2f075;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e7529b18e6814c19da6c485b025a1e88931f781123e7a1f17bda6611e42c23dd6f3294c523425a63b52d939560cf7a765f5a0a3726a91cff6d519aae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h869b416d16b5f6b6377ebe2dbd896000acdc39b8c87b6d120ddb420499313f57a39beb83053358deb8dc54ff1f4c3e8dc4fe812da2c44a47b9dbc867b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ac03aa68ef3325b25c4cabab2851113d5574798e3d972c5a9a0a9f074846cf7de7f301076e44dff5991afec65149cd69e41d7f567dddadbfa88a8163;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a5e32f1a65da54f912e6fa4894ae623c42457c2b2f09869abc799aea2d7b3a57f9fcaa2978c1d3dc227815868c0eccbb4e73030ab3629ce602cab338;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c8cd3321f4dd648252f621c97273f3d21a6cea52a57f856b0e9af610c73281f81024c790fee57e536d835de5dd4261956cd32445a02e719ea41a347;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7648d5e1f070d349cbcfb77ba9169022f18fd07904334b4d048c3a08217750525fb0985ffd1750dc2c3cb8f51959134e41e7997589fdf46cae9b2e2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42c8d19a8786e0981303e5b28f4d0a806574d2eed18bba615d7e5790a4ede2eeeb006ae9779bff34e463b1e1d23c2187f0209cd6da228ccbefcd1107a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74d5101a5807c652e9fffa282db4dbfe0dab4b19a64a8cc6fd52f46927e7ec74a87e025cfe03e48a7d27b00b56db2b1b4d77355828de8b826d8128a16;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5126751b3367829ade13ea9e3a4d79dc8c7a2d19895848a06e2bab5aa4eeafbd466fa3ca611ece2fd9fbe93460e1264c4811abd6aeaad6325ae98954;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5d30111d896bf860b82504c669d88a14a4007e8e72fb69de908cc4154c59ab0028d26ae4058e12733ad21d54fd2079f42e9bb01edd48618bb1f566ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h163115f7a5617c1eb71b051f43f4ecda3f7be2b7a2aae18c36a96738fc2c7e4b5999ee4886f67a5bc5b997a7525b4fe6b876cb657e15b8f5a485b3dc0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c2e22006e0b16dd01e80f97b6713eb7cc8b442147682a45832736a1530c8c354e207142ec8fabc688b7a19174c020776582118e5a1562b70ff30111a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h132787d39051b8caa75ba1fadd38d10bd048ac186eb4a91662d49bbf40492be193b3c15daf789e068bbf063808c18668096ca1f1f2b1b6f6c882481b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d5de7ae801f82200588a10fdc8793556698ce417eb35b9a7cfc6a5fd615495518ebcc0c0068f01289d662a83bc99cc8616f268821ccf060b19148030;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53bd7df001f28461a056e5f6da6c234565363326d792b706bfd16006bf0e7835fdf5a8274ec6dec7e608854c0ce9e86227073a277de75d30b4d0a0a13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he52352d9f204553fe8873bfc79fe209327d7fd7ad2a49f859058d3a30bace5af5a572581e11a0b80aeb8155ae9d915c9a0cf89bc8eb491fcc6a68082e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf35ed68efe251b4ba25242fb5bf4008d35b9f5aec1b1167fcc76ac2807e50d5f2e538d326ddfa8182ebf72166c14bd44f1f34f03461ed83725aafb024;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h438d2b416379cf9bd7218c71df008e0617e402f4489b35f23bb3304718ecfb4ca8a160fbc7942ce4e9004b120a4ea1b23bd7be0eacbe7071efa6e7cc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6c86091355f97e1ad6f0c58fff0d076b4584d1c94204ba1f8b10cb5c088c3e6c192886467e0058704ef0e1865974b93b55b237f462a1cfd47d4355a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccdab50e7a68450b3a36194885c0c9d06934d67ee22515452474f090119685b2cda86a91206964ee60eabc33b47444a26da6a257b6e4a884621dea0c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea70f095545d1f29d44fceb795e6422e417ada7541d430ea48e5c9596db03e6bb95d49b75852dcdc7fb0cc6f6a98a3fd20d38d4c008b39d999525a549;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd099d3dd25c623f4571f11ed16b027eee23bfdf36cdc7e1e6cbb513cf73ecd97c39f26964096eb0afa1950fc40a3721b8ab1b9c460773e37b93bc8e58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdba3e10c709da143683bb0e2384c866a9ab7d52751b01e91e2d97dc8b910ce30090568d61d7a16ba20451b3322b3bac77f064d5164bdf93d61c35b97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85771c6ddacfbed341f47f8cc9c22203e8d552f584365163039e40656c8a24001d064ecbffd413714f73515d4752cf6e8e490edd2f2e649f5f4ef5706;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f2c3186b1158232c36c85c08e15b000a4bcce6c31589b229c19adf05f79e401406058a96851005bc1cef48b41f34f422e6deef2a30a1d11a901f17c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bb4a8330b919cd47193734a0a1d22c988608394d8314efd6b37b7f178eace6a482b3be5369b14128371b6c680827bf050729f4468529f053583535c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1bce799729841243dc98f445c88f97f2546886b58319afce861690c6e8e5706cbf4feb79e461c4071b7f7eb229943a0e3efe23a697735b1109fe50a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9f7b6346f129bb2afca934697bdd16121d99d70811157b50c8f2fe4cc112ae3c9c9d0ca49d47ba01b529e054b032e1a819e352226aaedc07476501bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8b06be95bd2693a9191a67fb39adf25d8ae23b27af4639b6752e9a8057bf9a71a95b725ba5e2368e7bf3d6f9eb6b1dedaf6a376b66c92d32472bfd3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32846658c06453558cbce3abcc4dcecfd34b02b5d05652c8bcca91e18edbe85a217b5b1d823879c2110d0e284356ccc1dcb580252c1b3c0bec934c133;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d37e6addfbaf7156e34641e066c53a3a9831723638f3dcd990a66b3ea6db4fd912fbe862ff284cb1657fa1a4281b7b1483e164b94348ae7610a5aca6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31c29afcf03d96705da3c44c161aa46a782e7bc6dd7875a0f5111ae4de4c7e2d65aec21638b2a5e207f10f37d6bfca31ecc2e6d0774e2b884f08eaf95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbeee2cb2efe1c94c65b6e097563e6962de881d51cabf6435ea2f5915d41b218789cb4934c9c24b3371042d49b51b03999131105525ae187b3f9626beb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h979cec77c3e420834b65e9d1570ca2b75a6eac4836698b4e06dd37ab84bf72787c461800f81d2cc5381ce80a15378cdb58e1e3e0d7640454892df4418;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha09cdfe6d467dcfc38e6f02d826a5fa3a3db8e5c07ef7bc8a984368de912200fe704390aeb61ce4f06e03e7cf551301cc34834c5b1cb6345aa32d6458;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c8a76057378c0604b791d21bb6247e8435e2da4d60b0e4899e9a5397489a9e975f9a75fbeca806e096ab6b60d9683c6e8d719eafcb982ec9fbe87f3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b704c359915580e92d7874fbd430b0334ee6119479503e568ffc1a2ef6b1e8f74df01155e2fbaaaff8c1d7f5136c485cd04606c287f72362ce9d9b8e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f712e4bf171288ef8b57a196dae2464a096197b3d8c4bf28bcf4d13029393fdfc843d4c9a13327c5c4d103375219c047f531247c6a633dbf3bff1920;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59e45bfc00f1e9d1376b43a31377e3138b9d50612cdb4efaa499fb97d85a48759d833405a85619e0ce8da50cf9451a056a36d03cbf97e3f511560f675;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40fa930ba6c410a762b2b5f6b62c6957988a07373e26969a154743371a4dab5761c62a5d831053baafff21be9cf95a12408bbadfa842102d9835511f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f77b539d5bcac11a910f830de78a47858c6e66e184d1990302dbd8e10af5ce48b9e31c854254dfc964757d996d2027786c5b9a64f72368acdde094d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h699a749a4f0285f6491e5b18204d0007d3bf664509d65d9e823118fce5f3d131e1655d5007665cc78bf1d899257a1e9375c18234ed2414ac6e42ed850;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3c67a1a0944418a15ed4b857e06f30485b56d9e480733ae493829395f89ef291a7cfefb36171e7b3df3a0e94b949e5c07a50255b92a863f353c4bdfd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9f257fcb8bd284272d81997c7c24a47df05739e221faf3b9295f1a28e98ec310360b94ba6bcbc6b6134c70a0fb6ce3f884ed3b8325e41961e3380d30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he320ac197438341282e751d251140d782c1361176b2c0d4b86fa7d9b7f5d1b585dbe32035b0a3c4b76b0e1dd00b84557fbabd977e616e5ca19df2be1f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h584eb56ff3b51886b0b1990f501bd5b07b2b79dc08fb5142bba1f5a0ac181ad4bc7cb00e16c52c8dbfc71ce7e51b43e9d1bf0cf6452a2eb3c159d04ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69791618a63d2d83fd0a5f4705dbe56a6bb762dde8a078e2c740393cd76ab9124965449662b34aba5586f476d4bb5ec0150c9f30091ab6ff11ea7d959;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1858566e57eaf87ed1e9d92837af6a5af29a46c020d8c79c4960fbafd04587699a1b7ef4541b76f1bad1a8f1571bdbe18cb33c7af359731bcc064aeb2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f0751c5f31d40e1863717874efb1f64920235e45095ba8a7feb6bee574de5c459704bf94ad1f55c85f34f3134d477eba60c7ca7959a0b143b56c552c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf25513a70acff012d3b0fefa13ae86a6641c029d312bc9586c36e0f2fdb3eca2c0c266233b3c57f173302e363ee17feb6e9f696826eb926eddfc0e34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274f30080aff65df3841d7d47f3d0f727ff0c3ab77e93c6a22521967f1433c83e193e180cd1f97663469e8bc9e0c18f24615fb285740b07e72ba65b43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdb329aadedbc0856eb8592c14c8228bad9a249b8460486603bf72344ac199ec4c0df1f92389009b5dd41adb9c6f406fcaec7247cd9f1488dac401c9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd02e719474d439d72e02f583e8bb2a76f78a150f6402c10d8c60c430e9e930ff88e09552daf0f8f1cb6063e240a011d6debf641f8be872b33cfe0ebfb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2fcffcf815c8b614440a50b41f0f88c9c47cc7448cbf82aad1f73547aab993f284d8429626fab37fa4124d73b374b3fe46776819e6bbbd5fa70e3b1a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf039490106f630b9b50cffcea4e5c218fe196634cb1126fd2b4d71920a72101791ce8018649ecae4dd15e6f73bed6432565f33a508fb8e2788e363ac3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ef2f1cdff6cf37b7daa5634e97bf7b88baca75a11e2452a98e67d4e93a7ae20fab274207c16f113a37bcf54656d77fa4025513d37c19388c05e17516;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h707006c2fcb1d7a9deea6d0171857d698950fd9ecf9117038695179cf98dcc3cbfcbc7dfd3a4707fd6f3c38c9eec69aff2a56487675ffe39843cb37ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfae84b3b72cac74412e17d679210f324b1db9cec8ba214a0a82270ae5a5fa79c3cb28815ad6f3ab5c297b38a810f79856ede76c34c5398e189fca9454;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he438dc9556b1c8f055aa7b1eb71ab94dfc8e57fc5fd9b9758db1ff62d27ede9edf0896814c93e6f23be6c8d3e382c4b6cf5e3b9b1c471d15a237bb942;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ed38eacc6f103f7443db1aa95f9568dbb6c9b7055e24822fa441b2cb0211683d97d0bd1a28d7820ad4c97e4804c690da3a8a73408227a4aad0ba57ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec7a1792039f06193acc38a3ee0ea007c540318a1dd5bc32b69a1f5042d741b33af4ca413cb9e73a4381608eec694d322121765b6cf609ba8ab7262e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h102ea3971cd96eecf4acdaf0ad7b3dc2abaff09e7f146c601c48d9de75016d205a2e60dfe293f09201eadb0052f9cb522cd9af6d43d6ef6deb83a5aa7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1afd55d287e8366dc659382e2efdce7d1637e87c750c17367bafbd9f42fa31c5e1609fce82812b8fc2a02b67d60d53b4432e6c400669b9f0cfcb6162;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc78456a6702766cb972c9a4e08bde36e51567e70b4b0813ac770e7716eb4178524ef9101de876dd0ff82f87878353e86c1549cb563dd97f4ad0b32f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf01da95cbec037134ed260d37d0d3c9f624c424f37abca6116dadf08f2ca7097526010e9b0f982d6d29a254a6280930b364f2cd9999fd720a0367ab73;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13e7ff33fe58e60d1ecde77fd1bb9cfb66bba6e04f01dd6024d1c1b5f43a9ed2abcd6b1698844279a9266eed1f8a34b45a0113bae064fa4a50836c8c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h346873bf0f054fbd48cfc6bded9942d70a5115e51449eb27b1950adf70f1febcc9caabf59965b4de6c2565c21c14dc84625bdea3357cdb4a196165fb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8479da0ad9074fde89a55df0e8d5add064cc2e57bece3f241231510a967db7f295a5d0fd3dba0128f3b8c61b63610eeb2966a05ce0f8c2cd816f8a2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91891ad07d8af223049fda309737769aba3f7ef13513d04c28fa1424c28ed577eaf1746697a7589aaf7c1e666f3e59b8604abbf8441181d6594e6a34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c2895110cf946831be3faecde9731ffbb84f762c39c448232dd1ddbd4523d45e0ba4b00764deba45629aec0c4319739909625f3760359dc63826baa6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h223b23d979fc391773cae62ef97da56003e555f8586536962724ea39a4f02545aa5e54f2f5ab69bd8cf022a953b347fd5f34d739da08347ec99f68287;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4e1eb847f945fbd9b58ba0f4d0d0832ba1cc41fcd0ebd34e6a4425e3b03d7bb7ac27f7b656d4403bc6265f69d2d5285c35c6e6decd98c2197c809690;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6aabc53a17df41ae567e5b3e6625e7ce8709b7b5c6a531b2488659fe61d2019f3aae5de75e07c6014ea76a28118c6355710c619228fbaad13c2d8fc73;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f9b7938ea6a99550aa54896cb102f10c707ab9357085acd3f525dacc5fc8eaee24953caa6d3d81c10374fefc0d674865303633db89b671f3c9151847;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96b4c69a6365fc97f0b33510f2fdfb9c3962ee8a6afde8f6c033d67d7f9d4a369035183be724abe4bebf346016382f456c09e5383c67316a78fbfc222;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b129172d8d97f6af10807b17ed1922138243fc8a3762fabf79dbad8d88dca3158950557ac72df922f22b55f3a45ecb29a6cedb79c19203a792c7cb7d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37666126897f474e0763b619b5c4c973800bf0f9f03c9319855304e2c10e2ce7134aa88387db669aa9e75eb6dfee9fa369b48428263985179d553cca4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd12a5e58d2c515b51f7151a8c089a1e8f18406edf2d210c6c43b6c85d6a29247e6ee8fbd964ba957322867585ac9ba83edac3a75d013771e731cbe298;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha015efb81488cb01453e098b21a581824577f26d5cfadb8a70757a76fa90b00aabfabc57a5fd5ce469f765f11f8efec86584b4c13706eef0f9210ae2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b5bcfe7691e5bb0cd0ef89be72d0781c27cbe2d3790843367a40a849d3348824c4a9d5009a0a0cd09fbe74a6659f57e07770ba616593a7dfa8f197c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36637fbdb0d8fb7e445c81d1769e140ac9e3f5761b60c31a77200bf14fc40c8dda17459e18cea682b3293c14d78b26ea1eea53a71046119c572c7579b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef841df91db69c5c444d87eb15d72eeed38961d3d4dd9fc630f749ca8560af66128a2fdb093e5db436b2a111f843bf67e5ebac339c44e93c30fd38e44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had912b70911e5ed77338cba44fd4d4a4a91d25c0b37f12a969128d7ec7721048b70d43409509c48924f6f6d7b868d6cbf0e96a5aa1422a7165fd02fee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h601c4186bddfb7a7484c3d416db5fb4d24256e6b606012effa3d1ecb2f4b252b91be8d3298b19d5d5a0366be31528d78f0c66cef20e8a59bf95520719;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe6f719e8599db7ac06eb0567fb0503c2327e0c5d0d3c4c26fb89c53acd87508000930ef1fc49d7e63e5d4b3d63b786276e827427974615cc888d1eff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37de7e2625343c18526f83800ec78dbd6d4f694431a3fcefe19994072f87a76e95446b00e9c1fddcb600d60ad27f27b728e52fb262ff105a9ea0516df;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e37597a837a332cf33ee24b2235076b3c6a5569d7d4b97636ce6968506ba7c172d1fb5f0ca2eacc11df5ae507f1040aee73361001cdf3b55be43cec5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dc6bfb4066eaaf6acc860fcd57b85b6030e8a8b7550e52e0ac611a8ff34576fe3ec00591cc262cbeaf409f15c35df2d16368232f4f40d4c55ce5e844;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b9aa5a1e195f8db134f8932c030a8cdc2334504c524f5a6dff4da683e615f8be627deb725ebe01271ed596c4b2e63e6071df47f83d4417c3ab9a6785;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b307cfe8c7b374c8622da987e52b7025727a4de8d1243f13d9c473124dd9a1a75a142969b67bfe8e37a0fb550c5e1c39c0c3b17fbc57ceab0867603;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dce7b5d67925e4ae5a34cbece3f5fa2f95fcc7f1c32aae1ee1669d9091ccde5b9236db584408a0e2b092b75402f74cb1ddc0873c389d523c699ada18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf84743fae5675b3e4d12adb7af7efe12212fd8946ab740de9b606b710a953f288ddfb596c7bdd304f6b77f272c2444fc3819dff3fd14b9f71abd7cbdf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea47ac5ee46830cbf8927fc884d6c14615f3d8ebda6930622bcb7fa08cc15c798277e69a3d0744719f5aa89118faa7e4c167c2dbcdab91ac712247630;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h625ff5c7995228e37d1934bbbd652aaea2b715b7af89135de7d9bfcae6ef9b222e23dbb6da093a187da831b95785476da876953066446036facbc6c6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedcb204741323f2d78d692275c16994687712958353ed8fc719d38eefa4af33af1df57b73593ddb9d6b5129029e556179ec38d6e43d77a98335d62e15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e6d9dab7a4ead625a8683a3d1cec3cff221fbcf4d99d72307ebea539501985848094f66e6f09572c65652384e0d13f75c647d980e4faa9f8ba3420f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a8973b3fa980febe314405a2248b3777b5fa8ecbc96e20296e3bc53ca068f8c25f18cb055f46c14073ee18f4c223ef49e22ec9aff78565a866d0f842;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he05be50062a5b0cb762a3337b27e9fea0416e34bf268f22c0d2279b15e8d8645c963d95e238a5a77bee7b91d62a1888e149399c5b9a15f739cd8773bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbac6507163e7d5c6073fa7252e48d9be93645210a8da82e99a352b1ab15a45e557092c43176c2249024a4821b29be9b386b99f59b376ddc8169ca89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbdcec60dcde62f41d015ca01c59f775c122f8873395fecbc1706900937d3c6434e1ee4d4bc56ab542f0cc128332fe2511005b4425e83f381360446dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fdb85351fc7b1d997c18478a2192b3e0603bcfcac09dc90c9338ad3cd9e0a930f9c435b3a4e616c10e2a3f0fb5db90323d374b481cde9f1699831dd5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2de1db04d8c3441e56aec49cac4dcb96964bcb94daddbea292fe758de9c89fb57c425a6782f49cd42bcb606799ab3d189b5e5acdedd9be5a393413181;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52763092175c26d035e03350f0461b337f69794374613552826f916f677a0c74a1c4fb3987b8ffc3caaeaf9cb0feb6e2df992c2ae32caaa7a65538868;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1056ff73f24b0ef2e400171a2118313323a4d67d111c3093577fbbfb7e46f014ecb3a07b217904a311138b20659a4149f4900111d7d6254457b8e8a1c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69a3c76f00d5bec76d36bb6688ff29d96aad708d86fa0a3804d8345af3e6ebfe5bbac9eb540d2296d1069d5750a84bc0204e882500fa899110827de44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a9eb441a70e4626cccbebeace4fe8b81de6cfaebe3f449e1f321d3986fc6d958f3598bd262e850e074e86e491d3ad279dfcab6d5ef37309bd3bb4af7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8f9eb56a66702fd2df3d1e45cbfcb272de6a932d5de08c9412509a77265edfd591a42549e9fe0ea1f54f941d67790510b18ed04a07a1cbbf4b00693c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he855d5ce98a05c6819739d58f0a955ff6e7719de657af027c10e8edc920ee9cf06d09601af9f22f8a6d1bf1490c43a545f666159c32a521067160ed00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7610fcac347a9aa4817b833d9517475ea597a1e1505c37c0d941edca29bff441333cb91363f570faafeab649446533658e202c5619ff311e0addb13b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52b3d203d758143bbf3ad7a4eb7cb637aae0eb754f7c3608e1da475a62d3e59e5b9f38c5c1db7d64ff8f000b0b9e3d9f2f3413869d5f5ebc7ce6cc625;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9c3a12d330fa23ad69fe93ed5cbb5711d4d050a36f13fb5d3ad04d87bec529330950c9e3d3fb4877a12b4708015f18eb09c4225306316b87abb84621;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe88229b0c64c4f37e31f2afd19846b2fcc3a7fa52a20513c9b5a23f43275692d8a9af66a6d1441847aa7801101177ba8cd93e181a4c6361723d656ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d4c861b521a3a7509998602281fdec28f41c75e0b4b9b455498ad12832af9004a3eb0e157cf1ba32a7650ebd11bfca9637eccdf0ac8e6c1ab1c65c2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e455b62961404a11e062a24b47bfd4d601a358958a3ed0fb0c52bd0d258d2c8b332d26f2f47f444fd283923d160dc82ef387ce6bce090966346b1880;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c98c86d4b3b835692ce8ceb7a3cf664c76fd263f12e178dd18a024d092c0b2051217ddde7e73814ec106991922e0b5c0e12349065dc88f8afa16ee24;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76dfa296dd210d4aeeeae7062c6f866ed70da60d0ec5edbd2e466a8e1f7afe067ff6910d3fa742a8082921fcfce2f9a60ccd382930a9eca1fa019264a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h517282672b12a49de1f5d5e7f53f43a94bce1101c5c1b39b65bf470c0712b6d5feb21e93ea7e7213ca35d45914795e75618792da67c232bc146c6fefa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2eec2ac82357faac40e3d8f6739a294aaae6e1c9c4962e7657c7a1e787da784b14f8a40276932835abd1e683acd16cb3b08ba8f79d0762daa40ee6be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1588fbf2600793c80377a5e39cec8418e4c34cb3f7786b23bedcbf2f7be573f210fe91c19da86486fc55927cff0cde766bfe32964e771eaba4314baa6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h745e1840536d8c68867f5bfc69f74b079d809dc571c3e4b442968f427194acdbf742151b36e17405c66962a3408550c31af05e00f9877374fb63fcc2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28758f19380f055f74bb539ffcc24f20b614a4766c7c34272060ad789ce5212dc97dfc8e2644c183fc016701ef3bdc36566cc124c2ae60649a5d84a06;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6ae49fab47615285d11b30360ec548338d200c123e91fd739d332d71b62d89f9410e1f76f9253ffd678f0fa20d4f3dd65d2b85a6a70752adc87a78e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbab1a6422a0520e23448bfca64d47487f4881bf6664618b86f52843f3caa639aa64d3c7d027cc7a6c34b0801b5a9955ef96b0b7cf426f89a4315dbc2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe6cb65b85dd38d40262070f5adfb278424debfaf8dc4e5562aadbada3fcd5a03c88cb79e4152af5a52147b742c3aa7bcb08ca22cf2d9ce4f8f9091ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85733c818c749a135d71a2d1bc9d7367078212f33b8939ec5b4bb4cae5caa500d697d7a2257086d8af5beafaf118a31d091af7db688dfa83dd1b1c2b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h465034972a006464c7ec584b956d3486657de5757470f366367a49ff1678f822de855c23dc2b1fbddd99e9b616ad910d8124869fb2d897c453fe82d68;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he15515b9b74fe81f812dea4dab1dcad3aee232dd882a617e774b66343e45e1ce146b560639086f5e1af691862d3af10dcc123107063e15c94aef13498;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha320ecf780becc642846237a909de12358449ba905172e7b6a585f64251509b8f3b689b59cf769c5057d08089752525ba3b4472a7fe3e76e5bc527d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h908ff3ed55be95556501f36a8958f710c6e9a8246c776f3847b21b62eaa3d31b926bdd317d3c3f367235cb9943eeb0517ae559f54f3b8ab73a373317f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7ef5f4bb742ba0b3d0b3e8eec70b4bc75230b549d76d3b48f1a62a8607591042959ea0bab78361d21209b4d62bfb10d36a5d099ef1cff5394749b59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33557561b48d11af09d2a6d12515f9cb0814edfdc85ed37853920af1c071428070f9082bd954df60596c61c6f1367200887111f73b2aaaf24f6caf30e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7a059edee05c70450f2c8b393c708d4f89c3712280664d5e737013af8d217d9c983198601a07d7700f57b76291b48998a6c31bc0728c12827a0ea221;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h884cbda99e0d604b0c46dc68561a383796369c7dfb22b5e9595eb32f27a289d9dd95a4f40c000d10d199e9d08ee5464090dd1179ed5cc0e85105ec599;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2448a5818556088936e42f2b5693e9a29a9275c6043904354cbe0f6346f28329cebdcace5482b4ecc0ba6403c4da9ada97de00c9f6101efb8149d3442;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fbc8ad4df4476a19555bbef588cad78b8f022eecaf92fba6301eb941a3d2b709954d2720b35f120c1bce41a05349ba7795446e68b8f45df13fb66056;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82527e2540ce5c96de9b93207072b04e111137cf6da98141973667d48b94c128fb2a7394a95d6dd680a8d676cdc97d943c09ba4e7a66dc26e1430b698;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67a31ad4c3065da32cd6ad6fe02390fba5c16cc51645c9f2a510469eb9b70ca6b7efde7c6c2a58dc32b2c6d21968a3a33a9bef5364554692a50b5606f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea93023113f1cb14ed3d9429c890172b3a0025b240e2a35459acb812984dfac6c9a3887afd3e7a8fb30445da72389518595fc725f343895397e9bec97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1200f1d63c9654501b379044a9947e512caa0fe86d4c1a9b91e6c98d02a14fa70fe36e0cf7f9d27ae5f8ab6993808bc166954b49617f9124987137034;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69d47c027183bf8c4411702448aa6ee998f104ec428361cc2ba91e8564d08d5cf2bc5cadea10150fc15b5c1fe4abde4c5baa92ba03eff95617bdc044d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8782e2259478417329e24382282020d38771195a1eed220e55d228da18001c2d0a39a648277f6e2cfd3a746a1a12e96144b7bcc73d76388870f7d0f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h627a08a76550cef75c531de534be0b825bbce420d11a633f3ddfc1864401f9d1886136bd2d6308f8963c5ba439499d5f5af4330f18e2e2455010425b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f9f4774a7de02abc98ebb145d6add0744f124ee632181ba5d1651509e904266afb40923e7fd3768fd1d6c68c405cfdd300f3fdd50f0935980ddc844b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c2592bdd11cad933b4c75169178ea85299da0c65c1791084c13ff689deba64d28541761dd3829d0e54d2f9d321e6484e7508399ee9358240b155528;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84c89fac0fde92bcde5278552906d4043af25bb970dee6720401e26573f2d5744f4d162202dd2579f662e517c86edfc44f8aa532130cf2989ac99502a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27852dde72afd620855498fbdd22c26444204ef54c471e70e5f35011d2a74eceaf61433f6544c4fc4cf8fbdacbba8bd50e8f55b3615074438b77eb933;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbef71dfcb84d70b93cc29d704d7f0eefb9cae1c41f708f3504ae67871446a08319c138fe74f8e5f91368cddeada4e565fdbe0dfed2716080449ae36e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5df6a50a9cc5acbd0ffe2493184a2b03a175bf7ca1e7d92fb29d9c30d2de101945508f7eefc1baf55c2bd626746a03483e0b030b377720740f20c63c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2899b177c27ccb36cfa4574f276fc88e7992927c92efbb0effd2ca195ab4e87d0d6cf07fab5def39b57d848f030faf72971c7cb3bb99de42298dd0ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65b50362cb46be38974bb17e1d66c85329b5bb00c2ba0ac0bb8a24fa97215ae5ffe9718c4d64c647f9be088e7bad6927f39dc265c5799296211adaaa8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2129e12b10715084f8a187932c400d590e66e66d45df370d1d33ee1afe25e286491a0c5100c04d546c47ac7257243959af22c43555053ab2f50968be5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13b10d8fda741ebaa7eeac2fd40ce0dccc2b1d61e405432f59f6ff9dd2f82802ebdc7b730d17a0cd957df3d0c45e26bcf3a0ac658f453c95b5d107f71;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d3585a53f0049fa41e76b0015eee98fb45953257a6eac8b3e19a7a8b256fc113a8a97af313b95b675452fcbd456267e845c6a0c7eec8914c51707755;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he561bafe793ce56119b8ab02e26bba7996d38e76fab455242498b7a34ab91b08601e05a1665a3b1393b8fc51c8ef4e5dfa22a2439038839b2f2d8bda4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d71c90c7eb9718ee2b0849fd2b43f3ef00e8bcace42ecc28f140dd7d995e3932345d8a81918dbd2b68fb1c87be0a3372d7e8ccebbd52092e82b0cd57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he28bedc68cf7ed1b24a0472e77b43f59896feceeaa6fe1c5b924e7ca531b2f050d568ff54e0dec84fc1c5bdcafd0096fcaa5ac9782126336c6dba10ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb542625d4840cb4f021c73c6ff18d05baba2c8a9b4c533af74d2c221e55a48cabcecf0b72e2b1c7c68e439255559becd56b26ad93de70283186fdb27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e40c12bf8a7e32f04b03447380c8911ea43884664b2c31a6351f4dbff6d264db1eb7b670c9dcfd3142cc282fb58f02aadc918b82fe2a91703495a65b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbec2023c3a12ff069cd3fcd80b86240fc4246820e51dd340bfd3be79dc8134a5177516573ab05572101c029da7deb3ca45be8b9e290285596400946a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33813ded49e9b23526c01337323b66f194f5966a3c69f1ae8240be746499bf286e86d06a3b8242f49f136f15f6c356c260c7db917dcad7aa2c399c97b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf268c5d07e56544ac650494e366211a23f28442dad4d5d70d247ed21215c9f1656e7acae0eeb2e367285c9cce96987b553cfcc5b8f3ca6f9bb32ffef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32a6403da4b1cb8601db343bf8a4d030f2a72a7b3fd9e6aec23d1f8dea82277ef9ae48ae1e6971f61513739afc768b50b14808cedfb9a35963ed333f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd234f7585122a2fd16c67c945f6aaabbbc1740bad10229bf9c8faabceaa3346c823b0696ac1b694221ee6160256d663956dc7647a86db8e46ab105907;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2ed9b12b8e2df1fc592c904cc0bcec8559baf2cb4fb5a338e7abc68907460f7fd99e1a4844a38820f46bb66a7b5c9cd084dc3ec98191659a91db9b86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e391ca2de33e19d6cf2a42754e72a9a9c06f1a1141407c22cfe7fa5225473ee511f5537a87ee77d7f431a54333ea4b7672ab6af02c31037b0ead6aaa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h165a669472a57b076fca8b5222719464cf2d11320b24bbacde9860d355130bc76c4435577504498381ac6cbd8a7ca313f69899454efa2a034c912c9de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17de06cb986eea0e8b67d9b9df9f08fb8b38bf45858954590e50f5436e5de6415d0a9885f32c4bbc5ee9d612157cb8e31e3e8570f5dbffad311780f8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb61eb3a8a26602c63cda130cf847db6b00524473985116a1f19e56b853aec126294a63bb1ccc4b5f5e632afb63ab85252f4441f43f12e5b477ed046b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50e0b21d5cdad632458245e9d2570e1f11839158e5b649d7c7028146e51aee9f1d807029f5ae96ffd9c27eed2226f46a1507155f9919059e26bb0f113;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd7b1047760343d0ee440d35fde9881b6e137a66e40641ffe1c65551c4e52704ec4de063645b99c71164a1b39b20fda07d3dae39bfed0f923e4617db4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd68093a5122f2f6ff1c047e08149611fa1a452ba5d468de8a6e5f392a9f59b8c59b32fa0dfd0a3f2477e0bf48bf785c36455bb557f7dd5791d1f1dd2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e9a28abef725f7f39b1111fd3d51fb37a40f3077211d1ab085a4510539144d155b602ea0d893ff9a82cc84e2983e778f107e3d7a294369cf61374161;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1146214b1cb89520d60cdbaed9832842fd1dab2d985c5430224ed397eecd73af4fc30bd45bbe1958ffe51cdcd62f05e1289fd6092dd044cf7feeeca3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb83805cf3b4cbc6408e72c22e63e8e4609cd6a0a53bdca34e4b995eb702c3078fd281a1a895c227b1105d9192c24eb37844b71789284bb3be995c4a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2ad70846d5005e1ec4828b72935d8b2a547c2c5ad0a6db4ae5f1fd84f69bbd480b52ccd0abafe6a0db057d64ff7e3827a2247440850d48bf4bad5349;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7ff7e37371f86dd1c1e151740176991bbe148e5f17736b272b0db1678ed0d1058d4557df443c207b7a4755d19ca560b4c97eb16de20b049772f7a649;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa348d861228f0c6fc5873c85259d9c984455907624e07738c818a31a5fa6653a9f24a946d139638c244b777cb8c4b04f428f71edaab49ec3dcffdd3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ec0afd153dd4578427ffe4434c54760fa53a90a23481a1dc23cd3a66104f0d34895dcc77302d9e758b7e4dc2b1e2433142723c24d8e94efc287b0ecf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc250ee63920b432ed9ac1050597598a9a0fb7eadda52cdd967931a95cb861c9e179c0c5151293dcda667012145b8103ebeeab87deb9e03ae6452ae00e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26f667786e2a4e8c8333a42282b91bb03b48208ddb4a776a80a59e464cf2cd47b0668f0b88d97b5ef3efc911cbfce93b61334074756b991c2a40b224e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b4f763a4773f93e74bad4d8a08393d135911b4b5b4210ac143c6404ae6fb2e2cbc0437dcf3d5751c9d91096064311c5c6a6231de2607b5ba56b4bb06;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd1a3aa5b2a5fba637109a7f34ef112ed2a40bf06f7ec94f7d3e99dd7f1050c8566ad0a01a667c324af3b24bd84a10090c96b96f7b6cbceeefab677ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f276ba1c389a42d8640917869721b02d72a005d48f5416f30a13ed70db8fc7504cefd613334ef8a866d51fcbf069a76b33a38771827cd221690a79cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0a8cb2a8b8256566f87aa4974e38997b105137d415d41766f7c713a9fc3a39323761be19f5c589cd4ef63703e3b5410ea66af4f111e9bdebde90aece;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he29258b17134b8b359d5f262c339ab96b1a219a05b320ec5e6e0183ade1d7c61b5ecf391e0abcd26fbe9d040f6156da29569cdce35d264c1d74958186;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35087a8cfa9584c4061e064b2ac1c3b5305e791c3cabd41c6de84f226de37c0c0c52c245ca806d5b1fa205e6c742378adb069ead04998d1e743177546;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cdec906f623ee17f977ad957428d67ffae44932976090b71c7cef94af7c72b10ef03c2e848c36a7a101a23256dc417a85ba2e3383bd533fba3ae5497;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e5dbe1d52d420b6ee66e5dac8884911465eeee00ffcba18922a2dfab79e075b5faaad3073ff9db1e18e347745fef38cf804688357738bc3dd114b96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bc49d0ffc29b817337fb36d06ce83252328d38718ab8196d86b28b6e53e47e684b984d26945d53c6920a6e463db74989b45be6f4eb802a86048133e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9893d11192a1cc56269d3f576ad9ed5de9d3e5f5877eb0acee895f2ccced55912601b6fee7b8497666473c63acde8e70d14414ce4e89f384a80e356f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4d365d5d701508bd58c5fd71ac0126911f29eff48e8a4c0833d14e677d365734eed60430bf7aa187c2ce7cecb9401811463f7ed356f2fd94703929a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c19ae342a21b419ecf056f3fa1a97d0b979bd22680dd9bf37f74c1db69c4f8454ac6a317bdb413026000504c84dd541b18e2445e90b6f5410d217f44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3a68a73aa7f7f1b7e8fdfc30c3bc6988709661d6e19e95dbf6bfcd6e11d4baed6c285211b4738dd4c3a5258df23960d6a4da8809c99a5855f6e27ba1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17cd2ded38d6d7d8301d3701fae270030a75ce69dbd0da6922271bedc81886981821ee15839f8eb973c3a892dad1f064ad5eeff8e1936fa878bcc4b3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aa12111335474bfcadfba4ed9bce78946cddce3196038a3b461389c69016f224556183ad36f34d4d76b46143d9c7e6529aedfd4b42cb842907074ffb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfae5cf7a537dcb5ab8e4e2d3efc65be78caa6197e7fd55a369d6847495e729c81d0459f8617fca51ccfbf5c33e6123cfc976c95d49969c4fa93a4fbdf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha09b58094caf53952f2afce6d1bfa5ec014e579a6baf07aab7c383c753bef7a216295d886033357a85071d7b19259d91b11e291b2bc6f3dedc9f71a10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dd0edef28935a4bfcc0c21a1fd272fb8b3bd67c104c0997b0bc33930671f3b91910350880172a032b95588d0721cf47b35bb67887e6ef38a60a43a2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a8d69eb5723d3d7a81169c56355b600b756afd56e3f3ea53b733327af2f386c6fb65e16bfe10dea027a0cd38c19b9f873f6b1919afc878e7857831a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf34f6bd6277a6aa4f3e466e74e74d595855808afebf736ebc5106b66e493b8747876e2c36c9a2b8aae4f42712eb63953d64e43cc46deb4d01282e1b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61828886eeec11fd14ab26aa5c660e4c17ccb50c8e85617bcd4fd75c24eb041e70401361ace8e825792be9e1d45d653f70b8f8445755bd1b72cd05900;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h411362a0e89e6019b49717a9a2a4a2c7db02b2bb5ff1820c6b97eaa1de80cbb19e0bd5c7f86202ec8ea5902249dcdad9c4384333e00372da736565471;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3229a6f0871715813cafa0eacf2d8115023f9117a5394f0029a1e569476f8f9df6fe99333141b2fe29ea8ee091d3c73c2a3e11f33dbc37631196237e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h194e5b7c5cb9d47c4839d6c7b0340e31bd6bf94539ee9e2471f5a7670549334a2348b44745da79fbc9909f87e6304f5e251ecc3ffbd6ff14ce69fb820;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd1db8f306af2e56051b03d6d4bc285400fa3ab87a11eeaef1a1155e3b3d07ecf0ef71499d89e656b399668147d269554cd81a10482d85b806c022382;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb475b4c0a1511fb2c925d22ca6122fe4d479625d6629f2b7b9061f7c65767297ae70a7e33e719fe53f96e3790b3b755a762814a27de6d2e770c13c235;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21168d529feeca5541bd428414c8fdd609b54b118eaca1fa3f247b8c9dd49c46dd3d123a759247d60a5a58c3765b52ba404671dcae4b31914a95769c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3258ce682e04979cc5c9dde59a2712db57681184362e72a8da31b5ab973a72d032b8358738f2d6a755c19e590e809c2e3ba971fb587b27b5b72a1fa4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e60dac1ca963c59d4735863fd646e0222941f9f08095843affb44a5cafab9289be214379be2146c1e657df718f55d4caac1d5ba4f92927eea82d75fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf76b21ddf90a3d5e5eeb1342a007ad553670b1a1972ef5f885bc016a0157cf83813c425f34e676456c67ad17fa77b5e5555f6298da7e1ea4a6362a3e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ca9c840339c585b9d3a97a69bf232d93e02f22abef2cc2857ded2cd64cac183fb4e9ada01c579c621a1647b773f06b503c0e29976cb310c337918d0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd28877d8019da235bd39b89112d2adb244a6b831ba77f40b1d1c62969ebe255619a123a8057a384ff7f8a0da5d63b0afb72f1232c6c921cba441326d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he88a5576a38cdf5eb65fdee02c8b27f82edf29d46db2a1b0fe5e4a4da65e089e57fa2723c76742135d06d783779d448488618dd56509c303c45ad3653;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2572f385e1d24268cd933cc53da67fa97876791a45c33f7dbfa1ed6d796183af93ff929df5d17e8a4d74af9b42635444ca370568e623e3654cb22d09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2afb8e7bd560f5ff21de14c3a6cd4f799f286878427e14fad2ec952f9cda57a36c0b93ac5e4380c7948d25c33acb864019d9f488625ac9083a5b9df15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0f4ff57291658d22e5a883df37e663894151529d77b7effad7c14359646726ebb2675f870dd01462b60c9287f2721af6b42957487f0bb30fa1636d89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1b98308f356f34394e6b0ff183197df8723e13a1deab13e7991dcc856f1a0dfa53b0775bff7ed1da6a42e72b75775b93cff28c13d33d5d5baec644ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c6ddf0a065fcd5746aa74842f65056b60b787357a8ec6cc19a624b2929deacda1250e4b5411c68e2e04b24ce7cd9b533774ec7a70eec6c96c1535d37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8325683a7f9ed458ff044caf67d20e30f2ef6f974c7bc66c21260a578e995853e122f0fad898f99f4f8aa999bb2eef3268d9f638fd3a8a7804d40dc3e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd37c46a516cb9d84ec8f8fe4640e097840b16329d32d4f3efd5a440a566f4b40ed9e6071299c5be56fde2ce779978aeb7f6e56af0e123d21e5d74e5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4dcf992ae6ded3a4639c7f5cb424e7ddf35d409864ec3215f9bf0f3afcf557c523805f4cc9bf447d513328850c65c0b2fe22a6e929162e5cd888bde16;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd36faefc7683186e94c59a17b9622e7b16451eb8cac4b258580b7f015ee5b986b6708215af6aacf1043ecec1f889fbedf1837cecb12b0f8cfb3a29a11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3d686e4dd07902d3e2bc7a65dede5f9f2b5e68e53981ea23289b9dab52775f6e5d676ca7debd4aa87b1f243da1b144e5a532bd6e2081e71af29f2e3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc68c7c54ddf49816bb96f7f8f471aa9f075b3057eb2932a6d482fc20a6a3eed1bb9e49f460e0c518057b5434a1c31b3221d2d7ed1ee727b55092e3e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c4e16f822e4e5d37ea521daf6c68542a202aa3389ac65453db1c38b4085e0470d2b571d2f10c9b467858e413c1b441ee7e7c951b62574efe2377b317;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4c8c4e8f2e6677f3ebcbae30ecfa07ca86ee556cbb44ba5ed0c1ad732ef448bf850f8a1144c56696f9a5bd0dc1a64a576d94b72fe26aa6c69a6843fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa82f6c93a9433178c78396d1469c27dc47c7a9ea6961f7ede81905e50e973e201ed549775202590eb9eded763e98042635fc18850e2b512bce519ff0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc24667705d550f9de666d1fe962f6d4e3ba9823be9d6262a6dd438f072a79de2c9913b50b26e03fc9a54eb3ca74b9793a79589d65aadfa5b5decd3447;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5cc87e5a039b967c644671d004bbbae60879a5c31933c40f9c92026a2b335a79d90590c07af225e8d4a47017284d91cfac53997a404d920766542626;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67f6c9b508f56258ec461b837657ffa115b636f0e46617d89db20878d927f2a6b8c8221bd5a6280db661087b34a32993032d019102c556863e6df25da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f5e7d3b6cf31d5cbcf9591498f11f1fea51056eca88cefed971dc1f8e29780a979d6486630a17085081b67b57b87b468e25ecfe2da35d652a79e61c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2697bb0e3824b91699b8ce55cd57b8e20b135d6c441a5ef63d914a57f618b7523081fbe7e33cf3e4d7fb687e1b68760a807b596746c563d2adc094bc3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37b3e4c6236a58f4353314472d7b1cf1361b06d38634c28dfd69e342fb7616b5db7a651c92831da5d69e9072d5197431e6ce511f900714eedd7109032;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8610bde4bc957a4764db3e7e84e821cb6d0f604c6dbb1b6a0fbbfa4075e50368a30aaaddebb536043b6fd7e1d3be54c88b19c1d4cce2270d3ecc23473;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0563dbee83eae0bad4c91e607c2fc64f621a413ade6d5a823563bc87a96beee6c25d46973c9f179946526bcedad24712ecf34a198d9bf437be400656;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5816ac0334cd56784dec2e7cd40f943fbcf6cc43482a2cad65be9fdc8a733648fae332a68f11dd2681ea2aa35a14f7fee9b10a199cda94663822085ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba6400aa09ad0643f190b9a1dfc053eb02fd3df40aebfcbd2af2a0460a5ce9a77374a28309640870ef93381364bb5a2436978b7f59bf02131307cf859;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f5389edaa0e376dc531e645870861c977317e6b3d0c50a05a3cbc3785faccbb8575a6b1247f58d14a068e4f8d94e44fd077eb89e55a2a402205673c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92d4cb4cb9f7973955a87728b9fbd578053c2083507c41d19d010940ba5a6cd2a9df94df31647d4594d2fc74095fbc92b8282bcb9ae1d8a965eb8dc34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f92ded3d40f6adf15972e0ae6bd89a735f66024e84a70c662edb07a6688affa5d1326b124378abc0461da47573e133ac43ed18a21b417ff15fc8d157;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha852d6b419fb11ac5c02df89e0a7445db0e325ba2038912fa448352925c0e4d126597382fd8cf94e2689d8f6305403cf44d24372ab3c78a753d8ab6b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3e4c40c0d48f9549d5bd693b8958314494b01b050cea63547860b8072f551a50b1ddf24ece83052ee098bb592dbd56dec65cc7a662a1f6749b0f9a01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd78b34c0750ef078c1f513cab230976a70e822db6738ad4bda139432f6ce435724ffe83ce941ed9a0160550661f10571783f1f193cb9d5757c105179e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29321497fe62ff871dca86a6f3e02ae49842147f6a4982445760fcb424c26e15f5683ac3abd70b996d8e09b3a8fb581cc5c9f04833652ee1b566e713e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e8d5be2b65529b74ee39d9a167df490030e4d4a5322ee539cecb90dd9aeba239924baecf46f8b62376d8fdf07bec63b6ec10a37ce8c2cec65ba38f60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h912ac12f11cebeaf448898082e5e82fd776a7412fa4639b39c34341bce5f7dae44c8df1688ba850117b437b68f003c05b8bd9ed6bd9de19d5d430fa7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7913b28d9ceacf5b4c55cfdcbf152c6dcbecbb2293fe81b2474a5ff8b02f63497124147274a3ae9100fe5a17d9ba2647cf04bfedb8071e798b712616;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd03eb0c3ed3fc50113d7bbec92e790b89c1ef64616bad3a19be9cf865dbe5ea6bff2d9f7a65a0486712f25b43dbc0b3e5506f78b2394bd480b3f8b8c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc6c6ecdfbdee61bba7e7f085a1fae2e03c2319ff597351551fe86da830deca441284e23f2b1dd476e3f7deabe06f73477fb632c714be882954fe2fb8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95a40e1fd4ccd4d92846dfa9a62fd8b29738d5062c3241bdbadc92473f618e5e8be342b8c079cd62faa79246c2b44a7a8c1ac6d8e0474b1b9491e96f9;
        #1
        $finish();
    end
endmodule
